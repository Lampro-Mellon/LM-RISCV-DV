//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_188(
);
  wire [2:0] _EVAL;
  wire [31:0] _EVAL_0;
  wire [31:0] _EVAL_1;
  wire [31:0] _EVAL_2;
  wire [1:0] _EVAL_3;
  wire [31:0] _EVAL_4;
  wire [31:0] _EVAL_5;
  wire [31:0] _EVAL_6;
  wire [31:0] _EVAL_7;
  wire [2:0] _EVAL_8;
  wire [31:0] _EVAL_9;
  wire [31:0] _EVAL_10;
  wire  _EVAL_11;
  wire  _EVAL_12;
  wire  _EVAL_13;
  wire  _EVAL_14;
  wire [31:0] _EVAL_15;
  wire [31:0] _EVAL_16;
  wire [31:0] _EVAL_17;
  wire [31:0] _EVAL_18;
  wire [31:0] _EVAL_19;
  wire [31:0] _EVAL_20;
  wire [31:0] _EVAL_21;
  wire [31:0] _EVAL_22;
  wire [31:0] _EVAL_23;
  wire [31:0] _EVAL_24;
  wire [31:0] _EVAL_25;
  wire [31:0] _EVAL_26;
  wire  _EVAL_27;
  wire [31:0] _EVAL_28;
  wire [31:0] _EVAL_29;
  wire  _EVAL_30;
  wire [31:0] _EVAL_31;
  wire [31:0] _EVAL_32;
  wire  _EVAL_33;
  wire [31:0] _EVAL_34;
  wire [31:0] _EVAL_35;
  wire [31:0] _EVAL_36;
  wire [3:0] _EVAL_37;
  wire [31:0] MemTap_mem_0;
  wire [31:0] MemTap_mem_1;
  wire [31:0] MemTap_mem_2;
  wire [31:0] MemTap_mem_3;
  wire [31:0] MemTap_mem_4;
  wire [31:0] MemTap_mem_5;
  wire [31:0] MemTap_mem_6;
  wire [31:0] MemTap_mem_7;
  wire [31:0] MemTap_mem_8;
  wire [31:0] MemTap_mem_9;
  wire [31:0] MemTap_mem_10;
  wire [31:0] MemTap_mem_11;
  wire [31:0] MemTap_mem_12;
  wire [31:0] MemTap_mem_13;
  wire [31:0] MemTap_mem_14;
  wire [31:0] MemTap_mem_15;
  wire [31:0] MemTap_mem_16;
  wire [31:0] MemTap_mem_17;
  wire [31:0] MemTap_mem_18;
  wire [31:0] MemTap_mem_19;
  wire [31:0] MemTap_mem_20;
  wire [31:0] MemTap_mem_21;
  wire [31:0] MemTap_mem_22;
  wire [31:0] MemTap_mem_23;
  wire [31:0] MemTap_mem_24;
  wire [31:0] MemTap_mem_25;
  wire [31:0] MemTap_mem_26;
  wire [31:0] MemTap_mem_27;
  wire [31:0] MemTap_mem_28;
  wire [31:0] MemTap_mem_29;
  wire [31:0] MemTap_mem_30;
  wire [3:0] _EVAL_38;
  wire  _EVAL_39;
  wire [1:0] _EVAL_40;
  wire [31:0] _EVAL_41;
  wire [31:0] _EVAL_42;
  wire  _EVAL_43;
  wire [31:0] _EVAL_44;
  wire [31:0] _EVAL_45;
  wire [31:0] _EVAL_46;
  wire [2:0] _EVAL_47;
  wire [2:0] _EVAL_48;
  wire [31:0] _EVAL_49;
  wire [31:0] _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire [31:0] _EVAL_53;
  wire  _EVAL_54;
  wire [31:0] _EVAL_55;
  wire [31:0] _EVAL_56;
  wire [31:0] _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire [3:0] _EVAL_60;
  wire [31:0] _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire [31:0] _EVAL_64;
  wire [3:0] _EVAL_65;
  wire  _EVAL_66;
  wire [31:0] _EVAL_67;
  wire [31:0] _EVAL_68;
  wire [31:0] _EVAL_69;
  wire  _EVAL_70;
  wire [31:0] _EVAL_71;
  wire [3:0] _EVAL_72;
  wire  _EVAL_73;
  wire [31:0] _EVAL_74;
  wire [31:0] _EVAL_75;
  wire [31:0] _EVAL_76;
  wire [2:0] _EVAL_77;
  wire [31:0] _EVAL_78;
  wire [2:0] _EVAL_79;
  wire [3:0] _EVAL_80;
  wire [31:0] _EVAL_81;
  wire [31:0] _EVAL_82;
  wire [31:0] _EVAL_83;
  wire [31:0] _EVAL_84;
  wire [31:0] _EVAL_85;
  wire  DataTap_1_1__5;
  wire [31:0] DataTap_1_1__4;
  wire  DataTap_1_1__3;
  wire  DataTap_1_1__2;
  wire  DataTap_1_1__1;
  wire  DataTap_1_1__0;
  wire  DataTap_1__2;
  wire  DataTap_1__1;
  wire  DataTap_1__0;
  wire [31:0] _EVAL_86;
  wire [31:0] _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire [31:0] _EVAL_91;
  wire [31:0] _EVAL_92;
  wire [31:0] _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire [31:0] _EVAL_96;
  wire [31:0] _EVAL_97;
  wire [31:0] _EVAL_98;
  wire  _EVAL_99;
  wire [31:0] _EVAL_100;
  wire [31:0] _EVAL_101;
  wire  _EVAL_102;
  wire [31:0] _EVAL_103;
  wire  _EVAL_104;
  wire [31:0] _EVAL_105;
  wire  _EVAL_106;
  wire [31:0] _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire [31:0] _EVAL_110;
  wire  _EVAL_111;
  wire [31:0] _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire [31:0] _EVAL_115;
  wire [31:0] _EVAL_116;
  wire  _EVAL_117;
  SiFive_MemTap MemTap (
    .mem_0(MemTap_mem_0),
    .mem_1(MemTap_mem_1),
    .mem_2(MemTap_mem_2),
    .mem_3(MemTap_mem_3),
    .mem_4(MemTap_mem_4),
    .mem_5(MemTap_mem_5),
    .mem_6(MemTap_mem_6),
    .mem_7(MemTap_mem_7),
    .mem_8(MemTap_mem_8),
    .mem_9(MemTap_mem_9),
    .mem_10(MemTap_mem_10),
    .mem_11(MemTap_mem_11),
    .mem_12(MemTap_mem_12),
    .mem_13(MemTap_mem_13),
    .mem_14(MemTap_mem_14),
    .mem_15(MemTap_mem_15),
    .mem_16(MemTap_mem_16),
    .mem_17(MemTap_mem_17),
    .mem_18(MemTap_mem_18),
    .mem_19(MemTap_mem_19),
    .mem_20(MemTap_mem_20),
    .mem_21(MemTap_mem_21),
    .mem_22(MemTap_mem_22),
    .mem_23(MemTap_mem_23),
    .mem_24(MemTap_mem_24),
    .mem_25(MemTap_mem_25),
    .mem_26(MemTap_mem_26),
    .mem_27(MemTap_mem_27),
    .mem_28(MemTap_mem_28),
    .mem_29(MemTap_mem_29),
    .mem_30(MemTap_mem_30)
  );
  SiFive_Insight_hart_0_mapping SiFive_Insight_hart_0_mapping (
  );
  SiFive_DataTap_1_0 DataTap_1_1 (
    ._5(DataTap_1_1__5),
    ._4(DataTap_1_1__4),
    ._3(DataTap_1_1__3),
    ._2(DataTap_1_1__2),
    ._1(DataTap_1_1__1),
    ._0(DataTap_1_1__0)
  );
  SiFive_DataTap_1 DataTap_1 (
    ._2(DataTap_1__2),
    ._1(DataTap_1__1),
    ._0(DataTap_1__0)
  );
  assign _EVAL_46 = _EVAL_75;
  assign _EVAL_3 = 2'h0;
  assign _EVAL_34 = MemTap_mem_5;
  assign _EVAL_59 = 1'h0;
  assign _EVAL_103 = MemTap_mem_22;
  assign _EVAL_57 = MemTap_mem_12;
  assign _EVAL_13 = 1'h0;
  assign _EVAL_44 = 32'h0;
  assign _EVAL_78 = _EVAL_10;
  assign _EVAL_63 = DataTap_1__1;
  assign _EVAL_85 = _EVAL_49;
  assign _EVAL_21 = MemTap_mem_1;
  assign _EVAL = 3'h0;
  assign _EVAL_58 = 1'h0;
  assign _EVAL_117 = _EVAL_102 & _EVAL_63;
  assign _EVAL_4 = MemTap_mem_9;
  assign _EVAL_48 = 3'h0;
  assign _EVAL_18 = 32'h0;
  assign _EVAL_25 = MemTap_mem_21;
  assign _EVAL_84 = _EVAL_96;
  assign _EVAL_15 = _EVAL_20;
  assign _EVAL_33 = ~_EVAL_104;
  assign _EVAL_106 = _EVAL_88 & _EVAL_63;
  assign _EVAL_35 = _EVAL_98;
  assign _EVAL_20 = MemTap_mem_2;
  assign _EVAL_75 = MemTap_mem_24;
  assign _EVAL_65 = 4'h0;
  assign _EVAL_79 = 3'h0;
  assign _EVAL_60 = 4'h0;
  assign _EVAL_105 = 32'h0;
  assign _EVAL_5 = _EVAL_81;
  assign _EVAL_54 = 1'h0;
  assign _EVAL_31 = MemTap_mem_18;
  assign _EVAL_26 = 32'h0;
  assign _EVAL_6 = _EVAL_103;
  assign _EVAL_17 = _EVAL_21;
  assign _EVAL_107 = 32'h0;
  assign _EVAL_8 = 3'h0;
  assign _EVAL_12 = 1'h0;
  assign _EVAL_23 = _EVAL_4;
  assign _EVAL_50 = MemTap_mem_26;
  assign _EVAL_112 = MemTap_mem_16;
  assign _EVAL_108 = 1'h0;
  assign _EVAL_93 = _EVAL_0;
  assign _EVAL_102 = DataTap_1__2;
  assign _EVAL_1 = _EVAL_64;
  assign _EVAL_70 = _EVAL_99 & _EVAL_66;
  assign _EVAL_101 = 32'h0;
  assign _EVAL_68 = _EVAL_34;
  assign _EVAL_116 = _EVAL_67;
  assign _EVAL_27 = ~_EVAL_102;
  assign _EVAL_40 = 2'h0;
  assign _EVAL_52 = 1'h0;
  assign _EVAL_82 = MemTap_mem_3;
  assign _EVAL_29 = MemTap_mem_8;
  assign _EVAL_64 = MemTap_mem_27;
  assign _EVAL_61 = MemTap_mem_23;
  assign _EVAL_83 = _EVAL_19;
  assign _EVAL_0 = MemTap_mem_11;
  assign _EVAL_73 = _EVAL_33 & _EVAL_63;
  assign _EVAL_43 = 1'h0;
  assign _EVAL_99 = DataTap_1_1__3;
  assign _EVAL_80 = 4'h0;
  assign _EVAL_109 = 1'h0;
  assign _EVAL_51 = 1'h0;
  assign _EVAL_71 = _EVAL_31;
  assign _EVAL_95 = 1'h0;
  assign _EVAL_81 = MemTap_mem_14;
  assign _EVAL_16 = MemTap_mem_6;
  assign _EVAL_39 = 1'h0;
  assign _EVAL_86 = _EVAL_45;
  assign _EVAL_22 = _EVAL_16;
  assign _EVAL_36 = _EVAL_97;
  assign _EVAL_98 = MemTap_mem_0;
  assign _EVAL_113 = 1'h0;
  assign _EVAL_47 = 3'h0;
  assign _EVAL_38 = 4'h0;
  assign _EVAL_100 = MemTap_mem_15;
  assign _EVAL_55 = _EVAL_61;
  assign _EVAL_77 = 3'h0;
  assign _EVAL_90 = 1'h0;
  assign _EVAL_115 = _EVAL_9;
  assign _EVAL_89 = 1'h0;
  assign _EVAL_9 = MemTap_mem_13;
  assign _EVAL_41 = _EVAL_57;
  assign _EVAL_24 = 32'h0;
  assign _EVAL_62 = 1'h0;
  assign _EVAL_11 = 1'h0;
  assign _EVAL_66 = DataTap_1_1__5;
  assign _EVAL_28 = _EVAL_82;
  assign _EVAL_30 = 1'h0;
  assign _EVAL_96 = MemTap_mem_4;
  assign _EVAL_69 = _EVAL_25;
  assign _EVAL_19 = MemTap_mem_28;
  assign _EVAL_42 = MemTap_mem_30;
  assign _EVAL_88 = _EVAL_104 & _EVAL_27;
  assign _EVAL_67 = MemTap_mem_17;
  assign _EVAL_72 = 4'h0;
  assign _EVAL_7 = 32'h0;
  assign _EVAL_110 = 32'h0;
  assign _EVAL_94 = 1'h0;
  assign _EVAL_104 = DataTap_1__0;
  assign _EVAL_37 = 4'h0;
  assign _EVAL_10 = MemTap_mem_20;
  assign _EVAL_56 = _EVAL_42;
  assign _EVAL_53 = MemTap_mem_10;
  assign _EVAL_91 = _EVAL_53;
  assign _EVAL_97 = MemTap_mem_7;
  assign _EVAL_32 = _EVAL_112;
  assign _EVAL_76 = _EVAL_100;
  assign _EVAL_74 = _EVAL_29;
  assign _EVAL_111 = 1'h0;
  assign _EVAL_87 = _EVAL_50;
  assign _EVAL_114 = 1'h0;
  assign _EVAL_49 = MemTap_mem_29;
  assign _EVAL_45 = MemTap_mem_25;
  assign _EVAL_2 = MemTap_mem_19;
  assign _EVAL_92 = _EVAL_2;
  assign _EVAL_14 = 1'h0;
endmodule
