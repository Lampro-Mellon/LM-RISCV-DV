//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_182(
  input  [15:0] _EVAL,
  input  [3:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  output        _EVAL_4,
  input  [10:0] _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8
);
  reg  _EVAL_10;
  reg [31:0] _RAND_0;
  wire  _EVAL_12;
  wire  _EVAL_14;
  wire  _EVAL_15;
  reg  _EVAL_16;
  reg [31:0] _RAND_1;
  reg  _EVAL_17;
  reg [31:0] _RAND_2;
  wire  _EVAL_18;
  wire  _EVAL_19;
  reg  _EVAL_20;
  reg [31:0] _RAND_3;
  reg  _EVAL_21;
  reg [31:0] _RAND_4;
  reg  _EVAL_23;
  reg [31:0] _RAND_5;
  reg  _EVAL_25;
  reg [31:0] _RAND_6;
  reg  _EVAL_28;
  reg [31:0] _RAND_7;
  reg  _EVAL_29;
  reg [31:0] _RAND_8;
  reg  _EVAL_33;
  reg [31:0] _RAND_9;
  wire  _EVAL_36;
  wire  _EVAL_37;
  reg  _EVAL_39;
  reg [31:0] _RAND_10;
  wire  _EVAL_42;
  wire  _EVAL_43;
  reg  _EVAL_45;
  reg [31:0] _RAND_11;
  reg  _EVAL_46;
  reg [31:0] _RAND_12;
  reg  _EVAL_49;
  reg [31:0] _RAND_13;
  wire [31:0] _EVAL_53;
  wire  _EVAL_55;
  wire  _EVAL_56;
  reg  _EVAL_58;
  reg [31:0] _RAND_14;
  wire  _EVAL_60;
  wire  _EVAL_62;
  wire  _EVAL_63;
  reg  _EVAL_64;
  reg [31:0] _RAND_15;
  wire  _EVAL_65;
  wire  _EVAL_67;
  reg  _EVAL_68;
  reg [31:0] _RAND_16;
  wire  _EVAL_69;
  reg  _EVAL_73;
  reg [31:0] _RAND_17;
  reg  _EVAL_74;
  reg [31:0] _RAND_18;
  wire  _EVAL_75;
  wire  _EVAL_76;
  reg  _EVAL_77;
  reg [31:0] _RAND_19;
  reg  _EVAL_78;
  reg [31:0] _RAND_20;
  wire  _EVAL_82;
  reg  _EVAL_83;
  reg [31:0] _RAND_21;
  wire  _EVAL_84;
  reg  _EVAL_85;
  reg [31:0] _RAND_22;
  wire  _EVAL_86;
  wire  _EVAL_88;
  reg  _EVAL_91;
  reg [31:0] _RAND_23;
  reg  _EVAL_93;
  reg [31:0] _RAND_24;
  reg  _EVAL_97;
  reg [31:0] _RAND_25;
  reg  _EVAL_98;
  reg [31:0] _RAND_26;
  wire  _EVAL_99;
  reg  _EVAL_100;
  reg [31:0] _RAND_27;
  reg  _EVAL_101;
  reg [31:0] _RAND_28;
  wire  _EVAL_102;
  reg  _EVAL_104;
  reg [31:0] _RAND_29;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_113;
  reg  _EVAL_114;
  reg [31:0] _RAND_30;
  reg  _EVAL_115;
  reg [31:0] _RAND_31;
  wire  _EVAL_116;
  wire  _EVAL_117;
  assign _EVAL_53 = {_EVAL_0,_EVAL,_EVAL_5,1'h1};
  assign _EVAL_18 = _EVAL_53[3];
  assign _EVAL_67 = _EVAL_53[24];
  assign _EVAL_14 = _EVAL_53[13];
  assign _EVAL_69 = _EVAL_53[22];
  assign _EVAL_82 = _EVAL_53[5];
  assign _EVAL_55 = _EVAL_53[23];
  assign _EVAL_102 = _EVAL_53[12];
  assign _EVAL_60 = _EVAL_53[2];
  assign _EVAL_75 = _EVAL_53[21];
  assign _EVAL_42 = _EVAL_53[19];
  assign _EVAL_110 = _EVAL_53[10];
  assign _EVAL_111 = _EVAL_53[28];
  assign _EVAL_116 = _EVAL_53[8];
  assign _EVAL_84 = _EVAL_53[20];
  assign _EVAL_113 = _EVAL_53[18];
  assign _EVAL_117 = _EVAL_53[1];
  assign _EVAL_4 = _EVAL_49;
  assign _EVAL_76 = _EVAL_53[14];
  assign _EVAL_15 = _EVAL_53[6];
  assign _EVAL_12 = _EVAL_53[4];
  assign _EVAL_65 = _EVAL_53[17];
  assign _EVAL_63 = _EVAL_53[31];
  assign _EVAL_37 = _EVAL_53[9];
  assign _EVAL_88 = _EVAL_53[26];
  assign _EVAL_56 = _EVAL_53[15];
  assign _EVAL_43 = _EVAL_53[29];
  assign _EVAL_62 = _EVAL_53[30];
  assign _EVAL_107 = _EVAL_53[27];
  assign _EVAL_86 = _EVAL_53[7];
  assign _EVAL_106 = _EVAL_53[0];
  assign _EVAL_36 = _EVAL_53[11];
  assign _EVAL_19 = _EVAL_53[25];
  assign _EVAL_99 = _EVAL_53[16];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_10 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_16 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_17 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_20 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_21 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_23 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_25 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_28 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_29 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_33 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_39 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_45 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_46 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_49 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_58 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_64 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_68 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_73 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_74 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_77 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_78 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_83 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_85 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_91 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_93 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_97 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_98 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_100 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_101 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_104 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_114 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_115 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_7) begin
    if (_EVAL_6) begin
      _EVAL_10 <= _EVAL_110;
    end else if (_EVAL_3) begin
      _EVAL_10 <= _EVAL_16;
    end
    if (_EVAL_6) begin
      _EVAL_16 <= _EVAL_36;
    end else if (_EVAL_3) begin
      _EVAL_16 <= _EVAL_33;
    end
    if (_EVAL_6) begin
      _EVAL_17 <= _EVAL_107;
    end else if (_EVAL_3) begin
      _EVAL_17 <= _EVAL_20;
    end
    if (_EVAL_6) begin
      _EVAL_20 <= _EVAL_111;
    end else if (_EVAL_3) begin
      _EVAL_20 <= _EVAL_29;
    end
    if (_EVAL_6) begin
      _EVAL_21 <= _EVAL_12;
    end else if (_EVAL_3) begin
      _EVAL_21 <= _EVAL_97;
    end
    if (_EVAL_6) begin
      _EVAL_23 <= _EVAL_63;
    end else if (_EVAL_3) begin
      _EVAL_23 <= _EVAL_2;
    end
    if (_EVAL_6) begin
      _EVAL_25 <= _EVAL_42;
    end else if (_EVAL_3) begin
      _EVAL_25 <= _EVAL_39;
    end
    if (_EVAL_6) begin
      _EVAL_28 <= _EVAL_75;
    end else if (_EVAL_3) begin
      _EVAL_28 <= _EVAL_68;
    end
    if (_EVAL_6) begin
      _EVAL_29 <= _EVAL_43;
    end else if (_EVAL_3) begin
      _EVAL_29 <= _EVAL_85;
    end
    if (_EVAL_6) begin
      _EVAL_33 <= _EVAL_102;
    end else if (_EVAL_3) begin
      _EVAL_33 <= _EVAL_46;
    end
    if (_EVAL_6) begin
      _EVAL_39 <= _EVAL_84;
    end else if (_EVAL_3) begin
      _EVAL_39 <= _EVAL_28;
    end
    if (_EVAL_6) begin
      _EVAL_45 <= _EVAL_15;
    end else if (_EVAL_3) begin
      _EVAL_45 <= _EVAL_77;
    end
    if (_EVAL_6) begin
      _EVAL_46 <= _EVAL_14;
    end else if (_EVAL_3) begin
      _EVAL_46 <= _EVAL_58;
    end
    if (_EVAL_6) begin
      _EVAL_49 <= _EVAL_106;
    end else if (_EVAL_3) begin
      _EVAL_49 <= _EVAL_115;
    end
    if (_EVAL_6) begin
      _EVAL_58 <= _EVAL_76;
    end else if (_EVAL_3) begin
      _EVAL_58 <= _EVAL_114;
    end
    if (_EVAL_6) begin
      _EVAL_64 <= _EVAL_19;
    end else if (_EVAL_3) begin
      _EVAL_64 <= _EVAL_104;
    end
    if (_EVAL_6) begin
      _EVAL_68 <= _EVAL_69;
    end else if (_EVAL_3) begin
      _EVAL_68 <= _EVAL_100;
    end
    if (_EVAL_6) begin
      _EVAL_73 <= _EVAL_18;
    end else if (_EVAL_3) begin
      _EVAL_73 <= _EVAL_21;
    end
    if (_EVAL_6) begin
      _EVAL_74 <= _EVAL_67;
    end else if (_EVAL_3) begin
      _EVAL_74 <= _EVAL_64;
    end
    if (_EVAL_6) begin
      _EVAL_77 <= _EVAL_86;
    end else if (_EVAL_3) begin
      _EVAL_77 <= _EVAL_101;
    end
    if (_EVAL_6) begin
      _EVAL_78 <= _EVAL_60;
    end else if (_EVAL_3) begin
      _EVAL_78 <= _EVAL_73;
    end
    if (_EVAL_6) begin
      _EVAL_83 <= _EVAL_37;
    end else if (_EVAL_3) begin
      _EVAL_83 <= _EVAL_10;
    end
    if (_EVAL_6) begin
      _EVAL_85 <= _EVAL_62;
    end else if (_EVAL_3) begin
      _EVAL_85 <= _EVAL_23;
    end
    if (_EVAL_6) begin
      _EVAL_91 <= _EVAL_99;
    end else if (_EVAL_3) begin
      _EVAL_91 <= _EVAL_98;
    end
    if (_EVAL_6) begin
      _EVAL_93 <= _EVAL_113;
    end else if (_EVAL_3) begin
      _EVAL_93 <= _EVAL_25;
    end
    if (_EVAL_6) begin
      _EVAL_97 <= _EVAL_82;
    end else if (_EVAL_3) begin
      _EVAL_97 <= _EVAL_45;
    end
    if (_EVAL_6) begin
      _EVAL_98 <= _EVAL_65;
    end else if (_EVAL_3) begin
      _EVAL_98 <= _EVAL_93;
    end
    if (_EVAL_6) begin
      _EVAL_100 <= _EVAL_55;
    end else if (_EVAL_3) begin
      _EVAL_100 <= _EVAL_74;
    end
    if (_EVAL_6) begin
      _EVAL_101 <= _EVAL_116;
    end else if (_EVAL_3) begin
      _EVAL_101 <= _EVAL_83;
    end
    if (_EVAL_6) begin
      _EVAL_104 <= _EVAL_88;
    end else if (_EVAL_3) begin
      _EVAL_104 <= _EVAL_17;
    end
    if (_EVAL_6) begin
      _EVAL_114 <= _EVAL_56;
    end else if (_EVAL_3) begin
      _EVAL_114 <= _EVAL_91;
    end
    if (_EVAL_6) begin
      _EVAL_115 <= _EVAL_117;
    end else if (_EVAL_3) begin
      _EVAL_115 <= _EVAL_78;
    end
  end
endmodule
