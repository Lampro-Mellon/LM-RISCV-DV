//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_49(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [31:0] _EVAL_2,
  input  [31:0] _EVAL_3,
  output        _EVAL_4,
  output [3:0]  _EVAL_5,
  input         _EVAL_6,
  output        _EVAL_7,
  output        _EVAL_8,
  input  [1:0]  _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  input  [3:0]  _EVAL_12,
  input  [2:0]  _EVAL_13,
  output        _EVAL_14,
  input         _EVAL_15,
  output        _EVAL_16,
  output        _EVAL_17,
  output [31:0] _EVAL_18,
  input  [31:0] _EVAL_19,
  input         _EVAL_20,
  input         _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  output        _EVAL_25,
  output [31:0] _EVAL_26,
  output        _EVAL_27,
  output        _EVAL_28,
  input  [3:0]  _EVAL_29,
  output        _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_34,
  output        _EVAL_35,
  output [3:0]  _EVAL_36,
  output [2:0]  _EVAL_37,
  input         _EVAL_38,
  input  [3:0]  _EVAL_39,
  output        _EVAL_40,
  output [31:0] _EVAL_41
);
  assign _EVAL_17 = _EVAL;
  assign _EVAL_41 = _EVAL_19;
  assign _EVAL_16 = _EVAL_22;
  assign _EVAL_27 = _EVAL_33;
  assign _EVAL_26 = _EVAL_3;
  assign _EVAL_25 = _EVAL_23;
  assign _EVAL_14 = _EVAL_10;
  assign _EVAL_30 = _EVAL_38;
  assign _EVAL_36 = _EVAL_39;
  assign _EVAL_18 = _EVAL_2;
  assign _EVAL_37 = _EVAL_11;
  assign _EVAL_8 = _EVAL_31;
  assign _EVAL_7 = _EVAL_32;
  assign _EVAL_5 = _EVAL_29;
  assign _EVAL_4 = _EVAL_20;
  assign _EVAL_40 = _EVAL_21;
  assign _EVAL_28 = _EVAL_0;
  assign _EVAL_35 = _EVAL_24;
endmodule
