//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_22(
  input         _EVAL,
  output [31:0] _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [30:0] _EVAL_2,
  input         _EVAL_3,
  output        _EVAL_4,
  output [31:0] _EVAL_5,
  output [1:0]  _EVAL_6,
  output        _EVAL_7,
  output        _EVAL_8,
  input  [3:0]  _EVAL_9,
  output [1:0]  _EVAL_10,
  output [30:0] _EVAL_11,
  output [2:0]  _EVAL_12,
  input         _EVAL_13,
  input  [2:0]  _EVAL_14,
  output        _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19,
  input  [2:0]  _EVAL_20,
  output [2:0]  _EVAL_21,
  input         _EVAL_22,
  output        _EVAL_23,
  input         _EVAL_24,
  output [2:0]  _EVAL_25,
  input  [31:0] _EVAL_26,
  output [3:0]  _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  output [2:0]  _EVAL_30,
  input  [2:0]  _EVAL_31,
  output [2:0]  _EVAL_32,
  input  [31:0] _EVAL_33,
  input         _EVAL_34
);
  wire  _EVAL_35;
  wire  _EVAL_36;
  reg [2:0] _EVAL_37;
  reg [31:0] _RAND_0;
  reg  _EVAL_38;
  reg [31:0] _RAND_1;
  wire [30:0] _EVAL_39;
  reg [2:0] _EVAL_40;
  reg [31:0] _RAND_2;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire [30:0] _EVAL_43;
  wire [2:0] _EVAL_44;
  wire [30:0] _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire [3:0] _EVAL_49;
  wire [2:0] _EVAL_50;
  wire [2:0] _EVAL_53;
  wire [3:0] _EVAL_54;
  wire [2:0] Queue__EVAL;
  wire  Queue__EVAL_0;
  wire  Queue__EVAL_1;
  wire  Queue__EVAL_2;
  wire [1:0] Queue__EVAL_3;
  wire  Queue__EVAL_4;
  wire  Queue__EVAL_5;
  wire [2:0] Queue__EVAL_6;
  wire  Queue__EVAL_7;
  wire  Queue__EVAL_8;
  wire  Queue__EVAL_9;
  wire [2:0] Queue__EVAL_10;
  wire [2:0] Queue__EVAL_11;
  wire [2:0] Queue__EVAL_12;
  wire [31:0] Queue__EVAL_13;
  wire  Queue__EVAL_14;
  wire  Queue__EVAL_15;
  wire  Queue__EVAL_16;
  wire [2:0] Queue__EVAL_17;
  wire [31:0] Queue__EVAL_18;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  reg [2:0] _EVAL_60;
  reg [31:0] _RAND_3;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire [1:0] _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire [6:0] _EVAL_68;
  wire [3:0] _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire [5:0] _EVAL_74;
  wire  _EVAL_75;
  reg  _EVAL_76;
  reg [31:0] _RAND_4;
  wire [3:0] _EVAL_77;
  wire [30:0] _EVAL_78;
  wire [5:0] _EVAL_80;
  reg  _EVAL_81;
  reg [31:0] _RAND_5;
  wire [1:0] _EVAL_82;
  wire [2:0] _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_86;
  reg  _EVAL_88;
  reg [31:0] _RAND_6;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  reg [2:0] _EVAL_92;
  reg [31:0] _RAND_7;
  reg  _EVAL_93;
  reg [31:0] _RAND_8;
  wire  _EVAL_95;
  wire  _EVAL_96;
  reg  _EVAL_97;
  reg [31:0] _RAND_9;
  wire  _EVAL_98;
  wire [30:0] _EVAL_99;
  reg  _EVAL_100;
  reg [31:0] _RAND_10;
  wire  _EVAL_101;
  wire  _EVAL_102;
  reg  _EVAL_103;
  reg [31:0] _RAND_11;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  reg [31:0] _EVAL_107;
  reg [31:0] _RAND_12;
  wire [5:0] _EVAL_108;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire [2:0] _EVAL_120;
  wire  _EVAL_121;
  wire [1:0] _EVAL_122;
  wire  _EVAL_123;
  reg  _EVAL_124;
  reg [31:0] _RAND_13;
  wire [4:0] _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire [2:0] _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_131;
  wire [24:0] _EVAL_133;
  wire [1:0] _EVAL_134;
  wire [5:0] _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  reg [30:0] _EVAL_141;
  reg [31:0] _RAND_14;
  wire  _EVAL_143;
  wire [1:0] _EVAL_146;
  wire [3:0] _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  reg [31:0] _EVAL_152;
  reg [31:0] _RAND_15;
  wire [2:0] _EVAL_153;
  wire [12:0] _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire [1:0] _EVAL_161;
  wire  _EVAL_162;
  wire [3:0] _EVAL_163;
  wire [30:0] _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire [30:0] _EVAL_168;
  reg [2:0] _EVAL_170;
  reg [31:0] _RAND_16;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire [1:0] _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire [1:0] _EVAL_179;
  wire [3:0] _EVAL_180;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  reg  _EVAL_187;
  reg [31:0] _RAND_17;
  reg  _EVAL_188;
  reg [31:0] _RAND_18;
  wire [2:0] _EVAL_189;
  reg  _EVAL_190;
  reg [31:0] _RAND_19;
  wire  _EVAL_191;
  wire [1:0] _EVAL_192;
  wire [2:0] _EVAL_193;
  wire  _EVAL_194;
  wire [3:0] _EVAL_195;
  wire  _EVAL_196;
  wire [27:0] _EVAL_198;
  reg [2:0] _EVAL_199;
  reg [31:0] _RAND_20;
  wire [2:0] _EVAL_200;
  wire  _EVAL_201;
  reg  _EVAL_202;
  reg [31:0] _RAND_21;
  reg  _EVAL_203;
  reg [31:0] _RAND_22;
  wire  _EVAL_204;
  wire  _EVAL_205;
  reg [1:0] _EVAL_206;
  reg [31:0] _RAND_23;
  wire  _EVAL_207;
  wire  _EVAL_208;
  _EVAL_21 Queue (
    ._EVAL(Queue__EVAL),
    ._EVAL_0(Queue__EVAL_0),
    ._EVAL_1(Queue__EVAL_1),
    ._EVAL_2(Queue__EVAL_2),
    ._EVAL_3(Queue__EVAL_3),
    ._EVAL_4(Queue__EVAL_4),
    ._EVAL_5(Queue__EVAL_5),
    ._EVAL_6(Queue__EVAL_6),
    ._EVAL_7(Queue__EVAL_7),
    ._EVAL_8(Queue__EVAL_8),
    ._EVAL_9(Queue__EVAL_9),
    ._EVAL_10(Queue__EVAL_10),
    ._EVAL_11(Queue__EVAL_11),
    ._EVAL_12(Queue__EVAL_12),
    ._EVAL_13(Queue__EVAL_13),
    ._EVAL_14(Queue__EVAL_14),
    ._EVAL_15(Queue__EVAL_15),
    ._EVAL_16(Queue__EVAL_16),
    ._EVAL_17(Queue__EVAL_17),
    ._EVAL_18(Queue__EVAL_18)
  );
  assign _EVAL_151 = _EVAL_93 ? _EVAL_70 : _EVAL_205;
  assign _EVAL_64 = _EVAL_38 ? 2'h0 : 2'h1;
  assign _EVAL_110 = _EVAL_97 ? _EVAL_88 : _EVAL_102;
  assign _EVAL_177 = ~_EVAL_110;
  assign _EVAL_165 = _EVAL_176 | _EVAL_113;
  assign _EVAL_0 = Queue__EVAL_18;
  assign _EVAL_70 = _EVAL_185 & _EVAL_143;
  assign _EVAL_82 = {{1'd0}, _EVAL_166};
  assign _EVAL_83 = _EVAL_205 ? _EVAL_31 : _EVAL_40;
  assign _EVAL_149 = _EVAL_97 ? 1'h0 : _EVAL_151;
  assign _EVAL_7 = Queue__EVAL_16;
  assign _EVAL_72 = _EVAL_93 ? _EVAL_81 : _EVAL_150;
  assign _EVAL_78 = _EVAL_93 ? _EVAL_141 : _EVAL_99;
  assign _EVAL_143 = ~_EVAL_202;
  assign _EVAL_205 = _EVAL_116 & _EVAL_16;
  assign _EVAL_128 = _EVAL_97 ? _EVAL_40 : _EVAL_53;
  assign _EVAL_99 = _EVAL_160 ? _EVAL_2 : _EVAL_141;
  assign _EVAL_175 = {_EVAL_35,_EVAL_86};
  assign _EVAL_127 = _EVAL_95 | _EVAL_203;
  assign _EVAL_10 = Queue__EVAL_3;
  assign Queue__EVAL = _EVAL_37;
  assign _EVAL_207 = _EVAL_205 | _EVAL_93;
  assign _EVAL_171 = _EVAL_93 ? _EVAL_204 : _EVAL_129;
  assign _EVAL_47 = ~_EVAL_157;
  assign _EVAL_113 = _EVAL_162 | _EVAL_115;
  assign _EVAL_184 = _EVAL_160 ? _EVAL_47 : _EVAL_202;
  assign _EVAL_183 = _EVAL_97 ? _EVAL_76 : _EVAL_75;
  assign _EVAL_18 = _EVAL_97 ? _EVAL_202 : _EVAL_48;
  assign _EVAL_122 = _EVAL_200[1:0];
  assign _EVAL_176 = _EVAL_111 & _EVAL_73;
  assign _EVAL_95 = ~_EVAL_190;
  assign _EVAL_25 = _EVAL_97 ? _EVAL_199 : _EVAL_189;
  assign _EVAL_148 = {_EVAL_44, 1'h0};
  assign _EVAL_138 = _EVAL_97 ? _EVAL_187 : _EVAL_57;
  assign _EVAL_53 = _EVAL_93 ? _EVAL_40 : _EVAL_83;
  assign _EVAL_136 = _EVAL_68[5:0];
  assign _EVAL_46 = {{25'd0}, _EVAL_74};
  assign _EVAL_126 = _EVAL_97 ? _EVAL_202 : _EVAL_48;
  assign _EVAL_164 = ~_EVAL_168;
  assign _EVAL_35 = _EVAL_97 ? _EVAL_103 : _EVAL_90;
  assign _EVAL_116 = _EVAL_97 ? 1'h0 : _EVAL_101;
  assign _EVAL_68 = _EVAL_80 + 6'h4;
  assign _EVAL_112 = _EVAL_205 ? _EVAL_19 : _EVAL_103;
  assign _EVAL_119 = _EVAL_205 ? _EVAL_13 : _EVAL_188;
  assign _EVAL_198 = _EVAL_39[30:3];
  assign _EVAL_159 = Queue__EVAL_7;
  assign _EVAL_191 = _EVAL_205 ? _EVAL_123 : _EVAL_88;
  assign Queue__EVAL_0 = _EVAL_29;
  assign _EVAL_6 = _EVAL_91 ? _EVAL_134 : _EVAL_64;
  assign _EVAL_163 = _EVAL_97 ? {{1'd0}, _EVAL_60} : _EVAL_195;
  assign _EVAL_27 = {_EVAL_161,_EVAL_175};
  assign _EVAL_115 = _EVAL_62 & _EVAL_177;
  assign _EVAL_65 = _EVAL | _EVAL_121;
  assign _EVAL_192 = _EVAL_203 ? 2'h2 : {{1'd0}, _EVAL_158};
  assign _EVAL_75 = _EVAL_93 ? _EVAL_76 : _EVAL_118;
  assign _EVAL_44 = _EVAL_180[2:0];
  assign _EVAL_80 = _EVAL_168[5:0];
  assign _EVAL_153 = _EVAL_123 ? _EVAL_31 : 3'h2;
  assign _EVAL_160 = _EVAL_205 & _EVAL_98;
  assign _EVAL_21 = Queue__EVAL_12;
  assign _EVAL_168 = _EVAL_97 ? _EVAL_141 : _EVAL_78;
  assign _EVAL_54 = _EVAL_123 ? 4'h0 : _EVAL_69;
  assign _EVAL_180 = _EVAL_125[3:0];
  assign _EVAL_36 = ~_EVAL_104;
  assign _EVAL_118 = _EVAL_205 ? _EVAL_22 : _EVAL_76;
  assign _EVAL_11 = _EVAL_97 ? _EVAL_141 : _EVAL_78;
  assign _EVAL_57 = _EVAL_93 ? _EVAL_187 : _EVAL_105;
  assign _EVAL_158 = _EVAL_124 ? 1'h0 : 1'h1;
  assign _EVAL_155 = 13'h3f << _EVAL_128;
  assign _EVAL_195 = _EVAL_93 ? {{1'd0}, _EVAL_60} : _EVAL_77;
  assign _EVAL_161 = {_EVAL_186,_EVAL_183};
  assign _EVAL_8 = Queue__EVAL_14;
  assign Queue__EVAL_13 = _EVAL_33;
  assign _EVAL_42 = _EVAL_93 ? _EVAL_188 : _EVAL_119;
  assign _EVAL_178 = _EVAL_115 ? 1'h0 : 1'h1;
  assign _EVAL_139 = _EVAL_176 ? _EVAL_38 : _EVAL_58;
  assign _EVAL_73 = ~_EVAL_65;
  assign Queue__EVAL_15 = _EVAL_56 & _EVAL_167;
  assign _EVAL_96 = _EVAL_114 & _EVAL_65;
  assign _EVAL_121 = _EVAL_104 & _EVAL_127;
  assign _EVAL_137 = _EVAL_20 == 3'h5;
  assign _EVAL_89 = _EVAL_198 != 28'h0;
  assign _EVAL_4 = Queue__EVAL_2;
  assign _EVAL_193 = _EVAL_163[2:0];
  assign _EVAL_102 = _EVAL_93 ? _EVAL_88 : _EVAL_191;
  assign _EVAL_125 = _EVAL_49 - 4'h3;
  assign _EVAL_56 = _EVAL_140 & _EVAL_124;
  assign _EVAL_77 = _EVAL_160 ? _EVAL_54 : {{1'd0}, _EVAL_60};
  assign _EVAL_15 = Queue__EVAL_7;
  assign _EVAL_134 = _EVAL_38 ? 2'h2 : 2'h3;
  assign _EVAL_111 = _EVAL_97 ? _EVAL_97 : _EVAL_171;
  assign _EVAL_104 = _EVAL_97 ? _EVAL_81 : _EVAL_72;
  assign _EVAL_49 = {1'h0,_EVAL_31};
  assign _EVAL_189 = _EVAL_93 ? _EVAL_199 : _EVAL_120;
  assign _EVAL_131 = _EVAL_3 & _EVAL_84;
  assign Queue__EVAL_1 = _EVAL_190 & _EVAL_63;
  assign _EVAL_66 = _EVAL_65 & _EVAL_111;
  assign _EVAL_108 = _EVAL_155[5:0];
  assign _EVAL_91 = _EVAL_111 & _EVAL_36;
  assign _EVAL_120 = _EVAL_160 ? _EVAL_153 : _EVAL_199;
  assign _EVAL_61 = _EVAL_206 >= 2'h2;
  assign _EVAL_32 = Queue__EVAL_10;
  assign _EVAL_30 = Queue__EVAL_11;
  assign Queue__EVAL_17 = {{1'd0}, _EVAL_192};
  assign _EVAL_63 = _EVAL | _EVAL_203;
  assign _EVAL_133 = _EVAL_168[30:6];
  assign _EVAL_129 = _EVAL_205 | _EVAL_97;
  assign _EVAL_69 = _EVAL_148 | 4'h1;
  assign _EVAL_162 = _EVAL_62 & _EVAL_201;
  assign _EVAL_98 = ~_EVAL_137;
  assign _EVAL_166 = _EVAL_24 & _EVAL_159;
  assign _EVAL_39 = _EVAL_46 & _EVAL_164;
  assign Queue__EVAL_6 = _EVAL_92;
  assign _EVAL_114 = _EVAL_111 & _EVAL_41;
  assign Queue__EVAL_4 = _EVAL_24;
  assign _EVAL_179 = _EVAL_50[1:0];
  assign _EVAL_208 = ~_EVAL_126;
  assign _EVAL_150 = _EVAL_205 ? _EVAL_137 : _EVAL_81;
  assign Queue__EVAL_9 = _EVAL_17;
  assign _EVAL_86 = ~_EVAL_138;
  assign _EVAL_58 = _EVAL_162 ? _EVAL_38 : _EVAL_178;
  assign _EVAL_194 = _EVAL_185 & _EVAL_202;
  assign _EVAL_43 = {_EVAL_133,_EVAL_136};
  assign _EVAL_172 = ~_EVAL_89;
  assign _EVAL_84 = ~_EVAL_124;
  assign _EVAL_106 = _EVAL_143 | _EVAL_16;
  assign _EVAL_90 = _EVAL_93 ? _EVAL_103 : _EVAL_112;
  assign _EVAL_204 = _EVAL_185 & _EVAL_106;
  assign _EVAL_23 = _EVAL_97 ? 1'h0 : _EVAL_101;
  assign _EVAL_157 = _EVAL_20[2];
  assign _EVAL_156 = _EVAL_180[3];
  assign _EVAL_186 = _EVAL_97 ? _EVAL_188 : _EVAL_42;
  assign _EVAL_101 = _EVAL_93 ? _EVAL_194 : _EVAL_185;
  assign _EVAL_123 = _EVAL_137 | _EVAL_156;
  assign _EVAL_167 = ~_EVAL_203;
  assign _EVAL_74 = ~_EVAL_108;
  assign _EVAL_5 = _EVAL_152;
  assign _EVAL_12 = _EVAL_163[2:0];
  assign _EVAL_41 = _EVAL_110 | _EVAL_208;
  assign _EVAL_50 = _EVAL_206 + _EVAL_146;
  assign _EVAL_62 = _EVAL_97 ? _EVAL_93 : _EVAL_196;
  assign _EVAL_105 = _EVAL_205 ? _EVAL_28 : _EVAL_187;
  assign _EVAL_146 = {{1'd0}, _EVAL_149};
  assign _EVAL_48 = _EVAL_93 ? _EVAL_202 : _EVAL_184;
  assign _EVAL_185 = ~_EVAL_61;
  assign Queue__EVAL_8 = _EVAL_131 & _EVAL_167;
  assign _EVAL_201 = ~_EVAL_111;
  assign _EVAL_140 = _EVAL_3 | _EVAL_100;
  assign _EVAL_196 = _EVAL_93 ? _EVAL_93 : _EVAL_207;
  assign _EVAL_200 = _EVAL_179 - _EVAL_82;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_37 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_38 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_40 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_60 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_76 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_81 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_88 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_92 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_93 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_97 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_100 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_103 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_107 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_124 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_141 = _RAND_14[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_152 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_170 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_187 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_188 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_190 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_199 = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_202 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_203 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_206 = _RAND_23[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_17) begin
    if (_EVAL_66) begin
      if (_EVAL_97) begin
        _EVAL_37 <= _EVAL_170;
      end else if (_EVAL_93) begin
        _EVAL_37 <= _EVAL_170;
      end else if (_EVAL_205) begin
        _EVAL_37 <= _EVAL_14;
      end else begin
        _EVAL_37 <= _EVAL_170;
      end
    end
    _EVAL_38 <= _EVAL_29 | _EVAL_139;
    if (!(_EVAL_97)) begin
      if (!(_EVAL_93)) begin
        if (_EVAL_205) begin
          _EVAL_40 <= _EVAL_31;
        end
      end
    end
    if (_EVAL_29) begin
      _EVAL_60 <= 3'h0;
    end else begin
      _EVAL_60 <= _EVAL_193;
    end
    if (!(_EVAL_97)) begin
      if (!(_EVAL_93)) begin
        if (_EVAL_205) begin
          _EVAL_76 <= _EVAL_22;
        end
      end
    end
    if (!(_EVAL_97)) begin
      if (!(_EVAL_93)) begin
        if (_EVAL_205) begin
          _EVAL_81 <= _EVAL_137;
        end
      end
    end
    if (_EVAL_176) begin
      if (!(_EVAL_97)) begin
        if (!(_EVAL_93)) begin
          if (_EVAL_205) begin
            _EVAL_88 <= _EVAL_123;
          end
        end
      end
    end else if (_EVAL_162) begin
      if (!(_EVAL_97)) begin
        if (!(_EVAL_93)) begin
          if (_EVAL_205) begin
            _EVAL_88 <= _EVAL_123;
          end
        end
      end
    end else if (_EVAL_115) begin
      _EVAL_88 <= _EVAL_172;
    end else if (!(_EVAL_97)) begin
      if (!(_EVAL_93)) begin
        if (_EVAL_205) begin
          _EVAL_88 <= _EVAL_123;
        end
      end
    end
    if (_EVAL_66) begin
      if (_EVAL_97) begin
        _EVAL_92 <= _EVAL_40;
      end else if (_EVAL_93) begin
        _EVAL_92 <= _EVAL_40;
      end else if (_EVAL_205) begin
        _EVAL_92 <= _EVAL_31;
      end else begin
        _EVAL_92 <= _EVAL_40;
      end
    end
    if (_EVAL_29) begin
      _EVAL_93 <= 1'h0;
    end else begin
      _EVAL_93 <= _EVAL_165;
    end
    if (_EVAL_29) begin
      _EVAL_97 <= 1'h0;
    end else begin
      _EVAL_97 <= _EVAL_176;
    end
    if (_EVAL_63) begin
      if (_EVAL_38) begin
        _EVAL_100 <= 1'h0;
      end else begin
        _EVAL_100 <= _EVAL_140;
      end
    end
    if (!(_EVAL_97)) begin
      if (!(_EVAL_93)) begin
        if (_EVAL_205) begin
          _EVAL_103 <= _EVAL_19;
        end
      end
    end
    if (!(_EVAL_97)) begin
      if (_EVAL_93) begin
        _EVAL_107 <= _EVAL_26;
      end else if (_EVAL_160) begin
        _EVAL_107 <= _EVAL_26;
      end
    end
    if (_EVAL_66) begin
      if (_EVAL_97) begin
        _EVAL_124 <= _EVAL_202;
      end else if (_EVAL_93) begin
        _EVAL_124 <= _EVAL_202;
      end else if (_EVAL_160) begin
        _EVAL_124 <= _EVAL_47;
      end else begin
        _EVAL_124 <= _EVAL_202;
      end
    end
    if (_EVAL_29) begin
      _EVAL_141 <= 31'h0;
    end else if (_EVAL_176) begin
      if (!(_EVAL_97)) begin
        if (!(_EVAL_93)) begin
          if (_EVAL_160) begin
            _EVAL_141 <= _EVAL_2;
          end
        end
      end
    end else if (_EVAL_162) begin
      if (!(_EVAL_97)) begin
        if (!(_EVAL_93)) begin
          if (_EVAL_160) begin
            _EVAL_141 <= _EVAL_2;
          end
        end
      end
    end else if (_EVAL_115) begin
      _EVAL_141 <= _EVAL_43;
    end else if (!(_EVAL_97)) begin
      if (!(_EVAL_93)) begin
        if (_EVAL_160) begin
          _EVAL_141 <= _EVAL_2;
        end
      end
    end
    if (_EVAL_65) begin
      if (_EVAL_97) begin
        _EVAL_152 <= _EVAL_107;
      end else if (_EVAL_93) begin
        _EVAL_152 <= _EVAL_26;
      end else if (_EVAL_160) begin
        _EVAL_152 <= _EVAL_26;
      end else begin
        _EVAL_152 <= _EVAL_107;
      end
    end
    if (!(_EVAL_97)) begin
      if (!(_EVAL_93)) begin
        if (_EVAL_205) begin
          _EVAL_170 <= _EVAL_14;
        end
      end
    end
    if (!(_EVAL_97)) begin
      if (!(_EVAL_93)) begin
        if (_EVAL_205) begin
          _EVAL_187 <= _EVAL_28;
        end
      end
    end
    if (!(_EVAL_97)) begin
      if (!(_EVAL_93)) begin
        if (_EVAL_205) begin
          _EVAL_188 <= _EVAL_13;
        end
      end
    end
    if (_EVAL_29) begin
      _EVAL_190 <= 1'h0;
    end else if (_EVAL_63) begin
      _EVAL_190 <= _EVAL_96;
    end
    if (_EVAL_29) begin
      _EVAL_199 <= 3'h0;
    end else if (!(_EVAL_97)) begin
      if (!(_EVAL_93)) begin
        if (_EVAL_160) begin
          if (_EVAL_123) begin
            _EVAL_199 <= _EVAL_31;
          end else begin
            _EVAL_199 <= 3'h2;
          end
        end
      end
    end
    if (!(_EVAL_97)) begin
      if (!(_EVAL_93)) begin
        if (_EVAL_160) begin
          _EVAL_202 <= _EVAL_47;
        end
      end
    end
    if (_EVAL_66) begin
      if (_EVAL_97) begin
        _EVAL_203 <= _EVAL_81;
      end else if (_EVAL_93) begin
        _EVAL_203 <= _EVAL_81;
      end else if (_EVAL_205) begin
        _EVAL_203 <= _EVAL_137;
      end else begin
        _EVAL_203 <= _EVAL_81;
      end
    end
    if (_EVAL_29) begin
      _EVAL_206 <= 2'h0;
    end else begin
      _EVAL_206 <= _EVAL_122;
    end
  end
endmodule
