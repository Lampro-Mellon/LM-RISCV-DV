//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_90_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [1:0]  _EVAL_2,
  input  [1:0]  _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input  [1:0]  _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [3:0]  _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input  [29:0] _EVAL_16,
  input  [2:0]  _EVAL_17,
  input  [2:0]  _EVAL_18
);
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire [1:0] _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  reg [2:0] _EVAL_26;
  reg [31:0] _RAND_0;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  reg  _EVAL_34;
  reg [31:0] _RAND_1;
  wire [7:0] _EVAL_35;
  wire [4:0] _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire [1:0] _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  reg [29:0] _EVAL_50;
  reg [31:0] _RAND_2;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire [1:0] _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  reg [1:0] _EVAL_64;
  reg [31:0] _RAND_3;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire [3:0] _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire [7:0] _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire [31:0] _EVAL_86;
  reg [2:0] _EVAL_87;
  reg [31:0] _RAND_4;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire [30:0] _EVAL_96;
  wire  _EVAL_97;
  wire [1:0] _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  reg  _EVAL_102;
  reg [31:0] _RAND_5;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire [1:0] _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_111;
  wire [3:0] _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire [30:0] _EVAL_123;
  wire  _EVAL_124;
  reg  _EVAL_125;
  reg [31:0] _RAND_6;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire [32:0] _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  reg [2:0] _EVAL_139;
  reg [31:0] _RAND_7;
  wire [4:0] _EVAL_140;
  wire  _EVAL_141;
  wire [1:0] _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  reg  _EVAL_149;
  reg [31:0] _RAND_8;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  reg [2:0] _EVAL_155;
  reg [31:0] _RAND_9;
  wire  _EVAL_157;
  wire [4:0] _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire [29:0] _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire [4:0] _EVAL_177;
  reg  _EVAL_178;
  reg [31:0] _RAND_10;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  reg  _EVAL_184;
  reg [31:0] _RAND_11;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire [4:0] _EVAL_191;
  wire [3:0] _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire [29:0] _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire [3:0] _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  reg [1:0] _EVAL_210;
  reg [31:0] _RAND_12;
  wire [1:0] _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  reg [31:0] _EVAL_218;
  reg [31:0] _RAND_13;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire [29:0] _EVAL_222;
  wire  _EVAL_223;
  wire [1:0] _EVAL_224;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire [1:0] _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire [1:0] _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire [7:0] _EVAL_242;
  wire [7:0] _EVAL_243;
  wire  _EVAL_244;
  reg [1:0] _EVAL_245;
  reg [31:0] _RAND_14;
  wire  _EVAL_246;
  wire  _EVAL_247;
  reg [2:0] _EVAL_248;
  reg [31:0] _RAND_15;
  wire  _EVAL_249;
  wire [4:0] _EVAL_250;
  wire  _EVAL_251;
  wire [4:0] _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_255;
  wire [4:0] _EVAL_256;
  wire  _EVAL_257;
  wire [30:0] _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire [4:0] _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  reg [4:0] _EVAL_271;
  reg [31:0] _RAND_16;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_284;
  wire  _EVAL_285;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_206 = _EVAL_239 | _EVAL_124;
  assign _EVAL_222 = _EVAL_16 & _EVAL_203;
  assign _EVAL_131 = ~_EVAL_104;
  assign _EVAL_109 = _EVAL_5 == _EVAL_139;
  assign _EVAL_200 = _EVAL_12 == 3'h5;
  assign _EVAL_71 = ~_EVAL_273;
  assign _EVAL_224 = 2'h1 << _EVAL_169;
  assign _EVAL_108 = _EVAL_279 | _EVAL_10;
  assign _EVAL_183 = ~_EVAL_102;
  assign _EVAL_151 = _EVAL_18 <= 3'h4;
  assign _EVAL_38 = ~_EVAL_32;
  assign _EVAL_268 = ~_EVAL_231;
  assign _EVAL_282 = _EVAL_216 & _EVAL_182;
  assign _EVAL_143 = _EVAL_6 == _EVAL_64;
  assign _EVAL_247 = _EVAL_16 == _EVAL_50;
  assign _EVAL_214 = ~_EVAL_269;
  assign _EVAL_20 = ~_EVAL_126;
  assign _EVAL_40 = _EVAL_25 | _EVAL_45;
  assign _EVAL_78 = _EVAL_157 & _EVAL_282;
  assign _EVAL_104 = _EVAL_88 | _EVAL_10;
  assign _EVAL_177 = _EVAL_256 & _EVAL_36;
  assign _EVAL_29 = ~_EVAL_63;
  assign _EVAL_123 = $signed(_EVAL_259) & -31'sh2000;
  assign _EVAL_238 = _EVAL_11 == _EVAL_184;
  assign _EVAL_256 = _EVAL_271 | _EVAL_252;
  assign _EVAL_174 = _EVAL_116 | _EVAL_277;
  assign _EVAL_170 = _EVAL_206 | _EVAL_190;
  assign _EVAL_164 = _EVAL_31 | _EVAL_10;
  assign _EVAL_274 = _EVAL_7 == _EVAL_248;
  assign _EVAL_171 = _EVAL_114 | _EVAL_29;
  assign _EVAL_185 = _EVAL_130 | _EVAL_181;
  assign _EVAL_72 = _EVAL_151 | _EVAL_10;
  assign _EVAL_275 = _EVAL_202 | _EVAL_10;
  assign _EVAL_32 = _EVAL_247 | _EVAL_10;
  assign _EVAL_199 = ~_EVAL_236;
  assign _EVAL_122 = ~_EVAL_14;
  assign _EVAL_162 = _EVAL_116 | _EVAL_249;
  assign _EVAL_49 = _EVAL_9 & _EVAL_15;
  assign _EVAL_23 = _EVAL_7[2:1];
  assign _EVAL_63 = _EVAL_252 != 5'h0;
  assign _EVAL_261 = _EVAL_17 == 3'h5;
  assign _EVAL_265 = _EVAL_195 | _EVAL_10;
  assign _EVAL_58 = ~_EVAL_57;
  assign _EVAL_257 = _EVAL_107[0];
  assign _EVAL_43 = ~_EVAL_260;
  assign _EVAL_83 = _EVAL_266 | _EVAL_163;
  assign _EVAL_198 = _EVAL_175 | _EVAL_10;
  assign _EVAL_281 = _EVAL_12 == 3'h4;
  assign _EVAL_119 = _EVAL_2 >= 2'h2;
  assign _EVAL_285 = _EVAL_15 & _EVAL_59;
  assign _EVAL_213 = _EVAL_127 & _EVAL_182;
  assign _EVAL_215 = _EVAL_103 | _EVAL_10;
  assign _EVAL_67 = ~_EVAL_207;
  assign _EVAL_101 = _EVAL_4 & _EVAL_76;
  assign _EVAL_226 = ~_EVAL_178;
  assign _EVAL_33 = _EVAL_172 | _EVAL_10;
  assign _EVAL_128 = _EVAL_15 & _EVAL_138;
  assign _EVAL_53 = _EVAL_127 & _EVAL_217;
  assign _EVAL_107 = _EVAL_34 - 1'h1;
  assign _EVAL_231 = _EVAL_220 | _EVAL_10;
  assign _EVAL_74 = _EVAL_4 & _EVAL_137;
  assign _EVAL_194 = _EVAL_49 & _EVAL_253;
  assign _EVAL_189 = _EVAL_185 | _EVAL_10;
  assign _EVAL_175 = _EVAL_6 != 2'h2;
  assign _EVAL_85 = _EVAL_165 | _EVAL_10;
  assign _EVAL_239 = _EVAL_23 == 2'h1;
  assign _EVAL_284 = _EVAL_56 | _EVAL_10;
  assign _EVAL_150 = _EVAL_17 == 3'h2;
  assign _EVAL_36 = ~_EVAL_250;
  assign _EVAL_229 = _EVAL_171 | _EVAL_10;
  assign _EVAL_188 = _EVAL_66 | _EVAL_10;
  assign _EVAL_241 = ~_EVAL_70;
  assign _EVAL_242 = _EVAL_91 ? _EVAL_243 : 8'h0;
  assign _EVAL_272 = ~_EVAL_105;
  assign _EVAL_180 = _EVAL_15 & _EVAL_261;
  assign _EVAL_90 = ~_EVAL_215;
  assign _EVAL_59 = _EVAL_17 == 3'h1;
  assign _EVAL_140 = _EVAL_252 | _EVAL_271;
  assign _EVAL_209 = _EVAL_228 == 2'h1;
  assign _EVAL_260 = ~_EVAL_34;
  assign _EVAL_179 = _EVAL_17 == 3'h0;
  assign _EVAL_280 = _EVAL_221 | _EVAL_10;
  assign _EVAL_145 = ~_EVAL_108;
  assign _EVAL_44 = _EVAL_95 | _EVAL_10;
  assign _EVAL_230 = ~_EVAL_164;
  assign _EVAL_159 = _EVAL_49 & _EVAL_260;
  assign _EVAL_132 = _EVAL_152 | _EVAL_10;
  assign _EVAL_51 = _EVAL_18 != 3'h0;
  assign _EVAL_130 = _EVAL_209 | _EVAL_99;
  assign _EVAL_54 = _EVAL_106 | _EVAL_49;
  assign _EVAL_117 = _EVAL_94 | _EVAL_10;
  assign _EVAL_65 = _EVAL_271 != 5'h0;
  assign _EVAL_98 = _EVAL_102 - 1'h1;
  assign _EVAL_41 = _EVAL_55 | _EVAL_10;
  assign _EVAL_137 = ~_EVAL_183;
  assign _EVAL_81 = ~_EVAL_237;
  assign _EVAL_278 = _EVAL_40 | _EVAL_92;
  assign _EVAL_28 = _EVAL_4 & _EVAL_46;
  assign _EVAL_141 = _EVAL_4 & _EVAL_244;
  assign _EVAL_227 = ~_EVAL_132;
  assign _EVAL_138 = _EVAL_17 == 3'h4;
  assign _EVAL_186 = _EVAL_240 | _EVAL_10;
  assign _EVAL_47 = _EVAL_15 & _EVAL_264;
  assign _EVAL_133 = _EVAL_218 + 32'h1;
  assign _EVAL_115 = ~_EVAL_284;
  assign _EVAL_95 = _EVAL_18 == 3'h0;
  assign _EVAL_76 = _EVAL_12 == 3'h1;
  assign _EVAL_243 = 8'h1 << _EVAL_7;
  assign _EVAL_223 = _EVAL_15 & _EVAL_150;
  assign _EVAL_100 = _EVAL_191[0];
  assign _EVAL_203 = {{28'd0}, _EVAL_233};
  assign _EVAL_264 = _EVAL_17 == 3'h6;
  assign _EVAL_45 = _EVAL_234 & _EVAL_216;
  assign _EVAL_220 = ~_EVAL_84;
  assign _EVAL_99 = _EVAL_228 == 2'h0;
  assign _EVAL_35 = _EVAL_19 ? _EVAL_80 : 8'h0;
  assign _EVAL_89 = _EVAL_216 & _EVAL_217;
  assign _EVAL_196 = _EVAL_4 & _EVAL_281;
  assign _EVAL_111 = _EVAL_15 & _EVAL_179;
  assign _EVAL_172 = _EVAL_270 & _EVAL_144;
  assign _EVAL_22 = _EVAL_4 & _EVAL_24;
  assign _EVAL_211 = _EVAL_224 | 2'h1;
  assign _EVAL_106 = _EVAL_8 & _EVAL_4;
  assign _EVAL_24 = _EVAL_12 == 3'h0;
  assign _EVAL_263 = _EVAL_15 & _EVAL_43;
  assign _EVAL_120 = _EVAL_25 | _EVAL_10;
  assign _EVAL_202 = _EVAL_17 <= 3'h6;
  assign _EVAL_221 = _EVAL_18 <= 3'h2;
  assign _EVAL_91 = _EVAL_106 & _EVAL_226;
  assign _EVAL_252 = _EVAL_242[4:0];
  assign _EVAL_60 = _EVAL_178 - 1'h1;
  assign _EVAL_167 = ~_EVAL_205;
  assign _EVAL_86 = _EVAL_133[31:0];
  assign _EVAL_68 = _EVAL_106 & _EVAL_183;
  assign _EVAL_84 = _EVAL_262[0];
  assign _EVAL_73 = ~_EVAL_118;
  assign _EVAL_219 = ~_EVAL_10;
  assign _EVAL_27 = ~_EVAL_189;
  assign _EVAL_62 = ~_EVAL_275;
  assign _EVAL_250 = _EVAL_35[4:0];
  assign _EVAL_269 = _EVAL_134 | _EVAL_10;
  assign _EVAL_201 = ~_EVAL_85;
  assign _EVAL_207 = {_EVAL_176,_EVAL_278,_EVAL_162,_EVAL_174};
  assign _EVAL_142 = _EVAL_158[1:0];
  assign _EVAL_235 = _EVAL_98[0];
  assign _EVAL_166 = _EVAL_16 ^ 30'h20000000;
  assign _EVAL_77 = _EVAL_12 == 3'h3;
  assign _EVAL_105 = _EVAL_146 | _EVAL_10;
  assign _EVAL_204 = ~_EVAL_255;
  assign _EVAL_126 = _EVAL_274 | _EVAL_10;
  assign _EVAL_88 = _EVAL_13 == _EVAL_207;
  assign _EVAL_173 = _EVAL_60[0];
  assign _EVAL_191 = _EVAL_140 >> _EVAL_5;
  assign _EVAL_197 = ~_EVAL_280;
  assign _EVAL_148 = ~_EVAL_44;
  assign _EVAL_39 = _EVAL_125 - 1'h1;
  assign _EVAL_176 = _EVAL_40 | _EVAL_78;
  assign _EVAL_244 = _EVAL_12 == 3'h7;
  assign _EVAL_154 = ~_EVAL_229;
  assign _EVAL_262 = _EVAL_271 >> _EVAL_7;
  assign _EVAL_153 = ~_EVAL_129;
  assign _EVAL_57 = _EVAL_238 | _EVAL_10;
  assign _EVAL_25 = _EVAL_3 >= 2'h2;
  assign _EVAL_52 = ~_EVAL_41;
  assign _EVAL_97 = _EVAL_18 == _EVAL_26;
  assign _EVAL_31 = _EVAL_55 | _EVAL_14;
  assign _EVAL_259 = {1'b0,$signed(_EVAL_166)};
  assign _EVAL_66 = _EVAL_192 == 4'h0;
  assign _EVAL_267 = ~_EVAL_65;
  assign _EVAL_79 = _EVAL_4 & _EVAL_200;
  assign _EVAL_249 = _EVAL_157 & _EVAL_213;
  assign _EVAL_146 = _EVAL == _EVAL_149;
  assign _EVAL_114 = _EVAL_252 != _EVAL_250;
  assign _EVAL_56 = _EVAL_3 == _EVAL_245;
  assign _EVAL_124 = _EVAL_23 == 2'h0;
  assign _EVAL_168 = ~_EVAL_75;
  assign _EVAL_69 = _EVAL_2 == _EVAL_210;
  assign _EVAL_61 = ~_EVAL_120;
  assign _EVAL_246 = ~_EVAL_188;
  assign _EVAL_240 = _EVAL_222 == 30'h0;
  assign _EVAL_135 = ~_EVAL_72;
  assign _EVAL_193 = ~_EVAL_198;
  assign _EVAL_276 = ~_EVAL_265;
  assign _EVAL_234 = _EVAL_211[1];
  assign _EVAL_134 = _EVAL_18 <= 3'h1;
  assign _EVAL_273 = _EVAL_97 | _EVAL_10;
  assign _EVAL_216 = _EVAL_16[1];
  assign _EVAL_157 = _EVAL_211[0];
  assign _EVAL_75 = _EVAL_122 | _EVAL_10;
  assign _EVAL_165 = _EVAL_112 == 4'h0;
  assign _EVAL_113 = _EVAL_12 == 3'h2;
  assign _EVAL_136 = _EVAL_234 & _EVAL_127;
  assign _EVAL_205 = _EVAL_83 | _EVAL_10;
  assign _EVAL_266 = _EVAL_267 | _EVAL_37;
  assign _EVAL_255 = _EVAL_119 | _EVAL_10;
  assign _EVAL_212 = ~_EVAL_161;
  assign _EVAL_48 = ~_EVAL_264;
  assign _EVAL_182 = _EVAL_16[0];
  assign _EVAL_232 = _EVAL_4 & _EVAL_113;
  assign _EVAL_118 = _EVAL_69 | _EVAL_10;
  assign _EVAL_121 = ~_EVAL_33;
  assign _EVAL_147 = _EVAL_39[0];
  assign _EVAL_112 = ~_EVAL_13;
  assign _EVAL_127 = ~_EVAL_216;
  assign _EVAL_192 = _EVAL_13 & _EVAL_67;
  assign _EVAL_46 = _EVAL_12 == 3'h6;
  assign _EVAL_236 = _EVAL_170 | _EVAL_10;
  assign _EVAL_42 = ~_EVAL_186;
  assign _EVAL_279 = _EVAL_18 <= 3'h3;
  assign _EVAL_161 = _EVAL_251 | _EVAL_10;
  assign _EVAL_21 = _EVAL_4 & _EVAL_77;
  assign _EVAL_55 = ~_EVAL;
  assign _EVAL_116 = _EVAL_25 | _EVAL_136;
  assign _EVAL_152 = _EVAL_17 == _EVAL_155;
  assign _EVAL_80 = 8'h1 << _EVAL_5;
  assign _EVAL_208 = ~_EVAL_117;
  assign _EVAL_251 = _EVAL_6 <= 2'h2;
  assign _EVAL_70 = _EVAL_100 | _EVAL_10;
  assign _EVAL_233 = ~_EVAL_142;
  assign _EVAL_30 = _EVAL_51 | _EVAL_10;
  assign _EVAL_96 = _EVAL_123;
  assign _EVAL_195 = _EVAL_12 == _EVAL_87;
  assign _EVAL_270 = _EVAL_3 <= 2'h2;
  assign _EVAL_181 = _EVAL_5 == 3'h4;
  assign _EVAL_94 = ~_EVAL_1;
  assign _EVAL_163 = _EVAL_218 < plusarg_reader_out;
  assign _EVAL_144 = $signed(_EVAL_96) == 31'sh0;
  assign _EVAL_103 = _EVAL_6 == 2'h0;
  assign _EVAL_237 = _EVAL_109 | _EVAL_10;
  assign _EVAL_253 = ~_EVAL_125;
  assign _EVAL_19 = _EVAL_194 & _EVAL_48;
  assign _EVAL_129 = _EVAL_143 | _EVAL_10;
  assign _EVAL_92 = _EVAL_157 & _EVAL_89;
  assign _EVAL_228 = _EVAL_5[2:1];
  assign _EVAL_187 = ~_EVAL_30;
  assign _EVAL_169 = _EVAL_3[0];
  assign _EVAL_277 = _EVAL_157 & _EVAL_53;
  assign _EVAL_158 = 5'h3 << _EVAL_3;
  assign _EVAL_217 = ~_EVAL_182;
  assign _EVAL_190 = _EVAL_7 == 3'h4;
  assign _EVAL_37 = plusarg_reader_out == 32'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_26 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_34 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_50 = _RAND_2[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_64 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_87 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_102 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_125 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_139 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_149 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_155 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_178 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_184 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_210 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_218 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_245 = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_248 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_271 = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_0) begin
    if (_EVAL_68) begin
      _EVAL_26 <= _EVAL_18;
    end
    if (_EVAL_10) begin
      _EVAL_34 <= 1'h0;
    end else if (_EVAL_49) begin
      if (_EVAL_260) begin
        _EVAL_34 <= 1'h0;
      end else begin
        _EVAL_34 <= _EVAL_257;
      end
    end
    if (_EVAL_68) begin
      _EVAL_50 <= _EVAL_16;
    end
    if (_EVAL_159) begin
      _EVAL_64 <= _EVAL_6;
    end
    if (_EVAL_68) begin
      _EVAL_87 <= _EVAL_12;
    end
    if (_EVAL_10) begin
      _EVAL_102 <= 1'h0;
    end else if (_EVAL_106) begin
      if (_EVAL_183) begin
        _EVAL_102 <= 1'h0;
      end else begin
        _EVAL_102 <= _EVAL_235;
      end
    end
    if (_EVAL_10) begin
      _EVAL_125 <= 1'h0;
    end else if (_EVAL_49) begin
      if (_EVAL_253) begin
        _EVAL_125 <= 1'h0;
      end else begin
        _EVAL_125 <= _EVAL_147;
      end
    end
    if (_EVAL_159) begin
      _EVAL_139 <= _EVAL_5;
    end
    if (_EVAL_159) begin
      _EVAL_149 <= _EVAL;
    end
    if (_EVAL_159) begin
      _EVAL_155 <= _EVAL_17;
    end
    if (_EVAL_10) begin
      _EVAL_178 <= 1'h0;
    end else if (_EVAL_106) begin
      if (_EVAL_226) begin
        _EVAL_178 <= 1'h0;
      end else begin
        _EVAL_178 <= _EVAL_173;
      end
    end
    if (_EVAL_159) begin
      _EVAL_184 <= _EVAL_11;
    end
    if (_EVAL_159) begin
      _EVAL_210 <= _EVAL_2;
    end
    if (_EVAL_10) begin
      _EVAL_218 <= 32'h0;
    end else if (_EVAL_54) begin
      _EVAL_218 <= 32'h0;
    end else begin
      _EVAL_218 <= _EVAL_86;
    end
    if (_EVAL_68) begin
      _EVAL_245 <= _EVAL_3;
    end
    if (_EVAL_68) begin
      _EVAL_248 <= _EVAL_7;
    end
    if (_EVAL_10) begin
      _EVAL_271 <= 5'h0;
    end else begin
      _EVAL_271 <= _EVAL_177;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(726b05e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44271cc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3bec1f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c41d06e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80ada1b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46a0ba76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12e86ac5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15d417c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8ce2c91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be8f8114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed56c16b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3f446b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9131e715)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d3882b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7905c29b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c861b24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6d987)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d08f73d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdac62a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f67a31a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(697fbd56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a08790d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1dd1e2ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c27a21bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6325a59a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ff6fa1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4c36ec0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(328382e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b07d1f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b088f8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2cff6a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fce1b93a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ea95895)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(728f2b79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd24bd98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(485e1e34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(635d58ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44a85b46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8eb5ea00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(987cd782)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5955e8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3104f111)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(231b97c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4191dba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c85e4d15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c86fbd40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0e52375)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13f69272)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ac69f00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7389fc80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56f8918c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c56b9ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5988c15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f57ff1f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf6e173a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61fb6e6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb5a5293)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc37bca8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb1789e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd5ee101)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f85e98b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d1d2d58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f580d2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc215928)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2231626)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe0c14c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6eaec1ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2622ad6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e21e8066)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96963ed8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76ef0bd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f896d42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a459ac3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5736169c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1853b52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4cea21e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e79e0502)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5b8013)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f1eb87e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c26594a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd119746)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29636fe7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(feec364c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88440db0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4d35bab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7be5946)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7363448e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a11876f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84ff3c15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e471f2e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f68947c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(712a6637)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77a69c11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
