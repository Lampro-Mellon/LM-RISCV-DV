//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_165(
  input         _EVAL,
  output        _EVAL_0,
  input  [2:0]  _EVAL_1,
  output        _EVAL_2,
  input         _EVAL_3,
  input  [7:0]  _EVAL_4,
  output [31:0] _EVAL_5,
  input         _EVAL_6,
  output        _EVAL_7,
  output [31:0] _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  output        _EVAL_11,
  output [3:0]  _EVAL_12,
  output        _EVAL_13,
  input  [7:0]  _EVAL_14,
  input         _EVAL_15,
  output        _EVAL_16,
  input  [2:0]  _EVAL_17,
  input         _EVAL_18,
  output        _EVAL_19,
  output [31:0] _EVAL_20,
  input         _EVAL_21,
  output [3:0]  _EVAL_22,
  output        _EVAL_23,
  output        _EVAL_24,
  output        _EVAL_25,
  output [31:0] _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  output        _EVAL_30,
  output        _EVAL_31,
  input         _EVAL_32,
  output        _EVAL_33,
  output [2:0]  _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  output        _EVAL_38,
  input  [1:0]  _EVAL_39,
  output        _EVAL_40,
  output        _EVAL_41,
  output        _EVAL_42,
  input  [31:0] _EVAL_43,
  input  [1:0]  _EVAL_44,
  output [3:0]  _EVAL_45,
  output        _EVAL_46,
  output [2:0]  _EVAL_47,
  output        _EVAL_48,
  output [2:0]  _EVAL_49,
  output        _EVAL_50,
  input         _EVAL_51,
  input         _EVAL_52,
  input         _EVAL_53,
  input         _EVAL_54,
  output        _EVAL_55,
  input         _EVAL_56,
  output        _EVAL_57,
  input  [3:0]  _EVAL_58,
  input  [31:0] _EVAL_59,
  output [3:0]  _EVAL_60,
  input  [3:0]  _EVAL_61,
  output [2:0]  _EVAL_62,
  input         _EVAL_63,
  output        _EVAL_64,
  output        _EVAL_65,
  input  [31:0] _EVAL_66,
  output        _EVAL_67
);
  wire  _EVAL_68;
  wire [31:0] widget_1__EVAL;
  wire [2:0] widget_1__EVAL_0;
  wire  widget_1__EVAL_1;
  wire  widget_1__EVAL_2;
  wire  widget_1__EVAL_3;
  wire [1:0] widget_1__EVAL_4;
  wire  widget_1__EVAL_5;
  wire [3:0] widget_1__EVAL_6;
  wire  widget_1__EVAL_7;
  wire  widget_1__EVAL_8;
  wire [2:0] widget_1__EVAL_9;
  wire  widget_1__EVAL_10;
  wire  widget_1__EVAL_11;
  wire  widget_1__EVAL_12;
  wire [1:0] widget_1__EVAL_13;
  wire [2:0] widget_1__EVAL_14;
  wire [3:0] widget_1__EVAL_15;
  wire  widget_1__EVAL_16;
  wire  widget_1__EVAL_17;
  wire  widget_1__EVAL_18;
  wire  widget_1__EVAL_19;
  wire [31:0] widget_1__EVAL_20;
  wire [2:0] widget_1__EVAL_21;
  wire  widget_1__EVAL_22;
  wire  widget_1__EVAL_23;
  wire [2:0] widget_1__EVAL_24;
  wire  widget_1__EVAL_25;
  wire  widget_1__EVAL_26;
  wire [3:0] widget_1__EVAL_27;
  wire [31:0] widget_1__EVAL_28;
  wire [31:0] widget_1__EVAL_29;
  wire  widget_1__EVAL_30;
  wire [31:0] widget_1__EVAL_31;
  wire  widget_1__EVAL_32;
  wire  widget_1__EVAL_33;
  wire  widget_1__EVAL_34;
  wire  widget_1__EVAL_35;
  wire  widget_1__EVAL_36;
  wire [3:0] widget_1__EVAL_37;
  wire  widget_1__EVAL_38;
  wire  widget_1__EVAL_39;
  wire  widget_1__EVAL_40;
  wire  widget_1__EVAL_41;
  wire  widget_1__EVAL_42;
  wire  widget_1__EVAL_43;
  wire  widget_1__EVAL_44;
  wire [31:0] widget_1__EVAL_45;
  wire  widget_1__EVAL_46;
  wire  widget_1__EVAL_47;
  wire  widget_1__EVAL_48;
  wire [3:0] widget_1__EVAL_49;
  wire  widget_1__EVAL_50;
  wire [2:0] widget_1__EVAL_51;
  wire  widget_1__EVAL_52;
  wire  widget_1__EVAL_53;
  wire [3:0] widget_1__EVAL_54;
  wire  _EVAL_77;
  wire  _EVAL_78;
  reg  _EVAL_80;
  reg [31:0] _RAND_0;
  wire  _EVAL_81;
  wire  _EVAL_82;
  reg  _EVAL_83;
  reg [31:0] _RAND_1;
  wire  _EVAL_85;
  wire  _EVAL_90;
  wire  _EVAL_95;
  wire [3:0] _EVAL_98;
  reg  _EVAL_99;
  reg [31:0] _RAND_2;
  wire [2:0] buffer__EVAL;
  wire [3:0] buffer__EVAL_0;
  wire  buffer__EVAL_1;
  wire  buffer__EVAL_2;
  wire  buffer__EVAL_3;
  wire [3:0] buffer__EVAL_4;
  wire [3:0] buffer__EVAL_5;
  wire [31:0] buffer__EVAL_6;
  wire [31:0] buffer__EVAL_7;
  wire  buffer__EVAL_8;
  wire [31:0] buffer__EVAL_9;
  wire [2:0] buffer__EVAL_10;
  wire  buffer__EVAL_11;
  wire  buffer__EVAL_12;
  wire  buffer__EVAL_13;
  wire  buffer__EVAL_14;
  wire [2:0] buffer__EVAL_15;
  wire  buffer__EVAL_16;
  wire  buffer__EVAL_17;
  wire  buffer__EVAL_18;
  wire  buffer__EVAL_19;
  wire  buffer__EVAL_20;
  wire  buffer__EVAL_21;
  wire  buffer__EVAL_22;
  wire  buffer__EVAL_23;
  wire  buffer__EVAL_24;
  wire [3:0] buffer__EVAL_25;
  wire [3:0] buffer__EVAL_26;
  wire [31:0] buffer__EVAL_27;
  wire  buffer__EVAL_28;
  wire  buffer__EVAL_29;
  wire [2:0] buffer__EVAL_30;
  wire  buffer__EVAL_31;
  wire  buffer__EVAL_32;
  wire  buffer__EVAL_33;
  wire  buffer__EVAL_34;
  wire [31:0] buffer__EVAL_35;
  wire [31:0] buffer__EVAL_36;
  wire [31:0] buffer__EVAL_37;
  wire  buffer__EVAL_38;
  wire [1:0] buffer__EVAL_39;
  wire  buffer__EVAL_40;
  wire  buffer__EVAL_41;
  wire  buffer__EVAL_42;
  wire [31:0] buffer__EVAL_43;
  wire  buffer__EVAL_44;
  wire  buffer__EVAL_45;
  wire [2:0] buffer__EVAL_46;
  wire [3:0] buffer__EVAL_47;
  wire [2:0] buffer__EVAL_48;
  wire  buffer__EVAL_49;
  wire  buffer__EVAL_50;
  wire  buffer__EVAL_51;
  wire  buffer__EVAL_52;
  wire  buffer__EVAL_53;
  wire [1:0] buffer__EVAL_54;
  wire  buffer__EVAL_55;
  wire [2:0] buffer__EVAL_56;
  wire [31:0] buffer__EVAL_57;
  wire  buffer__EVAL_58;
  wire  buffer__EVAL_59;
  wire  buffer__EVAL_60;
  wire [3:0] buffer__EVAL_61;
  wire  buffer__EVAL_62;
  wire [31:0] buffer__EVAL_63;
  wire [3:0] buffer__EVAL_64;
  wire  buffer__EVAL_65;
  wire  buffer__EVAL_66;
  wire  buffer__EVAL_67;
  wire  buffer__EVAL_68;
  wire  buffer__EVAL_69;
  wire  buffer__EVAL_70;
  wire  buffer__EVAL_71;
  wire [2:0] buffer__EVAL_72;
  wire [2:0] buffer__EVAL_73;
  wire  buffer__EVAL_74;
  wire  buffer__EVAL_75;
  wire  buffer__EVAL_76;
  wire [3:0] buffer__EVAL_77;
  wire  buffer__EVAL_78;
  wire  buffer__EVAL_79;
  wire  buffer__EVAL_80;
  wire  buffer__EVAL_81;
  wire [1:0] buffer__EVAL_82;
  wire  buffer__EVAL_83;
  wire [3:0] buffer__EVAL_84;
  wire  buffer__EVAL_85;
  wire  buffer__EVAL_86;
  wire [2:0] buffer__EVAL_87;
  wire  buffer__EVAL_88;
  wire  buffer__EVAL_89;
  wire  buffer__EVAL_90;
  wire  buffer__EVAL_91;
  wire [31:0] buffer__EVAL_92;
  wire [3:0] buffer__EVAL_93;
  wire [2:0] buffer__EVAL_94;
  wire [1:0] buffer__EVAL_95;
  wire  buffer__EVAL_96;
  wire  buffer__EVAL_97;
  wire  buffer__EVAL_98;
  wire  buffer__EVAL_99;
  wire [3:0] buffer__EVAL_100;
  wire [2:0] buffer__EVAL_101;
  wire [31:0] buffer__EVAL_102;
  wire  buffer__EVAL_103;
  wire  buffer__EVAL_104;
  wire  buffer__EVAL_105;
  wire  buffer__EVAL_106;
  wire  buffer__EVAL_107;
  wire  buffer__EVAL_108;
  wire  _EVAL_101;
  reg [3:0] _EVAL_102;
  reg [31:0] _RAND_3;
  wire  widget__EVAL;
  wire  widget__EVAL_0;
  wire [2:0] widget__EVAL_1;
  wire  widget__EVAL_2;
  wire [3:0] widget__EVAL_3;
  wire  widget__EVAL_4;
  wire  widget__EVAL_5;
  wire  widget__EVAL_6;
  wire [31:0] widget__EVAL_7;
  wire  widget__EVAL_8;
  wire [1:0] widget__EVAL_9;
  wire [3:0] widget__EVAL_10;
  wire [1:0] widget__EVAL_11;
  wire [31:0] widget__EVAL_12;
  wire  widget__EVAL_13;
  wire  widget__EVAL_14;
  wire  widget__EVAL_15;
  wire  widget__EVAL_16;
  wire  widget__EVAL_17;
  wire  widget__EVAL_18;
  wire [31:0] widget__EVAL_19;
  wire  widget__EVAL_20;
  wire [3:0] widget__EVAL_21;
  wire [3:0] widget__EVAL_22;
  wire  widget__EVAL_23;
  wire  widget__EVAL_24;
  wire  widget__EVAL_25;
  wire [2:0] widget__EVAL_26;
  wire  widget__EVAL_27;
  wire [2:0] widget__EVAL_28;
  wire [3:0] widget__EVAL_29;
  wire [31:0] widget__EVAL_30;
  wire  widget__EVAL_31;
  wire  widget__EVAL_32;
  wire  widget__EVAL_33;
  wire [2:0] widget__EVAL_34;
  wire  widget__EVAL_35;
  wire  widget__EVAL_36;
  wire [2:0] widget__EVAL_37;
  wire [31:0] widget__EVAL_38;
  wire  widget__EVAL_39;
  wire  widget__EVAL_40;
  wire  widget__EVAL_41;
  wire  widget__EVAL_42;
  wire  widget__EVAL_43;
  wire [2:0] widget__EVAL_44;
  wire  widget__EVAL_45;
  wire  widget__EVAL_46;
  wire  widget__EVAL_47;
  wire  widget__EVAL_48;
  wire [31:0] widget__EVAL_49;
  wire  widget__EVAL_50;
  wire [3:0] widget__EVAL_51;
  wire  widget__EVAL_52;
  wire  widget__EVAL_53;
  wire  widget__EVAL_54;
  wire  tile_core_clock_gate_in;
  wire  tile_core_clock_gate_test_en;
  wire  tile_core_clock_gate_en;
  wire  tile_core_clock_gate_out;
  wire  _EVAL_107;
  wire  core__EVAL;
  wire  core__EVAL_0;
  wire [7:0] core__EVAL_1;
  wire [2:0] core__EVAL_2;
  wire  core__EVAL_3;
  wire  core__EVAL_4;
  wire  core__EVAL_5;
  wire [31:0] core__EVAL_6;
  wire [3:0] core__EVAL_7;
  wire  core__EVAL_8;
  wire [2:0] core__EVAL_9;
  wire  core__EVAL_10;
  wire  core__EVAL_11;
  wire  core__EVAL_12;
  wire  core__EVAL_13;
  wire [7:0] core__EVAL_14;
  wire  core__EVAL_15;
  wire  core__EVAL_16;
  wire  core__EVAL_17;
  wire  core__EVAL_18;
  wire [3:0] core__EVAL_19;
  wire  core__EVAL_20;
  wire [31:0] core__EVAL_21;
  wire  core__EVAL_22;
  wire  core__EVAL_23;
  wire  core__EVAL_24;
  wire [1:0] core__EVAL_25;
  wire [2:0] core__EVAL_26;
  wire [2:0] core__EVAL_27;
  wire  core__EVAL_28;
  wire  core__EVAL_29;
  wire  core__EVAL_30;
  wire  core__EVAL_31;
  wire  core__EVAL_32;
  wire  core__EVAL_33;
  wire  core__EVAL_34;
  wire  core__EVAL_35;
  wire  core__EVAL_36;
  wire  core__EVAL_37;
  wire  core__EVAL_38;
  wire  core__EVAL_39;
  wire  core__EVAL_40;
  wire  core__EVAL_41;
  wire  core__EVAL_42;
  wire  core__EVAL_43;
  wire  core__EVAL_44;
  wire [31:0] core__EVAL_45;
  wire  core__EVAL_46;
  wire  core__EVAL_47;
  wire [3:0] core__EVAL_48;
  wire [2:0] core__EVAL_49;
  wire  core__EVAL_50;
  wire [31:0] core__EVAL_51;
  wire  core__EVAL_52;
  wire [31:0] core__EVAL_53;
  wire  core__EVAL_54;
  wire  core__EVAL_55;
  wire [31:0] core__EVAL_56;
  wire  core__EVAL_57;
  wire [3:0] core__EVAL_58;
  wire [3:0] core__EVAL_59;
  wire [31:0] core__EVAL_60;
  wire [1:0] core__EVAL_61;
  wire [3:0] core__EVAL_62;
  wire  core__EVAL_63;
  wire  core__EVAL_64;
  wire  core__EVAL_65;
  wire  core__EVAL_66;
  wire  core__EVAL_67;
  wire [2:0] core__EVAL_68;
  wire  _EVAL_115;
  wire [4:0] _EVAL_116;
  wire  _EVAL_118;
  _EVAL_162 widget_1 (
    ._EVAL(widget_1__EVAL),
    ._EVAL_0(widget_1__EVAL_0),
    ._EVAL_1(widget_1__EVAL_1),
    ._EVAL_2(widget_1__EVAL_2),
    ._EVAL_3(widget_1__EVAL_3),
    ._EVAL_4(widget_1__EVAL_4),
    ._EVAL_5(widget_1__EVAL_5),
    ._EVAL_6(widget_1__EVAL_6),
    ._EVAL_7(widget_1__EVAL_7),
    ._EVAL_8(widget_1__EVAL_8),
    ._EVAL_9(widget_1__EVAL_9),
    ._EVAL_10(widget_1__EVAL_10),
    ._EVAL_11(widget_1__EVAL_11),
    ._EVAL_12(widget_1__EVAL_12),
    ._EVAL_13(widget_1__EVAL_13),
    ._EVAL_14(widget_1__EVAL_14),
    ._EVAL_15(widget_1__EVAL_15),
    ._EVAL_16(widget_1__EVAL_16),
    ._EVAL_17(widget_1__EVAL_17),
    ._EVAL_18(widget_1__EVAL_18),
    ._EVAL_19(widget_1__EVAL_19),
    ._EVAL_20(widget_1__EVAL_20),
    ._EVAL_21(widget_1__EVAL_21),
    ._EVAL_22(widget_1__EVAL_22),
    ._EVAL_23(widget_1__EVAL_23),
    ._EVAL_24(widget_1__EVAL_24),
    ._EVAL_25(widget_1__EVAL_25),
    ._EVAL_26(widget_1__EVAL_26),
    ._EVAL_27(widget_1__EVAL_27),
    ._EVAL_28(widget_1__EVAL_28),
    ._EVAL_29(widget_1__EVAL_29),
    ._EVAL_30(widget_1__EVAL_30),
    ._EVAL_31(widget_1__EVAL_31),
    ._EVAL_32(widget_1__EVAL_32),
    ._EVAL_33(widget_1__EVAL_33),
    ._EVAL_34(widget_1__EVAL_34),
    ._EVAL_35(widget_1__EVAL_35),
    ._EVAL_36(widget_1__EVAL_36),
    ._EVAL_37(widget_1__EVAL_37),
    ._EVAL_38(widget_1__EVAL_38),
    ._EVAL_39(widget_1__EVAL_39),
    ._EVAL_40(widget_1__EVAL_40),
    ._EVAL_41(widget_1__EVAL_41),
    ._EVAL_42(widget_1__EVAL_42),
    ._EVAL_43(widget_1__EVAL_43),
    ._EVAL_44(widget_1__EVAL_44),
    ._EVAL_45(widget_1__EVAL_45),
    ._EVAL_46(widget_1__EVAL_46),
    ._EVAL_47(widget_1__EVAL_47),
    ._EVAL_48(widget_1__EVAL_48),
    ._EVAL_49(widget_1__EVAL_49),
    ._EVAL_50(widget_1__EVAL_50),
    ._EVAL_51(widget_1__EVAL_51),
    ._EVAL_52(widget_1__EVAL_52),
    ._EVAL_53(widget_1__EVAL_53),
    ._EVAL_54(widget_1__EVAL_54)
  );
  _EVAL_164 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32),
    ._EVAL_33(buffer__EVAL_33),
    ._EVAL_34(buffer__EVAL_34),
    ._EVAL_35(buffer__EVAL_35),
    ._EVAL_36(buffer__EVAL_36),
    ._EVAL_37(buffer__EVAL_37),
    ._EVAL_38(buffer__EVAL_38),
    ._EVAL_39(buffer__EVAL_39),
    ._EVAL_40(buffer__EVAL_40),
    ._EVAL_41(buffer__EVAL_41),
    ._EVAL_42(buffer__EVAL_42),
    ._EVAL_43(buffer__EVAL_43),
    ._EVAL_44(buffer__EVAL_44),
    ._EVAL_45(buffer__EVAL_45),
    ._EVAL_46(buffer__EVAL_46),
    ._EVAL_47(buffer__EVAL_47),
    ._EVAL_48(buffer__EVAL_48),
    ._EVAL_49(buffer__EVAL_49),
    ._EVAL_50(buffer__EVAL_50),
    ._EVAL_51(buffer__EVAL_51),
    ._EVAL_52(buffer__EVAL_52),
    ._EVAL_53(buffer__EVAL_53),
    ._EVAL_54(buffer__EVAL_54),
    ._EVAL_55(buffer__EVAL_55),
    ._EVAL_56(buffer__EVAL_56),
    ._EVAL_57(buffer__EVAL_57),
    ._EVAL_58(buffer__EVAL_58),
    ._EVAL_59(buffer__EVAL_59),
    ._EVAL_60(buffer__EVAL_60),
    ._EVAL_61(buffer__EVAL_61),
    ._EVAL_62(buffer__EVAL_62),
    ._EVAL_63(buffer__EVAL_63),
    ._EVAL_64(buffer__EVAL_64),
    ._EVAL_65(buffer__EVAL_65),
    ._EVAL_66(buffer__EVAL_66),
    ._EVAL_67(buffer__EVAL_67),
    ._EVAL_68(buffer__EVAL_68),
    ._EVAL_69(buffer__EVAL_69),
    ._EVAL_70(buffer__EVAL_70),
    ._EVAL_71(buffer__EVAL_71),
    ._EVAL_72(buffer__EVAL_72),
    ._EVAL_73(buffer__EVAL_73),
    ._EVAL_74(buffer__EVAL_74),
    ._EVAL_75(buffer__EVAL_75),
    ._EVAL_76(buffer__EVAL_76),
    ._EVAL_77(buffer__EVAL_77),
    ._EVAL_78(buffer__EVAL_78),
    ._EVAL_79(buffer__EVAL_79),
    ._EVAL_80(buffer__EVAL_80),
    ._EVAL_81(buffer__EVAL_81),
    ._EVAL_82(buffer__EVAL_82),
    ._EVAL_83(buffer__EVAL_83),
    ._EVAL_84(buffer__EVAL_84),
    ._EVAL_85(buffer__EVAL_85),
    ._EVAL_86(buffer__EVAL_86),
    ._EVAL_87(buffer__EVAL_87),
    ._EVAL_88(buffer__EVAL_88),
    ._EVAL_89(buffer__EVAL_89),
    ._EVAL_90(buffer__EVAL_90),
    ._EVAL_91(buffer__EVAL_91),
    ._EVAL_92(buffer__EVAL_92),
    ._EVAL_93(buffer__EVAL_93),
    ._EVAL_94(buffer__EVAL_94),
    ._EVAL_95(buffer__EVAL_95),
    ._EVAL_96(buffer__EVAL_96),
    ._EVAL_97(buffer__EVAL_97),
    ._EVAL_98(buffer__EVAL_98),
    ._EVAL_99(buffer__EVAL_99),
    ._EVAL_100(buffer__EVAL_100),
    ._EVAL_101(buffer__EVAL_101),
    ._EVAL_102(buffer__EVAL_102),
    ._EVAL_103(buffer__EVAL_103),
    ._EVAL_104(buffer__EVAL_104),
    ._EVAL_105(buffer__EVAL_105),
    ._EVAL_106(buffer__EVAL_106),
    ._EVAL_107(buffer__EVAL_107),
    ._EVAL_108(buffer__EVAL_108)
  );
  _EVAL_160 widget (
    ._EVAL(widget__EVAL),
    ._EVAL_0(widget__EVAL_0),
    ._EVAL_1(widget__EVAL_1),
    ._EVAL_2(widget__EVAL_2),
    ._EVAL_3(widget__EVAL_3),
    ._EVAL_4(widget__EVAL_4),
    ._EVAL_5(widget__EVAL_5),
    ._EVAL_6(widget__EVAL_6),
    ._EVAL_7(widget__EVAL_7),
    ._EVAL_8(widget__EVAL_8),
    ._EVAL_9(widget__EVAL_9),
    ._EVAL_10(widget__EVAL_10),
    ._EVAL_11(widget__EVAL_11),
    ._EVAL_12(widget__EVAL_12),
    ._EVAL_13(widget__EVAL_13),
    ._EVAL_14(widget__EVAL_14),
    ._EVAL_15(widget__EVAL_15),
    ._EVAL_16(widget__EVAL_16),
    ._EVAL_17(widget__EVAL_17),
    ._EVAL_18(widget__EVAL_18),
    ._EVAL_19(widget__EVAL_19),
    ._EVAL_20(widget__EVAL_20),
    ._EVAL_21(widget__EVAL_21),
    ._EVAL_22(widget__EVAL_22),
    ._EVAL_23(widget__EVAL_23),
    ._EVAL_24(widget__EVAL_24),
    ._EVAL_25(widget__EVAL_25),
    ._EVAL_26(widget__EVAL_26),
    ._EVAL_27(widget__EVAL_27),
    ._EVAL_28(widget__EVAL_28),
    ._EVAL_29(widget__EVAL_29),
    ._EVAL_30(widget__EVAL_30),
    ._EVAL_31(widget__EVAL_31),
    ._EVAL_32(widget__EVAL_32),
    ._EVAL_33(widget__EVAL_33),
    ._EVAL_34(widget__EVAL_34),
    ._EVAL_35(widget__EVAL_35),
    ._EVAL_36(widget__EVAL_36),
    ._EVAL_37(widget__EVAL_37),
    ._EVAL_38(widget__EVAL_38),
    ._EVAL_39(widget__EVAL_39),
    ._EVAL_40(widget__EVAL_40),
    ._EVAL_41(widget__EVAL_41),
    ._EVAL_42(widget__EVAL_42),
    ._EVAL_43(widget__EVAL_43),
    ._EVAL_44(widget__EVAL_44),
    ._EVAL_45(widget__EVAL_45),
    ._EVAL_46(widget__EVAL_46),
    ._EVAL_47(widget__EVAL_47),
    ._EVAL_48(widget__EVAL_48),
    ._EVAL_49(widget__EVAL_49),
    ._EVAL_50(widget__EVAL_50),
    ._EVAL_51(widget__EVAL_51),
    ._EVAL_52(widget__EVAL_52),
    ._EVAL_53(widget__EVAL_53),
    ._EVAL_54(widget__EVAL_54)
  );
  EICG_wrapper tile_core_clock_gate (
    .in(tile_core_clock_gate_in),
    .test_en(tile_core_clock_gate_test_en),
    .en(tile_core_clock_gate_en),
    .out(tile_core_clock_gate_out)
  );
  _EVAL_158 core (
    ._EVAL(core__EVAL),
    ._EVAL_0(core__EVAL_0),
    ._EVAL_1(core__EVAL_1),
    ._EVAL_2(core__EVAL_2),
    ._EVAL_3(core__EVAL_3),
    ._EVAL_4(core__EVAL_4),
    ._EVAL_5(core__EVAL_5),
    ._EVAL_6(core__EVAL_6),
    ._EVAL_7(core__EVAL_7),
    ._EVAL_8(core__EVAL_8),
    ._EVAL_9(core__EVAL_9),
    ._EVAL_10(core__EVAL_10),
    ._EVAL_11(core__EVAL_11),
    ._EVAL_12(core__EVAL_12),
    ._EVAL_13(core__EVAL_13),
    ._EVAL_14(core__EVAL_14),
    ._EVAL_15(core__EVAL_15),
    ._EVAL_16(core__EVAL_16),
    ._EVAL_17(core__EVAL_17),
    ._EVAL_18(core__EVAL_18),
    ._EVAL_19(core__EVAL_19),
    ._EVAL_20(core__EVAL_20),
    ._EVAL_21(core__EVAL_21),
    ._EVAL_22(core__EVAL_22),
    ._EVAL_23(core__EVAL_23),
    ._EVAL_24(core__EVAL_24),
    ._EVAL_25(core__EVAL_25),
    ._EVAL_26(core__EVAL_26),
    ._EVAL_27(core__EVAL_27),
    ._EVAL_28(core__EVAL_28),
    ._EVAL_29(core__EVAL_29),
    ._EVAL_30(core__EVAL_30),
    ._EVAL_31(core__EVAL_31),
    ._EVAL_32(core__EVAL_32),
    ._EVAL_33(core__EVAL_33),
    ._EVAL_34(core__EVAL_34),
    ._EVAL_35(core__EVAL_35),
    ._EVAL_36(core__EVAL_36),
    ._EVAL_37(core__EVAL_37),
    ._EVAL_38(core__EVAL_38),
    ._EVAL_39(core__EVAL_39),
    ._EVAL_40(core__EVAL_40),
    ._EVAL_41(core__EVAL_41),
    ._EVAL_42(core__EVAL_42),
    ._EVAL_43(core__EVAL_43),
    ._EVAL_44(core__EVAL_44),
    ._EVAL_45(core__EVAL_45),
    ._EVAL_46(core__EVAL_46),
    ._EVAL_47(core__EVAL_47),
    ._EVAL_48(core__EVAL_48),
    ._EVAL_49(core__EVAL_49),
    ._EVAL_50(core__EVAL_50),
    ._EVAL_51(core__EVAL_51),
    ._EVAL_52(core__EVAL_52),
    ._EVAL_53(core__EVAL_53),
    ._EVAL_54(core__EVAL_54),
    ._EVAL_55(core__EVAL_55),
    ._EVAL_56(core__EVAL_56),
    ._EVAL_57(core__EVAL_57),
    ._EVAL_58(core__EVAL_58),
    ._EVAL_59(core__EVAL_59),
    ._EVAL_60(core__EVAL_60),
    ._EVAL_61(core__EVAL_61),
    ._EVAL_62(core__EVAL_62),
    ._EVAL_63(core__EVAL_63),
    ._EVAL_64(core__EVAL_64),
    ._EVAL_65(core__EVAL_65),
    ._EVAL_66(core__EVAL_66),
    ._EVAL_67(core__EVAL_67),
    ._EVAL_68(core__EVAL_68)
  );
  assign buffer__EVAL_24 = widget__EVAL_43;
  assign widget_1__EVAL_25 = core__EVAL_22;
  assign widget_1__EVAL_44 = buffer__EVAL_76;
  assign buffer__EVAL_98 = widget_1__EVAL_22;
  assign _EVAL_90 = _EVAL_102 >= 4'h8;
  assign _EVAL_67 = buffer__EVAL_80;
  assign core__EVAL_35 = widget__EVAL_33;
  assign buffer__EVAL_19 = widget__EVAL_40;
  assign widget__EVAL_29 = buffer__EVAL_64;
  assign widget_1__EVAL_28 = core__EVAL_6;
  assign buffer__EVAL_48 = _EVAL_17;
  assign buffer__EVAL_27 = widget_1__EVAL_45;
  assign buffer__EVAL_90 = _EVAL_6;
  assign widget_1__EVAL_21 = buffer__EVAL_87;
  assign _EVAL_85 = core__EVAL_54 | _EVAL_99;
  assign core__EVAL_53 = widget_1__EVAL_20;
  assign core__EVAL_32 = widget__EVAL_25;
  assign buffer__EVAL_58 = _EVAL_15;
  assign widget__EVAL_36 = core__EVAL_18;
  assign widget_1__EVAL_35 = buffer__EVAL_2;
  assign widget_1__EVAL_27 = buffer__EVAL_47;
  assign widget_1__EVAL_40 = buffer__EVAL_86;
  assign core__EVAL_67 = widget__EVAL_15;
  assign buffer__EVAL_34 = widget_1__EVAL_33;
  assign core__EVAL_8 = _EVAL_52;
  assign buffer__EVAL_96 = widget__EVAL_31;
  assign buffer__EVAL_15 = _EVAL_1;
  assign core__EVAL_57 = _EVAL_3;
  assign core__EVAL_47 = widget__EVAL_18;
  assign widget__EVAL_21 = core__EVAL_19;
  assign widget__EVAL_41 = core__EVAL_10;
  assign _EVAL_33 = _EVAL_83;
  assign core__EVAL_60 = widget__EVAL_19;
  assign _EVAL_95 = ~core__EVAL_34;
  assign widget_1__EVAL_7 = buffer__EVAL_99;
  assign buffer__EVAL_38 = widget_1__EVAL_41;
  assign buffer__EVAL_41 = _EVAL_29;
  assign _EVAL_45 = buffer__EVAL_93;
  assign _EVAL_8 = buffer__EVAL_9;
  assign widget_1__EVAL_29 = core__EVAL_45;
  assign _EVAL_115 = _EVAL_81 | _EVAL_82;
  assign widget__EVAL_49 = core__EVAL_21;
  assign _EVAL_7 = _EVAL_99;
  assign widget_1__EVAL_54 = core__EVAL_58;
  assign buffer__EVAL = widget__EVAL_44;
  assign core__EVAL_14 = _EVAL_14;
  assign _EVAL_30 = buffer__EVAL_32;
  assign _EVAL_5 = buffer__EVAL_36;
  assign widget__EVAL_38 = buffer__EVAL_57;
  assign core__EVAL_2 = widget__EVAL_34;
  assign buffer__EVAL_59 = widget_1__EVAL_48;
  assign _EVAL_20 = buffer__EVAL_63;
  assign widget__EVAL_37 = core__EVAL_9;
  assign _EVAL_62 = buffer__EVAL_30;
  assign core__EVAL_36 = tile_core_clock_gate_out;
  assign buffer__EVAL_61 = widget__EVAL_10;
  assign _EVAL_16 = buffer__EVAL_97;
  assign buffer__EVAL_100 = widget_1__EVAL_15;
  assign core__EVAL_31 = widget__EVAL_46;
  assign _EVAL_77 = _EVAL_4 != 8'h0;
  assign widget__EVAL_22 = core__EVAL_59;
  assign buffer__EVAL_75 = widget_1__EVAL_12;
  assign _EVAL_42 = buffer__EVAL_18;
  assign buffer__EVAL_105 = _EVAL_32;
  assign tile_core_clock_gate_test_en = _EVAL_10;
  assign widget__EVAL_47 = core__EVAL_5;
  assign core__EVAL_16 = _EVAL_51;
  assign widget__EVAL_27 = _EVAL_32;
  assign widget__EVAL_23 = buffer__EVAL_17;
  assign buffer__EVAL_66 = widget_1__EVAL_30;
  assign _EVAL_55 = _EVAL_102 >= 4'h8;
  assign widget_1__EVAL = buffer__EVAL_37;
  assign buffer__EVAL_71 = widget__EVAL;
  assign widget__EVAL_0 = core__EVAL_37;
  assign _EVAL_41 = buffer__EVAL_70;
  assign widget_1__EVAL_0 = core__EVAL_49;
  assign widget__EVAL_1 = core__EVAL_27;
  assign _EVAL_31 = buffer__EVAL_3;
  assign widget__EVAL_6 = core__EVAL_44;
  assign buffer__EVAL_16 = widget_1__EVAL_46;
  assign core__EVAL_40 = _EVAL;
  assign buffer__EVAL_43 = _EVAL_59;
  assign widget__EVAL_45 = buffer__EVAL_50;
  assign widget_1__EVAL_13 = buffer__EVAL_54;
  assign widget_1__EVAL_42 = core__EVAL_42;
  assign buffer__EVAL_84 = _EVAL_58;
  assign buffer__EVAL_21 = _EVAL_53;
  assign buffer__EVAL_62 = _EVAL_56;
  assign widget_1__EVAL_34 = buffer__EVAL_60;
  assign widget_1__EVAL_14 = core__EVAL_26;
  assign core__EVAL_13 = _EVAL_63;
  assign _EVAL_98 = _EVAL_116[3:0];
  assign buffer__EVAL_85 = _EVAL_21;
  assign core__EVAL_23 = widget_1__EVAL_17;
  assign widget__EVAL_2 = _EVAL_21;
  assign buffer__EVAL_26 = _EVAL_61;
  assign widget_1__EVAL_38 = core__EVAL_39;
  assign widget_1__EVAL_37 = core__EVAL_62;
  assign buffer__EVAL_0 = widget_1__EVAL_6;
  assign buffer__EVAL_102 = _EVAL_43;
  assign _EVAL_2 = buffer__EVAL_69;
  assign widget__EVAL_14 = core__EVAL_3;
  assign buffer__EVAL_92 = widget__EVAL_30;
  assign core__EVAL_68 = widget_1__EVAL_9;
  assign core__EVAL_12 = widget_1__EVAL_52;
  assign buffer__EVAL_35 = widget_1__EVAL_31;
  assign widget__EVAL_16 = core__EVAL_41;
  assign widget_1__EVAL_8 = core__EVAL_24;
  assign buffer__EVAL_106 = _EVAL_9;
  assign _EVAL_0 = buffer__EVAL_68;
  assign widget_1__EVAL_10 = core__EVAL_33;
  assign widget__EVAL_42 = buffer__EVAL_81;
  assign _EVAL_25 = buffer__EVAL_108;
  assign buffer__EVAL_14 = widget_1__EVAL_1;
  assign _EVAL_101 = _EVAL_68 | _EVAL_52;
  assign buffer__EVAL_44 = _EVAL_28;
  assign tile_core_clock_gate_in = _EVAL_21;
  assign buffer__EVAL_91 = widget__EVAL_48;
  assign core__EVAL_51 = _EVAL_66;
  assign buffer__EVAL_40 = _EVAL_54;
  assign widget__EVAL_11 = buffer__EVAL_95;
  assign _EVAL_60 = buffer__EVAL_5;
  assign widget__EVAL_13 = core__EVAL_66;
  assign buffer__EVAL_53 = widget__EVAL_35;
  assign _EVAL_12 = buffer__EVAL_4;
  assign widget__EVAL_24 = buffer__EVAL_22;
  assign buffer__EVAL_94 = widget_1__EVAL_51;
  assign buffer__EVAL_31 = widget_1__EVAL_5;
  assign buffer__EVAL_10 = widget__EVAL_26;
  assign buffer__EVAL_1 = widget_1__EVAL_43;
  assign core__EVAL_61 = widget_1__EVAL_4;
  assign core__EVAL_25 = widget__EVAL_9;
  assign widget__EVAL_4 = core__EVAL_52;
  assign _EVAL_81 = ~core__EVAL_28;
  assign buffer__EVAL_20 = widget__EVAL_5;
  assign _EVAL_22 = buffer__EVAL_77;
  assign _EVAL_19 = buffer__EVAL_49;
  assign core__EVAL_55 = widget_1__EVAL_32;
  assign _EVAL_68 = _EVAL_51 | _EVAL;
  assign buffer__EVAL_82 = _EVAL_39;
  assign widget__EVAL_53 = buffer__EVAL_51;
  assign buffer__EVAL_104 = widget__EVAL_50;
  assign buffer__EVAL_72 = widget_1__EVAL_24;
  assign buffer__EVAL_25 = widget__EVAL_3;
  assign widget_1__EVAL_47 = core__EVAL_0;
  assign widget_1__EVAL_36 = _EVAL_21;
  assign widget_1__EVAL_16 = core__EVAL_38;
  assign widget__EVAL_7 = core__EVAL_56;
  assign _EVAL_65 = buffer__EVAL_78;
  assign core__EVAL_64 = _EVAL_32;
  assign widget__EVAL_54 = buffer__EVAL_23;
  assign widget_1__EVAL_18 = buffer__EVAL_89;
  assign _EVAL_38 = buffer__EVAL_79;
  assign widget_1__EVAL_53 = core__EVAL_63;
  assign widget_1__EVAL_11 = _EVAL_32;
  assign _EVAL_107 = core__EVAL_34 & _EVAL_78;
  assign _EVAL_118 = _EVAL_101 | _EVAL_35;
  assign buffer__EVAL_52 = widget__EVAL_17;
  assign buffer__EVAL_28 = _EVAL_18;
  assign core__EVAL_7 = widget_1__EVAL_49;
  assign buffer__EVAL_74 = widget__EVAL_39;
  assign buffer__EVAL_45 = _EVAL_27;
  assign core__EVAL_1 = _EVAL_4;
  assign widget_1__EVAL_19 = core__EVAL_65;
  assign widget__EVAL_28 = buffer__EVAL_56;
  assign buffer__EVAL_6 = widget__EVAL_12;
  assign _EVAL_46 = buffer__EVAL_42;
  assign _EVAL_82 = _EVAL_118 | _EVAL_77;
  assign _EVAL_34 = buffer__EVAL_101;
  assign _EVAL_49 = buffer__EVAL_46;
  assign widget_1__EVAL_39 = core__EVAL_43;
  assign buffer__EVAL_11 = _EVAL_36;
  assign _EVAL_78 = ~_EVAL_90;
  assign core__EVAL = widget_1__EVAL_23;
  assign core__EVAL_17 = widget_1__EVAL_50;
  assign _EVAL_40 = buffer__EVAL_107;
  assign _EVAL_116 = _EVAL_102 + 4'h1;
  assign tile_core_clock_gate_en = _EVAL_115 | _EVAL_80;
  assign _EVAL_26 = buffer__EVAL_7;
  assign _EVAL_50 = buffer__EVAL_8;
  assign buffer__EVAL_65 = widget__EVAL_32;
  assign _EVAL_47 = buffer__EVAL_73;
  assign widget_1__EVAL_26 = core__EVAL_4;
  assign buffer__EVAL_39 = _EVAL_44;
  assign _EVAL_11 = buffer__EVAL_55;
  assign _EVAL_48 = buffer__EVAL_83;
  assign core__EVAL_11 = widget_1__EVAL_2;
  assign buffer__EVAL_67 = widget_1__EVAL_3;
  assign core__EVAL_29 = widget__EVAL_20;
  assign buffer__EVAL_103 = _EVAL_37;
  assign _EVAL_24 = buffer__EVAL_12;
  assign _EVAL_13 = buffer__EVAL_33;
  assign core__EVAL_20 = _EVAL_35;
  assign _EVAL_64 = buffer__EVAL_88;
  assign _EVAL_23 = buffer__EVAL_29;
  assign widget__EVAL_52 = core__EVAL_15;
  assign _EVAL_57 = buffer__EVAL_13;
  assign widget__EVAL_8 = core__EVAL_46;
  assign core__EVAL_48 = widget__EVAL_51;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_80 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_83 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_99 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_102 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_21) begin
    _EVAL_80 <= _EVAL_32;
    if (_EVAL_32) begin
      _EVAL_83 <= 1'h0;
    end else begin
      _EVAL_83 <= core__EVAL_28;
    end
    if (_EVAL_32) begin
      _EVAL_99 <= 1'h0;
    end else begin
      _EVAL_99 <= _EVAL_85;
    end
    if (_EVAL_32) begin
      _EVAL_102 <= 4'h0;
    end else if (_EVAL_107) begin
      _EVAL_102 <= _EVAL_98;
    end else if (_EVAL_95) begin
      _EVAL_102 <= 4'h0;
    end
  end
endmodule
