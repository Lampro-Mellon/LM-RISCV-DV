//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_166_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [31:0] _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [2:0]  _EVAL_8,
  input         _EVAL_9,
  input  [3:0]  _EVAL_10,
  input  [1:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input  [1:0]  _EVAL_14
);
  wire [4:0] _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  reg  _EVAL_21;
  reg [31:0] _RAND_0;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire [1:0] _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire [4:0] _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire [1:0] _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire [31:0] _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire [4:0] _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire [32:0] _EVAL_59;
  wire  _EVAL_60;
  wire [4:0] _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire [7:0] _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  reg [1:0] _EVAL_78;
  reg [31:0] _RAND_1;
  wire [32:0] _EVAL_79;
  reg [4:0] _EVAL_80;
  reg [31:0] _RAND_2;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire [4:0] _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire [7:0] _EVAL_88;
  wire  _EVAL_89;
  wire [1:0] _EVAL_90;
  wire  _EVAL_91;
  wire [32:0] _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire [32:0] _EVAL_105;
  wire [3:0] _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire [7:0] _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_113;
  wire [3:0] _EVAL_114;
  wire [3:0] _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  reg  _EVAL_125;
  reg [31:0] _RAND_3;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire [1:0] _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire [1:0] _EVAL_149;
  wire  _EVAL_150;
  wire [4:0] _EVAL_152;
  reg [2:0] _EVAL_153;
  reg [31:0] _RAND_4;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire [4:0] _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire [31:0] _EVAL_160;
  wire  _EVAL_161;
  reg [2:0] _EVAL_162;
  reg [31:0] _RAND_5;
  wire  _EVAL_163;
  wire [1:0] _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  reg  _EVAL_170;
  reg [31:0] _RAND_6;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  reg [2:0] _EVAL_176;
  reg [31:0] _RAND_7;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire [31:0] _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  reg [2:0] _EVAL_185;
  reg [31:0] _RAND_8;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire [3:0] _EVAL_193;
  reg [1:0] _EVAL_194;
  reg [31:0] _RAND_9;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire [1:0] _EVAL_199;
  wire [31:0] _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire [4:0] _EVAL_204;
  wire  _EVAL_205;
  reg [31:0] _EVAL_207;
  reg [31:0] _RAND_10;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  reg  _EVAL_217;
  reg [31:0] _RAND_11;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  reg [31:0] _EVAL_221;
  reg [31:0] _RAND_12;
  wire  _EVAL_222;
  wire  _EVAL_223;
  reg [2:0] _EVAL_224;
  reg [31:0] _RAND_13;
  wire [7:0] _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire [4:0] _EVAL_240;
  wire [1:0] _EVAL_241;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_227 = _EVAL_5 == _EVAL_221;
  assign _EVAL_203 = _EVAL_147 | _EVAL;
  assign _EVAL_140 = _EVAL_0 & _EVAL_135;
  assign _EVAL_117 = _EVAL_121 | _EVAL;
  assign _EVAL_229 = _EVAL_8 <= 3'h1;
  assign _EVAL_155 = ~_EVAL_21;
  assign _EVAL_238 = _EVAL_149[0];
  assign _EVAL_90 = ~_EVAL_199;
  assign _EVAL_45 = _EVAL_12 == 3'h6;
  assign _EVAL_181 = _EVAL_2 <= 3'h4;
  assign _EVAL_51 = ~_EVAL_47;
  assign _EVAL_173 = _EVAL_11 <= 2'h2;
  assign _EVAL_219 = _EVAL_208 | _EVAL_89;
  assign _EVAL_234 = ~_EVAL_75;
  assign _EVAL_96 = $signed(_EVAL_105) == 33'sh0;
  assign _EVAL_74 = _EVAL_8 <= 3'h3;
  assign _EVAL_68 = _EVAL_31 != 5'h0;
  assign _EVAL_47 = _EVAL_50 | _EVAL;
  assign _EVAL_26 = _EVAL_172 & _EVAL_35;
  assign _EVAL_22 = _EVAL_12 == 3'h2;
  assign _EVAL_113 = ~_EVAL_197;
  assign _EVAL_154 = _EVAL_0 & _EVAL_32;
  assign _EVAL_174 = _EVAL_3 & _EVAL_9;
  assign _EVAL_156 = _EVAL_130 & _EVAL_98;
  assign _EVAL_34 = _EVAL_43 | _EVAL;
  assign _EVAL_42 = _EVAL_59[31:0];
  assign _EVAL_169 = _EVAL_159 | _EVAL;
  assign _EVAL_215 = _EVAL_157[0];
  assign _EVAL_142 = _EVAL_4 == 3'h1;
  assign _EVAL_27 = ~_EVAL_223;
  assign _EVAL_188 = ~_EVAL_73;
  assign _EVAL_89 = _EVAL_178 & _EVAL_53;
  assign _EVAL_73 = _EVAL_181 | _EVAL;
  assign _EVAL_163 = _EVAL_15[0];
  assign _EVAL_187 = ~_EVAL_217;
  assign _EVAL_119 = ~_EVAL_203;
  assign _EVAL_64 = _EVAL_5[0];
  assign _EVAL_161 = _EVAL_178 & _EVAL_201;
  assign _EVAL_86 = _EVAL_230 | _EVAL;
  assign _EVAL_53 = _EVAL_130 & _EVAL_64;
  assign _EVAL_180 = {{30'd0}, _EVAL_90};
  assign _EVAL_226 = _EVAL_12 == 3'h5;
  assign _EVAL_92 = $signed(_EVAL_79) & -33'sh4000;
  assign _EVAL_108 = _EVAL_31 != _EVAL_240;
  assign _EVAL_93 = _EVAL_200 == 32'h0;
  assign _EVAL_208 = _EVAL_111 | _EVAL_124;
  assign _EVAL_56 = ~_EVAL_86;
  assign _EVAL_62 = _EVAL_207 < plusarg_reader_out;
  assign _EVAL_209 = plusarg_reader_out == 32'h0;
  assign _EVAL_81 = ~_EVAL_169;
  assign _EVAL_130 = _EVAL_5[1];
  assign _EVAL_134 = _EVAL_11 == _EVAL_78;
  assign _EVAL_36 = _EVAL_74 | _EVAL;
  assign _EVAL_123 = ~_EVAL_125;
  assign _EVAL_201 = _EVAL_55 & _EVAL_98;
  assign _EVAL_107 = _EVAL_55 & _EVAL_64;
  assign _EVAL_144 = _EVAL_0 & _EVAL_118;
  assign _EVAL_52 = ~_EVAL_40;
  assign _EVAL_103 = _EVAL_210 & _EVAL_187;
  assign _EVAL_149 = _EVAL_170 - 1'h1;
  assign _EVAL_60 = ~_EVAL_69;
  assign _EVAL_199 = _EVAL_152[1:0];
  assign _EVAL_16 = _EVAL_178 & _EVAL_107;
  assign _EVAL_33 = ~_EVAL_101;
  assign _EVAL_204 = _EVAL_61 & _EVAL_54;
  assign _EVAL_197 = _EVAL_177 | _EVAL;
  assign _EVAL_210 = _EVAL_13 & _EVAL_0;
  assign _EVAL_17 = _EVAL_229 | _EVAL;
  assign _EVAL_136 = _EVAL_134 | _EVAL;
  assign _EVAL_84 = _EVAL_31 | _EVAL_80;
  assign _EVAL_160 = _EVAL_5 ^ 32'h80000000;
  assign _EVAL_91 = _EVAL_137[0];
  assign _EVAL_72 = ~_EVAL_218;
  assign _EVAL_240 = _EVAL_225[4:0];
  assign _EVAL_70 = ~_EVAL_36;
  assign _EVAL_127 = _EVAL_163 | _EVAL;
  assign _EVAL_46 = _EVAL_233 | _EVAL_209;
  assign _EVAL_137 = _EVAL_217 - 1'h1;
  assign _EVAL_39 = ~_EVAL_127;
  assign _EVAL_183 = _EVAL_111 | _EVAL;
  assign _EVAL_23 = ~_EVAL_215;
  assign _EVAL_43 = _EVAL_7 <= 3'h4;
  assign _EVAL_212 = _EVAL_0 & _EVAL_182;
  assign _EVAL_94 = _EVAL_44 | _EVAL;
  assign _EVAL_57 = _EVAL_7 == _EVAL_176;
  assign _EVAL_31 = _EVAL_109[4:0];
  assign _EVAL_171 = ~_EVAL_117;
  assign _EVAL_152 = 5'h3 << _EVAL_11;
  assign _EVAL_100 = _EVAL_164[0];
  assign _EVAL_38 = ~_EVAL_95;
  assign _EVAL_29 = _EVAL_126 | _EVAL;
  assign _EVAL_205 = _EVAL_174 & _EVAL_158;
  assign _EVAL_223 = _EVAL_236 | _EVAL;
  assign _EVAL_216 = _EVAL_12 == 3'h7;
  assign _EVAL_111 = _EVAL_11 >= 2'h2;
  assign _EVAL_232 = ~_EVAL_1;
  assign _EVAL_99 = _EVAL_4 == 3'h5;
  assign _EVAL_101 = _EVAL_23 | _EVAL;
  assign _EVAL_37 = 2'h1 << _EVAL_175;
  assign _EVAL_87 = _EVAL_9 & _EVAL_216;
  assign _EVAL_190 = _EVAL_111 | _EVAL_49;
  assign _EVAL_121 = _EVAL_8 <= 3'h2;
  assign _EVAL_235 = _EVAL_46 | _EVAL_62;
  assign _EVAL_88 = 8'h1 << _EVAL_7;
  assign _EVAL_177 = _EVAL_173 & _EVAL_96;
  assign _EVAL_110 = _EVAL_178 & _EVAL_156;
  assign _EVAL_193 = ~_EVAL_114;
  assign _EVAL_189 = ~_EVAL_165;
  assign _EVAL_71 = ~_EVAL_68;
  assign _EVAL_115 = _EVAL_10 & _EVAL_193;
  assign _EVAL_50 = _EVAL_8 == _EVAL_224;
  assign _EVAL_132 = ~_EVAL_231;
  assign _EVAL_186 = ~_EVAL_94;
  assign _EVAL_95 = _EVAL_93 | _EVAL;
  assign _EVAL_104 = _EVAL_129 | _EVAL;
  assign _EVAL_141 = _EVAL_12 == 3'h1;
  assign _EVAL_239 = _EVAL_208 | _EVAL_110;
  assign _EVAL_85 = _EVAL_8 == 3'h0;
  assign _EVAL_114 = {_EVAL_219,_EVAL_239,_EVAL_220,_EVAL_133};
  assign _EVAL_150 = ~_EVAL;
  assign _EVAL_98 = ~_EVAL_64;
  assign _EVAL_109 = _EVAL_202 ? _EVAL_88 : 8'h0;
  assign _EVAL_126 = _EVAL_14 == _EVAL_194;
  assign _EVAL_133 = _EVAL_190 | _EVAL_161;
  assign _EVAL_24 = _EVAL_232 | _EVAL;
  assign _EVAL_106 = ~_EVAL_10;
  assign _EVAL_63 = _EVAL_0 & _EVAL_99;
  assign _EVAL_25 = _EVAL_28[0];
  assign _EVAL_218 = _EVAL_85 | _EVAL;
  assign _EVAL_59 = _EVAL_207 + 32'h1;
  assign _EVAL_172 = _EVAL_210 & _EVAL_155;
  assign _EVAL_76 = _EVAL_106 == 4'h0;
  assign _EVAL_138 = _EVAL_2 == _EVAL_153;
  assign _EVAL_230 = _EVAL_115 == 4'h0;
  assign _EVAL_157 = _EVAL_80 >> _EVAL_7;
  assign _EVAL_30 = ~_EVAL_34;
  assign _EVAL_61 = _EVAL_80 | _EVAL_31;
  assign _EVAL_131 = _EVAL_80 != 5'h0;
  assign _EVAL_178 = _EVAL_241[0];
  assign _EVAL_202 = _EVAL_174 & _EVAL_123;
  assign _EVAL_220 = _EVAL_190 | _EVAL_16;
  assign _EVAL_54 = ~_EVAL_240;
  assign _EVAL_184 = _EVAL_12 == 3'h4;
  assign _EVAL_35 = ~_EVAL_182;
  assign _EVAL_19 = ~_EVAL_158;
  assign _EVAL_175 = _EVAL_11[0];
  assign _EVAL_128 = _EVAL_18 | _EVAL;
  assign _EVAL_48 = ~_EVAL_17;
  assign _EVAL_145 = ~_EVAL_104;
  assign _EVAL_77 = _EVAL_0 & _EVAL_213;
  assign _EVAL_82 = ~_EVAL_24;
  assign _EVAL_15 = _EVAL_84 >> _EVAL_2;
  assign _EVAL_102 = _EVAL_9 & _EVAL_237;
  assign _EVAL_241 = _EVAL_37 | 2'h1;
  assign _EVAL_40 = _EVAL_227 | _EVAL;
  assign _EVAL_200 = _EVAL_5 & _EVAL_180;
  assign _EVAL_120 = ~_EVAL_136;
  assign _EVAL_158 = ~_EVAL_170;
  assign _EVAL_67 = ~_EVAL_183;
  assign _EVAL_18 = _EVAL_10 == _EVAL_114;
  assign _EVAL_166 = ~_EVAL_179;
  assign _EVAL_58 = ~_EVAL_196;
  assign _EVAL_143 = _EVAL_9 & _EVAL_228;
  assign _EVAL_129 = _EVAL_108 | _EVAL_71;
  assign _EVAL_83 = _EVAL_9 & _EVAL_184;
  assign _EVAL_159 = _EVAL_8 != 3'h0;
  assign _EVAL_233 = ~_EVAL_131;
  assign _EVAL_182 = _EVAL_4 == 3'h6;
  assign _EVAL_135 = _EVAL_4 == 3'h0;
  assign _EVAL_69 = _EVAL_138 | _EVAL;
  assign _EVAL_66 = _EVAL_9 & _EVAL_19;
  assign _EVAL_196 = _EVAL_76 | _EVAL;
  assign _EVAL_79 = {1'b0,$signed(_EVAL_160)};
  assign _EVAL_124 = _EVAL_222 & _EVAL_130;
  assign _EVAL_139 = _EVAL_174 | _EVAL_210;
  assign _EVAL_168 = _EVAL_9 & _EVAL_141;
  assign _EVAL_231 = _EVAL_57 | _EVAL;
  assign _EVAL_165 = _EVAL_146 | _EVAL;
  assign _EVAL_228 = _EVAL_12 == 3'h0;
  assign _EVAL_164 = _EVAL_125 - 1'h1;
  assign _EVAL_213 = ~_EVAL_187;
  assign _EVAL_222 = _EVAL_241[1];
  assign _EVAL_28 = _EVAL_21 - 1'h1;
  assign _EVAL_75 = _EVAL_235 | _EVAL;
  assign _EVAL_214 = ~_EVAL_128;
  assign _EVAL_225 = _EVAL_26 ? _EVAL_65 : 8'h0;
  assign _EVAL_105 = _EVAL_92;
  assign _EVAL_146 = _EVAL_4 <= 3'h6;
  assign _EVAL_32 = _EVAL_4 == 3'h2;
  assign _EVAL_97 = _EVAL_4 == _EVAL_185;
  assign _EVAL_147 = _EVAL_12 == _EVAL_162;
  assign _EVAL_49 = _EVAL_222 & _EVAL_55;
  assign _EVAL_236 = _EVAL_14 >= 2'h2;
  assign _EVAL_237 = _EVAL_12 == 3'h3;
  assign _EVAL_55 = ~_EVAL_130;
  assign _EVAL_122 = _EVAL_9 & _EVAL_45;
  assign _EVAL_211 = _EVAL_0 & _EVAL_142;
  assign _EVAL_116 = _EVAL_9 & _EVAL_226;
  assign _EVAL_118 = _EVAL_4 == 3'h4;
  assign _EVAL_65 = 8'h1 << _EVAL_2;
  assign _EVAL_167 = ~_EVAL_29;
  assign _EVAL_44 = _EVAL_8 <= 3'h4;
  assign _EVAL_179 = _EVAL_97 | _EVAL;
  assign _EVAL_20 = _EVAL_9 & _EVAL_22;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_21 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_78 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_80 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_125 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_153 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_162 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_170 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_176 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_185 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_194 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_207 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_217 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_221 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_224 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_6) begin
    if (_EVAL) begin
      _EVAL_21 <= 1'h0;
    end else if (_EVAL_210) begin
      if (_EVAL_155) begin
        _EVAL_21 <= 1'h0;
      end else begin
        _EVAL_21 <= _EVAL_25;
      end
    end
    if (_EVAL_205) begin
      _EVAL_78 <= _EVAL_11;
    end
    if (_EVAL) begin
      _EVAL_80 <= 5'h0;
    end else begin
      _EVAL_80 <= _EVAL_204;
    end
    if (_EVAL) begin
      _EVAL_125 <= 1'h0;
    end else if (_EVAL_174) begin
      if (_EVAL_123) begin
        _EVAL_125 <= 1'h0;
      end else begin
        _EVAL_125 <= _EVAL_100;
      end
    end
    if (_EVAL_103) begin
      _EVAL_153 <= _EVAL_2;
    end
    if (_EVAL_205) begin
      _EVAL_162 <= _EVAL_12;
    end
    if (_EVAL) begin
      _EVAL_170 <= 1'h0;
    end else if (_EVAL_174) begin
      if (_EVAL_158) begin
        _EVAL_170 <= 1'h0;
      end else begin
        _EVAL_170 <= _EVAL_238;
      end
    end
    if (_EVAL_205) begin
      _EVAL_176 <= _EVAL_7;
    end
    if (_EVAL_103) begin
      _EVAL_185 <= _EVAL_4;
    end
    if (_EVAL_103) begin
      _EVAL_194 <= _EVAL_14;
    end
    if (_EVAL) begin
      _EVAL_207 <= 32'h0;
    end else if (_EVAL_139) begin
      _EVAL_207 <= 32'h0;
    end else begin
      _EVAL_207 <= _EVAL_42;
    end
    if (_EVAL) begin
      _EVAL_217 <= 1'h0;
    end else if (_EVAL_210) begin
      if (_EVAL_187) begin
        _EVAL_217 <= 1'h0;
      end else begin
        _EVAL_217 <= _EVAL_91;
      end
    end
    if (_EVAL_205) begin
      _EVAL_221 <= _EVAL_5;
    end
    if (_EVAL_205) begin
      _EVAL_224 <= _EVAL_8;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(900fca35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5c490ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(719ec368)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16db8ef4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4144783a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c096dfd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3858f8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11005592)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74f24815)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a6a7cf8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d31429d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba1b75e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccf1561b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(655caa4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f20b596)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8cdd93f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acd6be12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcbce7ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(694b3aa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a440d73b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(614c2c58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6e37d56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7ddbad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3fa20ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(487a0621)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e8999da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f50de34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fe223f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56818047)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c444832)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc535e0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74ea9711)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(310649e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca7c1036)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef3e3366)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(766ca263)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12c23952)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89b2bbb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f5c9cc7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81d432d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31668ac4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57bf4dbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73eeb965)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32b4781e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd91cd68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1cb998a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99542aca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27398fe2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed4d2b11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cc28306)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(840dc32e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d63897cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87e983f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8eaf14a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f77a0b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3abde3a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa1ec43a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbee73ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7bc5bce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c07a360c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fab3db20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23af42bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6940c86b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ae8322f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(428b0ef7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1971cb10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd5e1c9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84ef941b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86076fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6540d3e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8742a04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dddfc867)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(205447f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
