//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_173_assert(
  input         _EVAL,
  input  [3:0]  _EVAL_0,
  input  [1:0]  _EVAL_1,
  input  [1:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [31:0] _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [2:0]  _EVAL_13,
  input  [2:0]  _EVAL_14
);
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire [7:0] _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire [31:0] plusarg_reader_out;
  wire [4:0] _EVAL_26;
  wire  _EVAL_27;
  wire [1:0] _EVAL_28;
  wire  _EVAL_29;
  reg [31:0] _EVAL_31;
  reg [31:0] _RAND_0;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire [1:0] _EVAL_34;
  wire  _EVAL_35;
  reg [1:0] _EVAL_36;
  reg [31:0] _RAND_1;
  wire  _EVAL_37;
  reg [4:0] _EVAL_38;
  reg [31:0] _RAND_2;
  wire [1:0] _EVAL_39;
  wire [1:0] _EVAL_40;
  wire  _EVAL_42;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire [7:0] _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  reg [31:0] _EVAL_56;
  reg [31:0] _RAND_3;
  wire  _EVAL_57;
  wire [4:0] _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  reg [2:0] _EVAL_61;
  reg [31:0] _RAND_4;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire [7:0] _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire [7:0] _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire [1:0] _EVAL_100;
  wire  _EVAL_101;
  wire [1:0] _EVAL_102;
  wire  _EVAL_103;
  wire [3:0] _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire [32:0] _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire [1:0] _EVAL_114;
  wire  _EVAL_115;
  wire [32:0] _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  reg  _EVAL_119;
  reg [31:0] _RAND_5;
  wire [4:0] _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire [32:0] _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  reg  _EVAL_144;
  reg [31:0] _RAND_6;
  wire  _EVAL_145;
  wire  _EVAL_146;
  reg  _EVAL_147;
  reg [31:0] _RAND_7;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire [3:0] _EVAL_151;
  wire [31:0] _EVAL_152;
  wire  _EVAL_153;
  wire [31:0] _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire [31:0] _EVAL_160;
  wire  _EVAL_161;
  wire [1:0] _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire [3:0] _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [4:0] _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire [4:0] _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire [32:0] _EVAL_195;
  wire  _EVAL_196;
  wire [4:0] _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  reg [2:0] _EVAL_201;
  reg [31:0] _RAND_8;
  wire [4:0] _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  reg  _EVAL_207;
  reg [31:0] _RAND_9;
  wire  _EVAL_208;
  wire  _EVAL_209;
  reg [2:0] _EVAL_210;
  reg [31:0] _RAND_10;
  reg [2:0] _EVAL_211;
  reg [31:0] _RAND_11;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  reg [2:0] _EVAL_215;
  reg [31:0] _RAND_12;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  reg [1:0] _EVAL_221;
  reg [31:0] _RAND_13;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire [31:0] _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire [4:0] _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire [3:0] _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire [4:0] _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_208 = _EVAL_14 == 3'h0;
  assign _EVAL_194 = _EVAL_139 | _EVAL_85;
  assign _EVAL_199 = _EVAL_165 & _EVAL_196;
  assign _EVAL_185 = _EVAL_58 != _EVAL_239;
  assign _EVAL_166 = _EVAL_1 >= 2'h2;
  assign _EVAL_100 = _EVAL_207 - 1'h1;
  assign _EVAL_136 = _EVAL_9 & _EVAL_21;
  assign _EVAL_200 = ~_EVAL_147;
  assign _EVAL_192 = _EVAL_140 | _EVAL_6;
  assign _EVAL_222 = ~_EVAL_99;
  assign _EVAL_97 = _EVAL_166 | _EVAL_6;
  assign _EVAL_229 = ~_EVAL_142;
  assign _EVAL_234 = _EVAL_12 == 3'h7;
  assign _EVAL_109 = $signed(_EVAL_123) & -33'sh4000;
  assign _EVAL_88 = ~_EVAL_130;
  assign _EVAL_226 = _EVAL_8 & _EVAL_154;
  assign _EVAL_65 = _EVAL_11 <= 3'h3;
  assign _EVAL_46 = _EVAL_10 & _EVAL_110;
  assign _EVAL_150 = _EVAL_7 <= 3'h4;
  assign _EVAL_19 = _EVAL_129 ? _EVAL_53 : 8'h0;
  assign _EVAL_165 = _EVAL_3 & _EVAL_10;
  assign _EVAL_187 = _EVAL_38 >> _EVAL_13;
  assign _EVAL_51 = ~_EVAL_52;
  assign _EVAL_103 = _EVAL_8[0];
  assign _EVAL_139 = ~_EVAL_180;
  assign _EVAL_209 = _EVAL_179 & _EVAL_103;
  assign _EVAL_57 = _EVAL_188 & _EVAL_103;
  assign _EVAL_129 = _EVAL_165 & _EVAL_198;
  assign _EVAL_78 = _EVAL_68 | _EVAL_108;
  assign _EVAL_130 = _EVAL_137 | _EVAL_6;
  assign _EVAL_113 = _EVAL_9 & _EVAL_208;
  assign _EVAL_232 = _EVAL_9 & _EVAL_75;
  assign _EVAL_89 = ~_EVAL_71;
  assign _EVAL_117 = _EVAL_9 & _EVAL_241;
  assign _EVAL_133 = _EVAL_9 & _EVAL_55;
  assign _EVAL_135 = _EVAL_115 & _EVAL_84;
  assign _EVAL_87 = _EVAL_11 <= 3'h1;
  assign _EVAL_121 = _EVAL_187[0];
  assign _EVAL_74 = ~_EVAL_103;
  assign _EVAL_155 = ~_EVAL_193;
  assign _EVAL_101 = _EVAL_204 & _EVAL_188;
  assign _EVAL_151 = ~_EVAL_0;
  assign _EVAL_241 = ~_EVAL_200;
  assign _EVAL_79 = _EVAL_10 & _EVAL_234;
  assign _EVAL_188 = ~_EVAL_179;
  assign _EVAL_131 = _EVAL_0 == _EVAL_104;
  assign _EVAL_112 = _EVAL_134 | _EVAL_6;
  assign _EVAL_145 = _EVAL_14 == _EVAL_215;
  assign _EVAL_143 = _EVAL_10 & _EVAL_124;
  assign _EVAL_198 = ~_EVAL_207;
  assign _EVAL_45 = _EVAL_141 | _EVAL_135;
  assign _EVAL_163 = _EVAL_147 - 1'h1;
  assign _EVAL_202 = _EVAL_120 & _EVAL_174;
  assign _EVAL_92 = _EVAL_10 & _EVAL_181;
  assign _EVAL_167 = _EVAL_141 | _EVAL_54;
  assign _EVAL_204 = _EVAL_34[1];
  assign _EVAL_240 = _EVAL_114[0];
  assign _EVAL_180 = _EVAL_38 != 5'h0;
  assign _EVAL_80 = 8'h1 << _EVAL_7;
  assign _EVAL_236 = _EVAL_0 & _EVAL_170;
  assign _EVAL_182 = _EVAL_188 & _EVAL_74;
  assign _EVAL_26 = _EVAL_197 >> _EVAL_7;
  assign _EVAL_153 = ~_EVAL_138;
  assign _EVAL_217 = _EVAL_27 | _EVAL_6;
  assign _EVAL_83 = _EVAL_13 <= 3'h4;
  assign _EVAL_193 = _EVAL_58 != 5'h0;
  assign _EVAL_195 = _EVAL_31 + 32'h1;
  assign _EVAL_23 = _EVAL_2 == _EVAL_36;
  assign _EVAL_32 = _EVAL_14 == 3'h1;
  assign _EVAL_168 = _EVAL_118 | _EVAL_6;
  assign _EVAL_16 = _EVAL_1 == _EVAL_221;
  assign _EVAL_60 = _EVAL_39[0];
  assign _EVAL_225 = _EVAL_185 | _EVAL_155;
  assign _EVAL_29 = _EVAL_164 | _EVAL_6;
  assign _EVAL_93 = ~_EVAL_4;
  assign _EVAL_17 = _EVAL_235 | _EVAL_6;
  assign _EVAL_138 = _EVAL_87 | _EVAL_6;
  assign _EVAL_15 = _EVAL_126 | _EVAL_6;
  assign _EVAL_27 = _EVAL_236 == 4'h0;
  assign _EVAL_18 = ~_EVAL_203;
  assign _EVAL_148 = _EVAL_14 == 3'h5;
  assign _EVAL_191 = _EVAL_63 & _EVAL_59;
  assign _EVAL_230 = _EVAL_12 == 3'h0;
  assign _EVAL_54 = _EVAL_115 & _EVAL_209;
  assign _EVAL_132 = $signed(_EVAL_116) == 33'sh0;
  assign _EVAL_84 = _EVAL_179 & _EVAL_74;
  assign _EVAL_98 = _EVAL_10 & _EVAL_127;
  assign _EVAL_49 = _EVAL_150 | _EVAL_6;
  assign _EVAL_223 = _EVAL_10 & _EVAL_230;
  assign _EVAL_237 = ~_EVAL_76;
  assign _EVAL_128 = ~_EVAL_97;
  assign _EVAL_37 = _EVAL_184 | _EVAL_6;
  assign _EVAL_99 = _EVAL_23 | _EVAL_6;
  assign _EVAL_214 = _EVAL_11 != 3'h0;
  assign _EVAL_55 = _EVAL_14 == 3'h4;
  assign _EVAL_213 = ~_EVAL_35;
  assign _EVAL_149 = _EVAL_14 <= 3'h6;
  assign _EVAL_114 = _EVAL_119 - 1'h1;
  assign _EVAL_179 = _EVAL_8[1];
  assign _EVAL_39 = _EVAL_144 - 1'h1;
  assign _EVAL_196 = ~_EVAL_144;
  assign _EVAL_35 = _EVAL_65 | _EVAL_6;
  assign _EVAL_238 = ~_EVAL_121;
  assign _EVAL_63 = _EVAL_5 & _EVAL_9;
  assign _EVAL_152 = _EVAL_195[31:0];
  assign _EVAL_94 = ~_EVAL_168;
  assign _EVAL_107 = ~_EVAL_15;
  assign _EVAL_90 = ~_EVAL_96;
  assign _EVAL_86 = _EVAL_1[0];
  assign _EVAL_105 = _EVAL_12 == _EVAL_61;
  assign _EVAL_123 = {1'b0,$signed(_EVAL_160)};
  assign _EVAL_124 = _EVAL_12 == 3'h6;
  assign _EVAL_44 = _EVAL_131 | _EVAL_6;
  assign _EVAL_111 = ~_EVAL_192;
  assign _EVAL_154 = {{30'd0}, _EVAL_28};
  assign _EVAL_157 = _EVAL_191 & _EVAL_228;
  assign _EVAL_20 = _EVAL_10 & _EVAL_218;
  assign _EVAL_231 = 5'h3 << _EVAL_1;
  assign _EVAL_53 = 8'h1 << _EVAL_13;
  assign _EVAL_67 = _EVAL_157 ? _EVAL_80 : 8'h0;
  assign _EVAL_91 = ~_EVAL_44;
  assign _EVAL_239 = _EVAL_67[4:0];
  assign _EVAL_156 = _EVAL_163[0];
  assign _EVAL_172 = _EVAL_178 | _EVAL_6;
  assign _EVAL_102 = _EVAL_231[1:0];
  assign _EVAL_85 = plusarg_reader_out == 32'h0;
  assign _EVAL_95 = _EVAL_149 | _EVAL_6;
  assign _EVAL_126 = _EVAL_11 == 3'h0;
  assign _EVAL_76 = _EVAL_238 | _EVAL_6;
  assign _EVAL_227 = _EVAL_63 & _EVAL_200;
  assign _EVAL_81 = _EVAL_115 & _EVAL_57;
  assign _EVAL_233 = ~_EVAL_37;
  assign _EVAL_75 = _EVAL_14 == 3'h2;
  assign _EVAL_106 = _EVAL_204 & _EVAL_179;
  assign _EVAL_160 = _EVAL_8 ^ 32'h80008000;
  assign _EVAL_169 = ~_EVAL_17;
  assign _EVAL_47 = ~_EVAL_186;
  assign _EVAL_104 = {_EVAL_167,_EVAL_45,_EVAL_219,_EVAL_78};
  assign _EVAL_218 = _EVAL_12 == 3'h4;
  assign _EVAL_66 = ~_EVAL_205;
  assign _EVAL_228 = ~_EVAL_21;
  assign _EVAL_96 = _EVAL_77 | _EVAL_6;
  assign _EVAL_42 = _EVAL_165 | _EVAL_63;
  assign _EVAL_159 = ~_EVAL_112;
  assign _EVAL_118 = _EVAL_11 == _EVAL_210;
  assign _EVAL_170 = ~_EVAL_104;
  assign _EVAL_34 = _EVAL_40 | 2'h1;
  assign _EVAL_216 = ~_EVAL_176;
  assign _EVAL_164 = _EVAL_11 <= 3'h2;
  assign _EVAL_186 = _EVAL_225 | _EVAL_6;
  assign _EVAL_184 = _EVAL_72 & _EVAL_132;
  assign _EVAL_134 = _EVAL_7 == _EVAL_201;
  assign _EVAL_178 = _EVAL_11 <= 3'h4;
  assign _EVAL_142 = _EVAL_105 | _EVAL_6;
  assign _EVAL_82 = _EVAL_100[0];
  assign _EVAL_137 = _EVAL_8 == _EVAL_56;
  assign _EVAL_212 = ~_EVAL_24;
  assign _EVAL_116 = _EVAL_109;
  assign _EVAL_171 = ~_EVAL_62;
  assign _EVAL_189 = _EVAL_2 >= 2'h2;
  assign _EVAL_71 = _EVAL_83 | _EVAL_6;
  assign _EVAL_110 = ~_EVAL_196;
  assign _EVAL_70 = _EVAL_151 == 4'h0;
  assign _EVAL_173 = _EVAL_10 & _EVAL_50;
  assign _EVAL_21 = _EVAL_14 == 3'h6;
  assign _EVAL_205 = _EVAL_161 | _EVAL_6;
  assign _EVAL_197 = _EVAL_58 | _EVAL_38;
  assign _EVAL_24 = _EVAL_189 | _EVAL_6;
  assign _EVAL_206 = ~_EVAL_190;
  assign _EVAL_120 = _EVAL_38 | _EVAL_58;
  assign _EVAL_235 = _EVAL_26[0];
  assign _EVAL_125 = ~_EVAL_6;
  assign _EVAL_50 = _EVAL_12 == 3'h5;
  assign _EVAL_33 = _EVAL_9 & _EVAL_32;
  assign _EVAL_77 = _EVAL_226 == 32'h0;
  assign _EVAL_72 = _EVAL_1 <= 2'h2;
  assign _EVAL_219 = _EVAL_68 | _EVAL_81;
  assign _EVAL_220 = _EVAL_12 == 3'h3;
  assign _EVAL_28 = ~_EVAL_102;
  assign _EVAL_203 = _EVAL_145 | _EVAL_6;
  assign _EVAL_140 = _EVAL_13 == _EVAL_211;
  assign _EVAL_190 = _EVAL_214 | _EVAL_6;
  assign _EVAL_68 = _EVAL_166 | _EVAL_101;
  assign _EVAL_108 = _EVAL_115 & _EVAL_182;
  assign _EVAL_177 = _EVAL_31 < plusarg_reader_out;
  assign _EVAL_176 = _EVAL_93 | _EVAL_6;
  assign _EVAL_40 = 2'h1 << _EVAL_86;
  assign _EVAL_181 = _EVAL_12 == 3'h1;
  assign _EVAL_127 = _EVAL_12 == 3'h2;
  assign _EVAL_175 = _EVAL_10 & _EVAL_220;
  assign _EVAL_59 = ~_EVAL_119;
  assign _EVAL_64 = ~_EVAL_172;
  assign _EVAL_224 = ~_EVAL_95;
  assign _EVAL_69 = ~_EVAL_49;
  assign _EVAL_58 = _EVAL_19[4:0];
  assign _EVAL_174 = ~_EVAL_239;
  assign _EVAL_146 = ~_EVAL_217;
  assign _EVAL_52 = _EVAL_16 | _EVAL_6;
  assign _EVAL_115 = _EVAL_34[0];
  assign _EVAL_161 = _EVAL_194 | _EVAL_177;
  assign _EVAL_158 = ~_EVAL_29;
  assign _EVAL_122 = _EVAL_9 & _EVAL_148;
  assign _EVAL_141 = _EVAL_166 | _EVAL_106;
  assign _EVAL_62 = _EVAL_70 | _EVAL_6;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_31 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_36 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_38 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_56 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_61 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_119 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_144 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_147 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_201 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_207 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_210 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_211 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_215 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_221 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL) begin
    if (_EVAL_6) begin
      _EVAL_31 <= 32'h0;
    end else if (_EVAL_42) begin
      _EVAL_31 <= 32'h0;
    end else begin
      _EVAL_31 <= _EVAL_152;
    end
    if (_EVAL_227) begin
      _EVAL_36 <= _EVAL_2;
    end
    if (_EVAL_6) begin
      _EVAL_38 <= 5'h0;
    end else begin
      _EVAL_38 <= _EVAL_202;
    end
    if (_EVAL_199) begin
      _EVAL_56 <= _EVAL_8;
    end
    if (_EVAL_199) begin
      _EVAL_61 <= _EVAL_12;
    end
    if (_EVAL_6) begin
      _EVAL_119 <= 1'h0;
    end else if (_EVAL_63) begin
      if (_EVAL_59) begin
        _EVAL_119 <= 1'h0;
      end else begin
        _EVAL_119 <= _EVAL_240;
      end
    end
    if (_EVAL_6) begin
      _EVAL_144 <= 1'h0;
    end else if (_EVAL_165) begin
      if (_EVAL_196) begin
        _EVAL_144 <= 1'h0;
      end else begin
        _EVAL_144 <= _EVAL_60;
      end
    end
    if (_EVAL_6) begin
      _EVAL_147 <= 1'h0;
    end else if (_EVAL_63) begin
      if (_EVAL_200) begin
        _EVAL_147 <= 1'h0;
      end else begin
        _EVAL_147 <= _EVAL_156;
      end
    end
    if (_EVAL_227) begin
      _EVAL_201 <= _EVAL_7;
    end
    if (_EVAL_6) begin
      _EVAL_207 <= 1'h0;
    end else if (_EVAL_165) begin
      if (_EVAL_198) begin
        _EVAL_207 <= 1'h0;
      end else begin
        _EVAL_207 <= _EVAL_82;
      end
    end
    if (_EVAL_199) begin
      _EVAL_210 <= _EVAL_11;
    end
    if (_EVAL_199) begin
      _EVAL_211 <= _EVAL_13;
    end
    if (_EVAL_227) begin
      _EVAL_215 <= _EVAL_14;
    end
    if (_EVAL_199) begin
      _EVAL_221 <= _EVAL_1;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9113b407)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f153b933)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(531165f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8597974)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92cef5d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62eed0c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e66a53d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(781a99a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb37614c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(209fe8e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b3e5b7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc494ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78e6c073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1a4c508)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8a85551)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7e138bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f723c44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28121978)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25cd420f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78aaf8e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(616a730b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f00fc8dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fded497)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31c50a9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6a7b77a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48b8e9df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d75f6d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a735556)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27ffe693)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(503bd64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1be3f668)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df275cb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(928493d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea9e0e51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa4ecc49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a307cb1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e98919b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e54899f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1df7baef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dcbc300)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9432dfc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef800dd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea510d66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2604eba2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abbdbe1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(288f7fe0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(151db744)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(809a9c60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fa40640)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d70a4bf0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d97fde5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7f38a3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50b3dba2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24bbc2e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a88941c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(588ee2fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84d0092a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bd11c33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d296070e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(832a2f23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(161a701e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef72ccf1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae542bd9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9f56510)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61ff4225)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c661c3ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b04a078a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4d3bbf0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e797217)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2f1b03f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26ba438d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b50cd0a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d4d2e22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
