//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_77_assert(
  input  [1:0]  _EVAL,
  input         _EVAL_0,
  input  [25:0] _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [1:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [3:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [2:0]  _EVAL_13,
  input         _EVAL_14
);
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire [26:0] _EVAL_20;
  wire [1:0] _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire [1:0] _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire [7:0] _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire [26:0] _EVAL_44;
  wire [1:0] _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire [4:0] _EVAL_48;
  wire [4:0] _EVAL_49;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_55;
  reg [2:0] _EVAL_56;
  reg [31:0] _RAND_0;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  reg [1:0] _EVAL_68;
  reg [31:0] _RAND_1;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire [31:0] _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  reg [1:0] _EVAL_79;
  reg [31:0] _RAND_2;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire [1:0] _EVAL_85;
  wire [4:0] _EVAL_86;
  reg  _EVAL_87;
  reg [31:0] _RAND_3;
  reg  _EVAL_88;
  reg [31:0] _RAND_4;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  reg [31:0] _EVAL_95;
  reg [31:0] _RAND_5;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire [4:0] _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire [25:0] _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  reg [2:0] _EVAL_113;
  reg [31:0] _RAND_6;
  wire [3:0] _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  reg  _EVAL_119;
  reg [31:0] _RAND_7;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire [7:0] _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire [4:0] _EVAL_131;
  wire [7:0] _EVAL_132;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  reg [2:0] _EVAL_138;
  reg [31:0] _RAND_8;
  wire  _EVAL_140;
  wire  _EVAL_141;
  reg [4:0] _EVAL_143;
  reg [31:0] _RAND_9;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire [25:0] _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire [3:0] _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire [1:0] _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire [26:0] _EVAL_161;
  wire  _EVAL_162;
  reg [2:0] _EVAL_163;
  reg [31:0] _RAND_10;
  wire [1:0] _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire [3:0] _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire [32:0] _EVAL_175;
  wire  _EVAL_177;
  wire  _EVAL_178;
  reg  _EVAL_180;
  reg [31:0] _RAND_11;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire [25:0] _EVAL_183;
  wire  _EVAL_184;
  wire [4:0] _EVAL_185;
  wire  _EVAL_186;
  wire [3:0] _EVAL_187;
  wire [4:0] _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire [1:0] _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire [1:0] _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  reg [25:0] _EVAL_210;
  reg [31:0] _RAND_12;
  wire [4:0] _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  reg [2:0] _EVAL_226;
  reg [31:0] _RAND_13;
  wire  _EVAL_229;
  wire [7:0] _EVAL_230;
  wire [1:0] _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire [4:0] _EVAL_243;
  wire  _EVAL_244;
  wire [1:0] _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_174 = _EVAL_98 & _EVAL_39;
  assign _EVAL_202 = _EVAL_3 == 3'h7;
  assign _EVAL_204 = _EVAL_2 == 3'h4;
  assign _EVAL_125 = _EVAL_107 ? _EVAL_38 : 8'h0;
  assign _EVAL_188 = 5'h3 << _EVAL_4;
  assign _EVAL_146 = _EVAL_5 & _EVAL_11;
  assign _EVAL_107 = _EVAL_146 & _EVAL_83;
  assign _EVAL_171 = _EVAL_43 | _EVAL_6;
  assign _EVAL_109 = _EVAL_134 | _EVAL_6;
  assign _EVAL_75 = _EVAL_11 & _EVAL_156;
  assign _EVAL_43 = ~_EVAL_239;
  assign _EVAL_47 = _EVAL_164 == 2'h0;
  assign _EVAL_192 = _EVAL_200 & _EVAL_59;
  assign _EVAL_26 = 2'h1 << _EVAL_128;
  assign _EVAL_121 = _EVAL_220 & _EVAL_192;
  assign _EVAL_126 = _EVAL_117 | _EVAL_6;
  assign _EVAL_23 = _EVAL_9 & _EVAL_215;
  assign _EVAL_31 = _EVAL_13 == 3'h4;
  assign _EVAL_209 = ~_EVAL_80;
  assign _EVAL_154 = _EVAL_11 & _EVAL_72;
  assign _EVAL_251 = _EVAL_12 == _EVAL_226;
  assign _EVAL_38 = 8'h1 << _EVAL_10;
  assign _EVAL_220 = _EVAL_45[0];
  assign _EVAL_61 = _EVAL_231[0];
  assign _EVAL_244 = _EVAL_157[0];
  assign _EVAL_53 = _EVAL_18 | _EVAL_6;
  assign _EVAL_149 = ~_EVAL_224;
  assign _EVAL_20 = _EVAL_44;
  assign _EVAL_248 = _EVAL_136 | _EVAL_6;
  assign _EVAL_93 = _EVAL_247 | _EVAL_6;
  assign _EVAL_198 = _EVAL_45[1];
  assign _EVAL_224 = _EVAL_160 | _EVAL_6;
  assign _EVAL_110 = ~_EVAL_59;
  assign _EVAL_25 = _EVAL_40 | _EVAL_6;
  assign _EVAL_90 = ~_EVAL_93;
  assign _EVAL_62 = ~_EVAL_63;
  assign _EVAL_232 = ~_EVAL_34;
  assign _EVAL_46 = _EVAL_9 & _EVAL_189;
  assign _EVAL_48 = _EVAL_211 >> _EVAL_13;
  assign _EVAL_106 = _EVAL_1 ^ 26'h2000000;
  assign _EVAL_101 = _EVAL_2 == 3'h1;
  assign _EVAL_117 = _EVAL_12 != 3'h0;
  assign _EVAL_225 = _EVAL_199 == 2'h1;
  assign _EVAL_240 = _EVAL_11 & _EVAL_202;
  assign _EVAL_30 = ~_EVAL_25;
  assign _EVAL_181 = _EVAL_10 == 3'h4;
  assign _EVAL_127 = _EVAL_2 == 3'h6;
  assign _EVAL_41 = _EVAL_76 | _EVAL_6;
  assign _EVAL_114 = ~_EVAL_7;
  assign _EVAL_153 = _EVAL_35 | _EVAL_130;
  assign _EVAL_170 = _EVAL_82 | _EVAL_6;
  assign _EVAL_250 = _EVAL_64 | _EVAL_6;
  assign _EVAL_111 = ~_EVAL_104;
  assign _EVAL_28 = _EVAL_3 == 3'h6;
  assign _EVAL_70 = _EVAL_9 & _EVAL_124;
  assign _EVAL_45 = _EVAL_26 | 2'h1;
  assign _EVAL_131 = _EVAL_230[4:0];
  assign _EVAL_246 = _EVAL_178 | _EVAL_6;
  assign _EVAL_128 = _EVAL_4[0];
  assign _EVAL_124 = _EVAL_2 == 3'h0;
  assign _EVAL_185 = ~_EVAL_131;
  assign _EVAL_112 = ~_EVAL_200;
  assign _EVAL_76 = _EVAL == _EVAL_79;
  assign _EVAL_187 = {_EVAL_94,_EVAL_221,_EVAL_135,_EVAL_105};
  assign _EVAL_37 = ~_EVAL_89;
  assign _EVAL_64 = _EVAL_1 == _EVAL_210;
  assign _EVAL_196 = ~_EVAL_126;
  assign _EVAL_63 = _EVAL_100 | _EVAL_6;
  assign _EVAL_51 = _EVAL_11 & _EVAL_249;
  assign _EVAL_67 = _EVAL_122 & _EVAL_169;
  assign _EVAL_212 = ~_EVAL_119;
  assign _EVAL_231 = _EVAL_88 - 1'h1;
  assign _EVAL_97 = _EVAL_9 & _EVAL_204;
  assign _EVAL_169 = $signed(_EVAL_20) == 27'sh0;
  assign _EVAL_186 = _EVAL_67 | _EVAL_6;
  assign _EVAL_217 = _EVAL_98 & _EVAL_212;
  assign _EVAL_161 = {1'b0,$signed(_EVAL_106)};
  assign _EVAL_105 = _EVAL_223 | _EVAL_15;
  assign _EVAL_85 = ~_EVAL_193;
  assign _EVAL_18 = _EVAL_129 | _EVAL_181;
  assign _EVAL_208 = ~_EVAL_184;
  assign _EVAL_108 = ~_EVAL_246;
  assign _EVAL_77 = _EVAL_95 < plusarg_reader_out;
  assign _EVAL_140 = _EVAL_199 == 2'h0;
  assign _EVAL_152 = _EVAL_112 & _EVAL_59;
  assign _EVAL_249 = _EVAL_3 == 3'h2;
  assign _EVAL_98 = _EVAL_14 & _EVAL_9;
  assign _EVAL_118 = _EVAL_21[0];
  assign _EVAL_159 = ~_EVAL_214;
  assign _EVAL_100 = _EVAL_137 | _EVAL_77;
  assign _EVAL_177 = _EVAL_12 <= 3'h4;
  assign _EVAL_178 = _EVAL_10 == _EVAL_163;
  assign _EVAL_213 = _EVAL_225 | _EVAL_140;
  assign _EVAL_211 = _EVAL_243 | _EVAL_143;
  assign _EVAL_33 = ~_EVAL_248;
  assign _EVAL_123 = _EVAL_198 & _EVAL_112;
  assign _EVAL_83 = ~_EVAL_88;
  assign _EVAL_156 = _EVAL_3 == 3'h5;
  assign _EVAL_207 = _EVAL_55 | _EVAL_6;
  assign _EVAL_233 = _EVAL_16 | _EVAL_6;
  assign _EVAL_173 = _EVAL_7 == _EVAL_187;
  assign _EVAL_71 = _EVAL_3 == 3'h0;
  assign _EVAL_94 = _EVAL_78 | _EVAL_121;
  assign _EVAL_191 = ~_EVAL_158;
  assign _EVAL_218 = _EVAL_3 == 3'h3;
  assign _EVAL_205 = _EVAL_3 == _EVAL_113;
  assign _EVAL_92 = ~_EVAL_53;
  assign _EVAL_50 = ~_EVAL_250;
  assign _EVAL_148 = plusarg_reader_out == 32'h0;
  assign _EVAL_167 = _EVAL_245[0];
  assign _EVAL_59 = _EVAL_1[0];
  assign _EVAL_182 = _EVAL_220 & _EVAL_152;
  assign _EVAL_194 = ~_EVAL_39;
  assign _EVAL_130 = ~_EVAL_229;
  assign _EVAL_40 = _EVAL_4 >= 2'h2;
  assign _EVAL_162 = _EVAL_2 == _EVAL_138;
  assign _EVAL_19 = _EVAL_13 == _EVAL_56;
  assign _EVAL_157 = _EVAL_180 - 1'h1;
  assign _EVAL_145 = ~_EVAL_127;
  assign _EVAL_72 = ~_EVAL_165;
  assign _EVAL_22 = ~_EVAL_60;
  assign _EVAL_147 = _EVAL_1 & _EVAL_183;
  assign _EVAL_229 = _EVAL_243 != 5'h0;
  assign _EVAL_27 = _EVAL_11 & _EVAL_218;
  assign _EVAL_66 = _EVAL_3 == 3'h4;
  assign _EVAL_29 = _EVAL_9 & _EVAL_101;
  assign _EVAL_73 = _EVAL_175[31:0];
  assign _EVAL_24 = ~_EVAL_41;
  assign _EVAL_243 = _EVAL_125[4:0];
  assign _EVAL_197 = _EVAL_11 & _EVAL_71;
  assign _EVAL_49 = _EVAL_86 & _EVAL_185;
  assign _EVAL_120 = ~_EVAL_6;
  assign _EVAL_237 = ~_EVAL_207;
  assign _EVAL_17 = ~_EVAL_186;
  assign _EVAL_184 = _EVAL_177 | _EVAL_6;
  assign _EVAL_60 = _EVAL_251 | _EVAL_6;
  assign _EVAL_158 = _EVAL_236 | _EVAL_6;
  assign _EVAL_234 = _EVAL_162 | _EVAL_6;
  assign _EVAL_168 = ~_EVAL_170;
  assign _EVAL_216 = _EVAL_200 & _EVAL_110;
  assign _EVAL_144 = _EVAL_42 | _EVAL_6;
  assign _EVAL_34 = _EVAL_153 | _EVAL_6;
  assign _EVAL_150 = _EVAL_198 & _EVAL_200;
  assign _EVAL_137 = _EVAL_81 | _EVAL_148;
  assign _EVAL_89 = _EVAL_19 | _EVAL_6;
  assign _EVAL_69 = _EVAL_36 | _EVAL_6;
  assign _EVAL_236 = _EVAL_151 == 4'h0;
  assign _EVAL_215 = _EVAL_2 == 3'h2;
  assign _EVAL_172 = ~_EVAL_187;
  assign _EVAL_86 = _EVAL_143 | _EVAL_243;
  assign _EVAL_201 = _EVAL_164 == 2'h1;
  assign _EVAL_230 = _EVAL_190 ? _EVAL_132 : 8'h0;
  assign _EVAL_91 = _EVAL_173 | _EVAL_6;
  assign _EVAL_135 = _EVAL_223 | _EVAL_182;
  assign _EVAL_82 = _EVAL_12 <= 3'h3;
  assign _EVAL_42 = _EVAL_4 == _EVAL_68;
  assign _EVAL_160 = ~_EVAL_0;
  assign _EVAL_175 = _EVAL_95 + 32'h1;
  assign _EVAL_57 = _EVAL_11 & _EVAL_195;
  assign _EVAL_129 = _EVAL_201 | _EVAL_47;
  assign _EVAL_155 = _EVAL_84 | _EVAL_6;
  assign _EVAL_134 = _EVAL_48[0];
  assign _EVAL_96 = _EVAL_9 & _EVAL_127;
  assign _EVAL_222 = ~_EVAL_144;
  assign _EVAL_141 = _EVAL_12 <= 3'h2;
  assign _EVAL_102 = _EVAL_146 | _EVAL_98;
  assign _EVAL_206 = _EVAL_114 == 4'h0;
  assign _EVAL_214 = _EVAL_205 | _EVAL_6;
  assign _EVAL_65 = ~_EVAL_171;
  assign _EVAL_223 = _EVAL_40 | _EVAL_123;
  assign _EVAL_103 = _EVAL_220 & _EVAL_216;
  assign _EVAL_44 = $signed(_EVAL_161) & -27'sh1000000;
  assign _EVAL_122 = _EVAL_4 <= 2'h2;
  assign _EVAL_238 = _EVAL_9 & _EVAL_194;
  assign _EVAL_80 = _EVAL_141 | _EVAL_6;
  assign _EVAL_99 = _EVAL_143 >> _EVAL_10;
  assign _EVAL_245 = _EVAL_119 - 1'h1;
  assign _EVAL_195 = _EVAL_3 == 3'h1;
  assign _EVAL_115 = ~_EVAL_69;
  assign _EVAL_235 = ~_EVAL_234;
  assign _EVAL_221 = _EVAL_78 | _EVAL_103;
  assign _EVAL_39 = ~_EVAL_87;
  assign _EVAL_239 = _EVAL_99[0];
  assign _EVAL_104 = _EVAL_206 | _EVAL_6;
  assign _EVAL_183 = {{24'd0}, _EVAL_85};
  assign _EVAL_132 = 8'h1 << _EVAL_13;
  assign _EVAL_55 = _EVAL_2 <= 3'h6;
  assign _EVAL_151 = _EVAL_7 & _EVAL_172;
  assign _EVAL_78 = _EVAL_40 | _EVAL_150;
  assign _EVAL_200 = _EVAL_1[1];
  assign _EVAL_193 = _EVAL_188[1:0];
  assign _EVAL_35 = _EVAL_243 != _EVAL_131;
  assign _EVAL_242 = ~_EVAL_109;
  assign _EVAL_81 = ~_EVAL_166;
  assign _EVAL_116 = ~_EVAL_233;
  assign _EVAL_36 = _EVAL_12 <= 3'h1;
  assign _EVAL_32 = _EVAL_11 & _EVAL_66;
  assign _EVAL_16 = _EVAL_147 == 26'h0;
  assign _EVAL_219 = ~_EVAL_91;
  assign _EVAL_247 = _EVAL >= 2'h2;
  assign _EVAL_136 = _EVAL_213 | _EVAL_31;
  assign _EVAL_241 = ~_EVAL_155;
  assign _EVAL_74 = _EVAL_11 & _EVAL_28;
  assign _EVAL_84 = _EVAL_12 == 3'h0;
  assign _EVAL_199 = _EVAL_13[2:1];
  assign _EVAL_166 = _EVAL_143 != 5'h0;
  assign _EVAL_21 = _EVAL_87 - 1'h1;
  assign _EVAL_165 = ~_EVAL_180;
  assign _EVAL_58 = _EVAL_112 & _EVAL_110;
  assign _EVAL_189 = _EVAL_2 == 3'h5;
  assign _EVAL_52 = _EVAL_146 & _EVAL_165;
  assign _EVAL_15 = _EVAL_220 & _EVAL_58;
  assign _EVAL_190 = _EVAL_217 & _EVAL_145;
  assign _EVAL_164 = _EVAL_10[2:1];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_56 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_68 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_79 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_87 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_88 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_95 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_113 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_119 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_138 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_143 = _RAND_9[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_163 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_180 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_210 = _RAND_12[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_226 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_8) begin
    if (_EVAL_174) begin
      _EVAL_56 <= _EVAL_13;
    end
    if (_EVAL_52) begin
      _EVAL_68 <= _EVAL_4;
    end
    if (_EVAL_174) begin
      _EVAL_79 <= _EVAL;
    end
    if (_EVAL_6) begin
      _EVAL_87 <= 1'h0;
    end else if (_EVAL_98) begin
      if (_EVAL_39) begin
        _EVAL_87 <= 1'h0;
      end else begin
        _EVAL_87 <= _EVAL_118;
      end
    end
    if (_EVAL_6) begin
      _EVAL_88 <= 1'h0;
    end else if (_EVAL_146) begin
      if (_EVAL_83) begin
        _EVAL_88 <= 1'h0;
      end else begin
        _EVAL_88 <= _EVAL_61;
      end
    end
    if (_EVAL_6) begin
      _EVAL_95 <= 32'h0;
    end else if (_EVAL_102) begin
      _EVAL_95 <= 32'h0;
    end else begin
      _EVAL_95 <= _EVAL_73;
    end
    if (_EVAL_52) begin
      _EVAL_113 <= _EVAL_3;
    end
    if (_EVAL_6) begin
      _EVAL_119 <= 1'h0;
    end else if (_EVAL_98) begin
      if (_EVAL_212) begin
        _EVAL_119 <= 1'h0;
      end else begin
        _EVAL_119 <= _EVAL_167;
      end
    end
    if (_EVAL_174) begin
      _EVAL_138 <= _EVAL_2;
    end
    if (_EVAL_6) begin
      _EVAL_143 <= 5'h0;
    end else begin
      _EVAL_143 <= _EVAL_49;
    end
    if (_EVAL_52) begin
      _EVAL_163 <= _EVAL_10;
    end
    if (_EVAL_6) begin
      _EVAL_180 <= 1'h0;
    end else if (_EVAL_146) begin
      if (_EVAL_165) begin
        _EVAL_180 <= 1'h0;
      end else begin
        _EVAL_180 <= _EVAL_244;
      end
    end
    if (_EVAL_52) begin
      _EVAL_210 <= _EVAL_1;
    end
    if (_EVAL_52) begin
      _EVAL_226 <= _EVAL_12;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1101092f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1c50339)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1274980e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86d14985)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b49ef97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90762cf8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a003657)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f40266d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d210bb82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(311eee2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(658efa04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53aff583)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7564ea71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81addba4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(261e3381)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4044799d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc5e9b7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bec9dfad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fb0ef47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(496c9f8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5c4f8fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e0e474c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af80ba55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d505b27f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e032816c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2879286a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(817c67c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de733f55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eae819d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1855039)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25f864b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ed80e57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4381f4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ba925f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c595cfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85f10ada)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33c9d678)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b25ac4d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6fb9fc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ef08d03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(804d65d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33ea9b03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(782fd51b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59d9e878)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39eabb47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38883ab1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(319aa0f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e1606d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af58263d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75e8505e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e960f713)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c965720)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bafe397)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67e7cbf6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81820a56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a057deb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5efc9b35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41d19fa3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ca687c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6714076)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5fbdba2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15ed91b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24daadc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3ec247)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc6e426f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(428bbb38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77ec2df3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7702c67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(171a54dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9458019)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82e15d91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37d09dfc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ad6a323)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
