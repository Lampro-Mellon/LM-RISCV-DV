//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_92_assert(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [29:0] _EVAL_4,
  input         _EVAL_5,
  input  [3:0]  _EVAL_6,
  input         _EVAL_7,
  input  [1:0]  _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  input  [1:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input  [1:0]  _EVAL_15,
  input         _EVAL_16,
  input  [2:0]  _EVAL_17,
  input         _EVAL_18
);
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire [4:0] _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  reg [2:0] _EVAL_27;
  reg [31:0] _RAND_0;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire [1:0] _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  reg  _EVAL_34;
  reg [31:0] _RAND_1;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire [1:0] _EVAL_42;
  wire  _EVAL_43;
  reg [4:0] _EVAL_44;
  reg [31:0] _RAND_2;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire [31:0] plusarg_reader_out;
  wire [3:0] _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_53;
  reg [2:0] _EVAL_54;
  reg [31:0] _RAND_3;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire [4:0] _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  reg [29:0] _EVAL_70;
  reg [31:0] _RAND_4;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire [1:0] _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire [4:0] _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire [3:0] _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire [7:0] _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  reg [1:0] _EVAL_99;
  reg [31:0] _RAND_5;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire [1:0] _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire [32:0] _EVAL_113;
  wire [30:0] _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire [29:0] _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire [30:0] _EVAL_128;
  wire [30:0] _EVAL_129;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire [1:0] _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire [3:0] _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire [7:0] _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  reg  _EVAL_161;
  reg [31:0] _RAND_6;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire [1:0] _EVAL_172;
  wire  _EVAL_173;
  wire [1:0] _EVAL_174;
  wire [7:0] _EVAL_175;
  wire  _EVAL_176;
  reg  _EVAL_177;
  reg [31:0] _RAND_7;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  reg [2:0] _EVAL_184;
  reg [31:0] _RAND_8;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  reg  _EVAL_193;
  reg [31:0] _RAND_9;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  reg  _EVAL_197;
  reg [31:0] _RAND_10;
  wire  _EVAL_198;
  wire  _EVAL_199;
  reg [2:0] _EVAL_200;
  reg [31:0] _RAND_11;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  reg [31:0] _EVAL_211;
  reg [31:0] _RAND_12;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire [29:0] _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire [1:0] _EVAL_222;
  wire [1:0] _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  reg [1:0] _EVAL_229;
  reg [31:0] _RAND_13;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire [4:0] _EVAL_239;
  wire [3:0] _EVAL_240;
  wire  _EVAL_241;
  wire [4:0] _EVAL_242;
  wire  _EVAL_243;
  wire [29:0] _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  reg [1:0] _EVAL_253;
  reg [31:0] _RAND_14;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_259;
  wire [4:0] _EVAL_260;
  wire  _EVAL_261;
  wire [31:0] _EVAL_262;
  wire  _EVAL_263;
  wire [4:0] _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire [1:0] _EVAL_269;
  reg  _EVAL_270;
  reg [31:0] _RAND_15;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire [4:0] _EVAL_273;
  wire  _EVAL_274;
  reg [2:0] _EVAL_275;
  reg [31:0] _RAND_16;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire [4:0] _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire [7:0] _EVAL_285;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_170 = _EVAL_159 | _EVAL_168;
  assign _EVAL_203 = ~_EVAL_257;
  assign _EVAL_202 = _EVAL_143 | _EVAL_2;
  assign _EVAL_64 = _EVAL_188 | _EVAL_2;
  assign _EVAL_41 = _EVAL_42 == 2'h0;
  assign _EVAL_176 = _EVAL_86 & _EVAL_249;
  assign _EVAL_155 = _EVAL_189 | _EVAL_215;
  assign _EVAL_214 = ~_EVAL_121;
  assign _EVAL_196 = _EVAL_174 == 2'h0;
  assign _EVAL_201 = _EVAL_8 == 2'h0;
  assign _EVAL_273 = _EVAL_285[4:0];
  assign _EVAL_137 = _EVAL_8 != 2'h2;
  assign _EVAL_247 = _EVAL_13 & _EVAL_87;
  assign _EVAL_215 = _EVAL_17 == 3'h4;
  assign _EVAL_224 = _EVAL_172 | 2'h1;
  assign _EVAL_262 = _EVAL_113[31:0];
  assign _EVAL_261 = _EVAL_85 | _EVAL_2;
  assign _EVAL_145 = _EVAL_84 & _EVAL_25;
  assign _EVAL_103 = ~_EVAL_216;
  assign _EVAL_107 = _EVAL_8 <= 2'h2;
  assign _EVAL_142 = _EVAL_6 & _EVAL_240;
  assign _EVAL_237 = _EVAL_44 != 5'h0;
  assign _EVAL_147 = _EVAL_15 >= 2'h2;
  assign _EVAL_63 = plusarg_reader_out == 32'h0;
  assign _EVAL_31 = _EVAL_34 - 1'h1;
  assign _EVAL_265 = _EVAL_12 >= 2'h2;
  assign _EVAL_84 = _EVAL_15 <= 2'h2;
  assign _EVAL_206 = ~_EVAL_153;
  assign _EVAL_218 = _EVAL_190 | _EVAL_63;
  assign _EVAL_221 = _EVAL_12 == _EVAL_99;
  assign _EVAL_38 = _EVAL_10 == _EVAL_200;
  assign _EVAL_33 = ~_EVAL_2;
  assign _EVAL_28 = ~_EVAL_64;
  assign _EVAL_267 = _EVAL_224[1];
  assign _EVAL_39 = _EVAL_164 & _EVAL_167;
  assign _EVAL_59 = _EVAL_5 & _EVAL_72;
  assign _EVAL_76 = _EVAL_147 | _EVAL_179;
  assign _EVAL_241 = ~_EVAL_182;
  assign _EVAL_132 = ~_EVAL_156;
  assign _EVAL_35 = ~_EVAL_161;
  assign _EVAL_65 = _EVAL_211 < plusarg_reader_out;
  assign _EVAL_199 = ~_EVAL_20;
  assign _EVAL_278 = _EVAL_13 & _EVAL_127;
  assign _EVAL_120 = _EVAL_15[0];
  assign _EVAL_228 = ~_EVAL_53;
  assign _EVAL_256 = ~_EVAL_90;
  assign _EVAL_185 = _EVAL_66 | _EVAL_2;
  assign _EVAL_136 = ~_EVAL_45;
  assign _EVAL_102 = _EVAL_11 == 3'h6;
  assign _EVAL_244 = _EVAL_4 ^ 30'h20000000;
  assign _EVAL_105 = ~_EVAL_251;
  assign _EVAL_180 = _EVAL_69 | _EVAL_2;
  assign _EVAL_210 = _EVAL_142 == 4'h0;
  assign _EVAL_187 = _EVAL_8 == _EVAL_229;
  assign _EVAL_75 = _EVAL_3 == 3'h3;
  assign _EVAL_115 = {1'b0,$signed(_EVAL_244)};
  assign _EVAL_83 = ~_EVAL_140;
  assign _EVAL_264 = _EVAL_239 | _EVAL_44;
  assign _EVAL_43 = _EVAL_210 | _EVAL_2;
  assign _EVAL_73 = _EVAL_161 - 1'h1;
  assign _EVAL_29 = ~_EVAL_98;
  assign _EVAL_280 = _EVAL_55 & _EVAL_243;
  assign _EVAL_95 = ~_EVAL_185;
  assign _EVAL_101 = _EVAL_26 | _EVAL_2;
  assign _EVAL_125 = ~_EVAL_261;
  assign _EVAL_32 = ~_EVAL_96;
  assign _EVAL_21 = _EVAL_171 & _EVAL_35;
  assign _EVAL_216 = _EVAL_239 != 5'h0;
  assign _EVAL_226 = ~_EVAL_18;
  assign _EVAL_157 = _EVAL_11 <= 3'h6;
  assign _EVAL_42 = _EVAL_10[2:1];
  assign _EVAL_68 = ~_EVAL_101;
  assign _EVAL_254 = _EVAL_228 & _EVAL_232;
  assign _EVAL_149 = _EVAL_5 & _EVAL_36;
  assign _EVAL_227 = _EVAL_268 | _EVAL_2;
  assign _EVAL_153 = _EVAL_231 | _EVAL_2;
  assign _EVAL_109 = _EVAL_5 & _EVAL_141;
  assign _EVAL_55 = _EVAL_86 & _EVAL_30;
  assign _EVAL_191 = _EVAL_11 == 3'h2;
  assign _EVAL_77 = _EVAL_145 | _EVAL_2;
  assign _EVAL_53 = _EVAL_4[1];
  assign _EVAL_274 = _EVAL_3 == _EVAL_184;
  assign _EVAL_150 = _EVAL_4 == _EVAL_70;
  assign _EVAL_282 = _EVAL_53 & _EVAL_232;
  assign _EVAL_36 = _EVAL_3 == 3'h2;
  assign _EVAL_46 = _EVAL_239 != _EVAL_273;
  assign _EVAL_164 = _EVAL_224[0];
  assign _EVAL_154 = _EVAL_73[0];
  assign _EVAL_88 = ~_EVAL_93;
  assign _EVAL_135 = _EVAL_177 - 1'h1;
  assign _EVAL_159 = _EVAL_147 | _EVAL_272;
  assign _EVAL_284 = _EVAL_79[0];
  assign _EVAL_152 = 8'h1 << _EVAL_17;
  assign _EVAL_207 = _EVAL_107 | _EVAL_2;
  assign _EVAL_89 = _EVAL_15 == _EVAL_253;
  assign _EVAL_242 = _EVAL_260 & _EVAL_281;
  assign _EVAL_174 = _EVAL_17[2:1];
  assign _EVAL_194 = _EVAL_259 | _EVAL_41;
  assign _EVAL_20 = _EVAL_187 | _EVAL_2;
  assign _EVAL_25 = $signed(_EVAL_129) == 31'sh0;
  assign _EVAL_245 = ~_EVAL_34;
  assign _EVAL_189 = _EVAL_110 | _EVAL_196;
  assign _EVAL_110 = _EVAL_174 == 2'h1;
  assign _EVAL_173 = _EVAL_160 | _EVAL_2;
  assign _EVAL_56 = _EVAL_5 & _EVAL_116;
  assign _EVAL_144 = _EVAL_76 | _EVAL_186;
  assign _EVAL_40 = _EVAL_11 == 3'h1;
  assign _EVAL_240 = ~_EVAL_82;
  assign _EVAL_252 = _EVAL_13 & _EVAL_40;
  assign _EVAL_175 = _EVAL_266 ? _EVAL_152 : 8'h0;
  assign _EVAL_230 = _EVAL_71 | _EVAL_2;
  assign _EVAL_104 = ~_EVAL_148;
  assign _EVAL_74 = _EVAL_5 & _EVAL_75;
  assign _EVAL_82 = {_EVAL_50,_EVAL_144,_EVAL_195,_EVAL_170};
  assign _EVAL_58 = _EVAL_5 & _EVAL_225;
  assign _EVAL_117 = _EVAL_13 & _EVAL_102;
  assign _EVAL_219 = _EVAL_139 | _EVAL_2;
  assign _EVAL_263 = _EVAL_3 == 3'h4;
  assign _EVAL_182 = _EVAL_80 | _EVAL_2;
  assign _EVAL_146 = ~_EVAL_207;
  assign _EVAL_257 = _EVAL_166 | _EVAL_2;
  assign _EVAL_118 = ~_EVAL_162;
  assign _EVAL_217 = _EVAL_4 & _EVAL_123;
  assign _EVAL_111 = _EVAL_13 & _EVAL_283;
  assign _EVAL_60 = ~_EVAL_208;
  assign _EVAL_66 = _EVAL_194 | _EVAL_126;
  assign _EVAL_71 = _EVAL_49 == 4'h0;
  assign _EVAL_246 = _EVAL_226 | _EVAL_2;
  assign _EVAL_158 = ~_EVAL_271;
  assign _EVAL_183 = _EVAL == 3'h0;
  assign _EVAL_162 = _EVAL_151 | _EVAL_2;
  assign _EVAL_138 = _EVAL_228 & _EVAL_124;
  assign _EVAL_87 = _EVAL_11 == 3'h4;
  assign _EVAL_123 = {{28'd0}, _EVAL_269};
  assign _EVAL_255 = _EVAL_221 | _EVAL_2;
  assign _EVAL_209 = _EVAL_9 == _EVAL_270;
  assign _EVAL_129 = _EVAL_128;
  assign _EVAL_156 = _EVAL_89 | _EVAL_2;
  assign _EVAL_23 = _EVAL_5 & _EVAL_169;
  assign _EVAL_167 = _EVAL_53 & _EVAL_124;
  assign _EVAL_93 = _EVAL_157 | _EVAL_2;
  assign _EVAL_81 = ~_EVAL_230;
  assign _EVAL_281 = ~_EVAL_273;
  assign _EVAL_192 = _EVAL_11 == 3'h5;
  assign _EVAL_231 = _EVAL_57[0];
  assign _EVAL_47 = ~_EVAL_43;
  assign _EVAL_222 = _EVAL_197 - 1'h1;
  assign _EVAL_232 = ~_EVAL_124;
  assign _EVAL_96 = _EVAL_131 | _EVAL_2;
  assign _EVAL_139 = _EVAL_46 | _EVAL_103;
  assign _EVAL_113 = _EVAL_211 + 32'h1;
  assign _EVAL_276 = ~_EVAL_236;
  assign _EVAL_133 = ~_EVAL_227;
  assign _EVAL_234 = _EVAL_5 & _EVAL_37;
  assign _EVAL_140 = _EVAL_248 | _EVAL_2;
  assign _EVAL_225 = _EVAL_3 == 3'h0;
  assign _EVAL_22 = ~_EVAL_246;
  assign _EVAL_85 = _EVAL_17 == _EVAL_54;
  assign _EVAL_116 = _EVAL_3 == 3'h7;
  assign _EVAL_186 = _EVAL_164 & _EVAL_282;
  assign _EVAL_269 = ~_EVAL_108;
  assign _EVAL_127 = _EVAL_11 == 3'h0;
  assign _EVAL_266 = _EVAL_171 & _EVAL_245;
  assign _EVAL_49 = ~_EVAL_6;
  assign _EVAL_279 = _EVAL_137 | _EVAL_2;
  assign _EVAL_163 = ~_EVAL_9;
  assign _EVAL_160 = _EVAL_6 == _EVAL_82;
  assign _EVAL_151 = _EVAL <= 3'h2;
  assign _EVAL_271 = _EVAL_209 | _EVAL_2;
  assign _EVAL_250 = ~_EVAL_173;
  assign _EVAL_171 = _EVAL_0 & _EVAL_5;
  assign _EVAL_260 = _EVAL_44 | _EVAL_239;
  assign _EVAL_45 = _EVAL_150 | _EVAL_2;
  assign _EVAL_141 = _EVAL_3 == 3'h1;
  assign _EVAL_67 = ~_EVAL_180;
  assign _EVAL_168 = _EVAL_164 & _EVAL_254;
  assign _EVAL_238 = ~_EVAL_219;
  assign _EVAL_108 = _EVAL_24[1:0];
  assign _EVAL_26 = _EVAL_218 | _EVAL_65;
  assign _EVAL_236 = _EVAL_163 | _EVAL_2;
  assign _EVAL_188 = ~_EVAL_1;
  assign _EVAL_272 = _EVAL_267 & _EVAL_228;
  assign _EVAL_166 = _EVAL_163 | _EVAL_18;
  assign _EVAL_251 = _EVAL_19 | _EVAL_2;
  assign _EVAL_50 = _EVAL_76 | _EVAL_39;
  assign _EVAL_233 = _EVAL_171 | _EVAL_86;
  assign _EVAL_220 = _EVAL <= 3'h1;
  assign _EVAL_169 = _EVAL_3 == 3'h6;
  assign _EVAL_213 = _EVAL_222[0];
  assign _EVAL_69 = _EVAL <= 3'h3;
  assign _EVAL_131 = _EVAL == _EVAL_27;
  assign _EVAL_92 = _EVAL_13 & _EVAL_192;
  assign _EVAL_190 = ~_EVAL_237;
  assign _EVAL_277 = _EVAL_31[0];
  assign _EVAL_19 = _EVAL_11 == _EVAL_275;
  assign _EVAL_285 = _EVAL_280 ? _EVAL_91 : 8'h0;
  assign _EVAL_119 = _EVAL_135[0];
  assign _EVAL_30 = ~_EVAL_177;
  assign _EVAL_208 = _EVAL_155 | _EVAL_2;
  assign _EVAL_268 = _EVAL_217 == 30'h0;
  assign _EVAL_134 = ~_EVAL_284;
  assign _EVAL_243 = ~_EVAL_102;
  assign _EVAL_235 = ~_EVAL_77;
  assign _EVAL_106 = ~_EVAL_181;
  assign _EVAL_205 = ~_EVAL_100;
  assign _EVAL_72 = _EVAL_3 == 3'h5;
  assign _EVAL_124 = _EVAL_4[0];
  assign _EVAL_90 = _EVAL_147 | _EVAL_2;
  assign _EVAL_98 = _EVAL_201 | _EVAL_2;
  assign _EVAL_62 = _EVAL_13 & _EVAL_191;
  assign _EVAL_112 = ~_EVAL_198;
  assign _EVAL_181 = _EVAL_220 | _EVAL_2;
  assign _EVAL_128 = $signed(_EVAL_115) & -31'sh2000;
  assign _EVAL_51 = ~_EVAL_202;
  assign _EVAL_143 = _EVAL <= 3'h4;
  assign _EVAL_48 = _EVAL_38 | _EVAL_2;
  assign _EVAL_37 = ~_EVAL_35;
  assign _EVAL_204 = _EVAL_5 & _EVAL_263;
  assign _EVAL_239 = _EVAL_175[4:0];
  assign _EVAL_165 = ~_EVAL_279;
  assign _EVAL_283 = ~_EVAL_249;
  assign _EVAL_148 = _EVAL_274 | _EVAL_2;
  assign _EVAL_79 = _EVAL_44 >> _EVAL_17;
  assign _EVAL_94 = ~_EVAL_255;
  assign _EVAL_57 = _EVAL_264 >> _EVAL_10;
  assign _EVAL_172 = 2'h1 << _EVAL_120;
  assign _EVAL_100 = _EVAL_265 | _EVAL_2;
  assign _EVAL_91 = 8'h1 << _EVAL_10;
  assign _EVAL_86 = _EVAL_7 & _EVAL_13;
  assign _EVAL_179 = _EVAL_267 & _EVAL_53;
  assign _EVAL_259 = _EVAL_42 == 2'h1;
  assign _EVAL_126 = _EVAL_10 == 3'h4;
  assign _EVAL_121 = _EVAL_183 | _EVAL_2;
  assign _EVAL_195 = _EVAL_159 | _EVAL_78;
  assign _EVAL_198 = _EVAL_134 | _EVAL_2;
  assign _EVAL_24 = 5'h3 << _EVAL_15;
  assign _EVAL_248 = _EVAL_16 == _EVAL_193;
  assign _EVAL_80 = _EVAL != 3'h0;
  assign _EVAL_78 = _EVAL_164 & _EVAL_138;
  assign _EVAL_249 = ~_EVAL_197;
  assign _EVAL_97 = ~_EVAL_48;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_27 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_34 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_44 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_54 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_70 = _RAND_4[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_99 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_161 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_177 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_184 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_193 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_197 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_200 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_211 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_229 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_253 = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_270 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_275 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_14) begin
    if (_EVAL_21) begin
      _EVAL_27 <= _EVAL;
    end
    if (_EVAL_2) begin
      _EVAL_34 <= 1'h0;
    end else if (_EVAL_171) begin
      if (_EVAL_245) begin
        _EVAL_34 <= 1'h0;
      end else begin
        _EVAL_34 <= _EVAL_277;
      end
    end
    if (_EVAL_2) begin
      _EVAL_44 <= 5'h0;
    end else begin
      _EVAL_44 <= _EVAL_242;
    end
    if (_EVAL_21) begin
      _EVAL_54 <= _EVAL_17;
    end
    if (_EVAL_21) begin
      _EVAL_70 <= _EVAL_4;
    end
    if (_EVAL_176) begin
      _EVAL_99 <= _EVAL_12;
    end
    if (_EVAL_2) begin
      _EVAL_161 <= 1'h0;
    end else if (_EVAL_171) begin
      if (_EVAL_35) begin
        _EVAL_161 <= 1'h0;
      end else begin
        _EVAL_161 <= _EVAL_154;
      end
    end
    if (_EVAL_2) begin
      _EVAL_177 <= 1'h0;
    end else if (_EVAL_86) begin
      if (_EVAL_30) begin
        _EVAL_177 <= 1'h0;
      end else begin
        _EVAL_177 <= _EVAL_119;
      end
    end
    if (_EVAL_21) begin
      _EVAL_184 <= _EVAL_3;
    end
    if (_EVAL_176) begin
      _EVAL_193 <= _EVAL_16;
    end
    if (_EVAL_2) begin
      _EVAL_197 <= 1'h0;
    end else if (_EVAL_86) begin
      if (_EVAL_249) begin
        _EVAL_197 <= 1'h0;
      end else begin
        _EVAL_197 <= _EVAL_213;
      end
    end
    if (_EVAL_176) begin
      _EVAL_200 <= _EVAL_10;
    end
    if (_EVAL_2) begin
      _EVAL_211 <= 32'h0;
    end else if (_EVAL_233) begin
      _EVAL_211 <= 32'h0;
    end else begin
      _EVAL_211 <= _EVAL_262;
    end
    if (_EVAL_176) begin
      _EVAL_229 <= _EVAL_8;
    end
    if (_EVAL_21) begin
      _EVAL_253 <= _EVAL_15;
    end
    if (_EVAL_176) begin
      _EVAL_270 <= _EVAL_9;
    end
    if (_EVAL_176) begin
      _EVAL_275 <= _EVAL_11;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1596d71e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56fb871d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d11108a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9f23fbc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(377bdbda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9ae872c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8260212a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9921198)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bc196e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e1d648a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3769b33d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e18389ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ab63fca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d34aaab9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f4bb00b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e9e6fc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce15ec2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0ce27d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(820af394)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79808ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29289122)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b892417e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3183cec0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa571a8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d15d71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86546731)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8a380b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6aac8835)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(697593cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8818e591)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(947e8384)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f00616ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b848bd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b883bdff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9bfbef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f0e8c3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f731a641)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2658ee53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(feace9d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5504eb2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e05b7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(956592c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48f86f2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80625db7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bef25851)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fae2013)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cd7d0c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45ffb970)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5368afcb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa6623e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5ca522c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0159ecf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d3e8929)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91277150)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6197d9e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a5d4de1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d83b4d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(689f50d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f787914c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e386f58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e8ae8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13822e39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7c27495)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8daed546)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccdf4eee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(679676c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17e3ee7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56fd5752)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e0adf3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3057aa6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed114575)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(600bd221)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(456a8953)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49a5db30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc30db05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19a5616c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d0b319a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(643a8060)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fcf5c44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d2fcae8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bb5bb12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f8ad5eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bffdaca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6eed72f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2797d7a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7bf5969)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b45e7ecd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cf3a629)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(881615a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdbc5cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70690027)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12f120)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a5170f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
