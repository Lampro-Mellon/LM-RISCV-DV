//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_176_assert(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [14:0] _EVAL_3,
  input  [3:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [1:0]  _EVAL_7,
  input  [2:0]  _EVAL_8,
  input  [1:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13
);
  wire  _EVAL_14;
  wire  _EVAL_15;
  reg  _EVAL_16;
  reg [31:0] _RAND_0;
  wire [4:0] _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  reg [2:0] _EVAL_22;
  reg [31:0] _RAND_1;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire [7:0] _EVAL_25;
  wire [1:0] _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  reg [2:0] _EVAL_29;
  reg [31:0] _RAND_2;
  wire [7:0] _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  reg  _EVAL_36;
  reg [31:0] _RAND_3;
  wire  _EVAL_37;
  wire [4:0] _EVAL_38;
  reg [2:0] _EVAL_39;
  reg [31:0] _RAND_4;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire [4:0] _EVAL_42;
  wire  _EVAL_43;
  wire [1:0] _EVAL_44;
  wire  _EVAL_45;
  reg  _EVAL_46;
  reg [31:0] _RAND_5;
  wire  _EVAL_47;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire [4:0] _EVAL_58;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire [15:0] _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire [32:0] _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  reg [2:0] _EVAL_73;
  reg [31:0] _RAND_6;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  reg [4:0] _EVAL_84;
  reg [31:0] _RAND_7;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire [14:0] _EVAL_91;
  wire [1:0] _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire [14:0] _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  reg [1:0] _EVAL_107;
  reg [31:0] _RAND_8;
  wire  _EVAL_108;
  wire [1:0] _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire [3:0] _EVAL_117;
  wire  _EVAL_118;
  wire [4:0] _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire [7:0] _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  reg [14:0] _EVAL_127;
  reg [31:0] _RAND_9;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  reg [2:0] _EVAL_138;
  reg [31:0] _RAND_10;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire [4:0] _EVAL_142;
  reg [31:0] _EVAL_143;
  reg [31:0] _RAND_11;
  wire  _EVAL_144;
  wire [14:0] _EVAL_145;
  wire  _EVAL_146;
  reg  _EVAL_147;
  reg [31:0] _RAND_12;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire [7:0] _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire [3:0] _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire [1:0] _EVAL_169;
  wire [4:0] _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire [15:0] _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire [15:0] _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire [3:0] _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire [31:0] _EVAL_184;
  wire [4:0] _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire [1:0] _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire [1:0] _EVAL_194;
  reg [1:0] _EVAL_195;
  reg [31:0] _RAND_13;
  wire  _EVAL_196;
  wire [1:0] _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire [3:0] _EVAL_203;
  wire  _EVAL_204;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_106 = ~_EVAL_188;
  assign _EVAL_193 = _EVAL_1 <= 3'h4;
  assign _EVAL_128 = _EVAL_162 & _EVAL_187;
  assign _EVAL_149 = ~_EVAL_24;
  assign _EVAL_100 = {{13'd0}, _EVAL_197};
  assign _EVAL_54 = _EVAL_0 & _EVAL_37;
  assign _EVAL_53 = ~_EVAL_49;
  assign _EVAL_64 = _EVAL_60 | _EVAL_140;
  assign _EVAL_38 = _EVAL_84 >> _EVAL_2;
  assign _EVAL_141 = _EVAL_6 & _EVAL_11;
  assign _EVAL_181 = _EVAL_12 == _EVAL_22;
  assign _EVAL_88 = ~_EVAL_131;
  assign _EVAL_159 = _EVAL_4 & _EVAL_179;
  assign _EVAL_157 = _EVAL_162 & _EVAL_111;
  assign _EVAL_162 = _EVAL_194[1];
  assign _EVAL_115 = _EVAL_8 == 3'h4;
  assign _EVAL_45 = ~_EVAL_166;
  assign _EVAL_31 = ~_EVAL_37;
  assign _EVAL_131 = _EVAL_1 <= 3'h1;
  assign _EVAL_179 = ~_EVAL_203;
  assign _EVAL_65 = _EVAL_11 & _EVAL_43;
  assign _EVAL_49 = ~_EVAL_147;
  assign _EVAL_191 = _EVAL_111 & _EVAL_14;
  assign _EVAL_167 = _EVAL_11 & _EVAL_20;
  assign _EVAL_71 = _EVAL_180 | _EVAL_112;
  assign _EVAL_94 = _EVAL_58 != _EVAL_119;
  assign _EVAL_180 = _EVAL_164 | _EVAL_157;
  assign _EVAL_135 = _EVAL_1 <= 3'h3;
  assign _EVAL_189 = _EVAL_7 >= 2'h2;
  assign _EVAL_87 = _EVAL_7 == _EVAL_195;
  assign _EVAL_81 = _EVAL_143 < plusarg_reader_out;
  assign _EVAL_153 = _EVAL_141 & _EVAL_113;
  assign _EVAL_185 = _EVAL_42 >> _EVAL;
  assign _EVAL_102 = ~_EVAL_87;
  assign _EVAL_145 = _EVAL_3 ^ 15'h4000;
  assign _EVAL_69 = _EVAL_141 | _EVAL_75;
  assign _EVAL_161 = _EVAL_2 == _EVAL_138;
  assign _EVAL_125 = _EVAL_75 & _EVAL_49;
  assign _EVAL_101 = _EVAL_11 & _EVAL_52;
  assign _EVAL_76 = ~_EVAL_57;
  assign _EVAL_196 = _EVAL_180 | _EVAL_183;
  assign _EVAL_175 = _EVAL_89 & _EVAL_163;
  assign _EVAL_190 = _EVAL_36 - 1'h1;
  assign _EVAL_112 = _EVAL_136 & _EVAL_133;
  assign _EVAL_118 = _EVAL_9[0];
  assign _EVAL_79 = _EVAL_64 | _EVAL_81;
  assign _EVAL_34 = ~_EVAL_193;
  assign _EVAL_122 = _EVAL_185[0];
  assign _EVAL_170 = 5'h3 << _EVAL_9;
  assign _EVAL_97 = ~_EVAL_175;
  assign _EVAL_61 = ~_EVAL_13;
  assign _EVAL_105 = _EVAL_12 == 3'h7;
  assign _EVAL_44 = _EVAL_46 - 1'h1;
  assign _EVAL_150 = ~_EVAL_149;
  assign _EVAL_155 = _EVAL_0 & _EVAL_27;
  assign _EVAL_37 = _EVAL_8 == 3'h6;
  assign _EVAL_151 = _EVAL_136 & _EVAL_77;
  assign _EVAL_95 = _EVAL_75 & _EVAL_55;
  assign _EVAL_99 = _EVAL_0 & _EVAL_115;
  assign _EVAL_130 = _EVAL_58 != 5'h0;
  assign _EVAL_186 = _EVAL_95 & _EVAL_31;
  assign _EVAL_28 = _EVAL_8 == _EVAL_39;
  assign _EVAL_25 = 8'h1 << _EVAL_2;
  assign _EVAL_20 = _EVAL_12 == 3'h1;
  assign _EVAL_117 = ~_EVAL_4;
  assign _EVAL_176 = $signed(_EVAL_173) & -16'sh1000;
  assign _EVAL_113 = ~_EVAL_16;
  assign _EVAL_123 = _EVAL_8 == 3'h2;
  assign _EVAL_82 = _EVAL_26[0];
  assign _EVAL_55 = ~_EVAL_36;
  assign _EVAL_146 = _EVAL_12 == 3'h2;
  assign _EVAL_188 = _EVAL_4 == _EVAL_203;
  assign _EVAL_120 = ~_EVAL_199;
  assign _EVAL_18 = _EVAL_12 == 3'h0;
  assign _EVAL_136 = _EVAL_194[0];
  assign _EVAL_111 = _EVAL_3[1];
  assign _EVAL_32 = _EVAL_178 | _EVAL_72;
  assign _EVAL_66 = _EVAL_44[0];
  assign _EVAL_56 = ~_EVAL_161;
  assign _EVAL_156 = _EVAL_94 | _EVAL_40;
  assign _EVAL_21 = _EVAL_190[0];
  assign _EVAL_42 = _EVAL_58 | _EVAL_84;
  assign _EVAL_201 = _EVAL_178 | _EVAL_151;
  assign _EVAL_198 = _EVAL_141 & _EVAL_108;
  assign _EVAL_62 = _EVAL_109[0];
  assign _EVAL_121 = ~_EVAL_122;
  assign _EVAL_103 = ~_EVAL_156;
  assign _EVAL_158 = _EVAL_187 & _EVAL_14;
  assign _EVAL_67 = _EVAL_2 <= 3'h4;
  assign _EVAL_197 = ~_EVAL_169;
  assign _EVAL_90 = ~_EVAL_68;
  assign _EVAL_19 = _EVAL_84 != 5'h0;
  assign _EVAL_93 = _EVAL_8 == 3'h0;
  assign _EVAL_139 = ~_EVAL_164;
  assign _EVAL_114 = _EVAL_11 & _EVAL_146;
  assign _EVAL_152 = _EVAL_198 ? _EVAL_25 : 8'h0;
  assign _EVAL_178 = _EVAL_164 | _EVAL_128;
  assign _EVAL_58 = _EVAL_152[4:0];
  assign _EVAL_86 = ~_EVAL_113;
  assign _EVAL_43 = _EVAL_12 == 3'h5;
  assign _EVAL_140 = plusarg_reader_out == 32'h0;
  assign _EVAL_52 = _EVAL_12 == 3'h6;
  assign _EVAL_177 = ~_EVAL_189;
  assign _EVAL_192 = ~_EVAL_28;
  assign _EVAL_169 = _EVAL_170[1:0];
  assign _EVAL_68 = _EVAL_1 == _EVAL_29;
  assign _EVAL_174 = ~_EVAL_137;
  assign _EVAL_116 = _EVAL_11 & _EVAL_15;
  assign _EVAL_40 = ~_EVAL_130;
  assign _EVAL_80 = _EVAL_9 == _EVAL_107;
  assign _EVAL_204 = _EVAL_159 == 4'h0;
  assign _EVAL_35 = _EVAL_3[0];
  assign _EVAL_51 = _EVAL_8 == 3'h5;
  assign _EVAL_194 = _EVAL_92 | 2'h1;
  assign _EVAL_129 = _EVAL_11 & _EVAL_18;
  assign _EVAL_166 = _EVAL_91 == 15'h0;
  assign _EVAL_33 = _EVAL_1 <= 3'h2;
  assign _EVAL_60 = ~_EVAL_19;
  assign _EVAL_142 = ~_EVAL_119;
  assign _EVAL_110 = ~_EVAL_33;
  assign _EVAL_91 = _EVAL_3 & _EVAL_100;
  assign _EVAL_199 = _EVAL == _EVAL_73;
  assign _EVAL_63 = _EVAL_176;
  assign _EVAL_89 = _EVAL_9 <= 2'h2;
  assign _EVAL_144 = ~_EVAL_135;
  assign _EVAL_85 = ~_EVAL_67;
  assign _EVAL_108 = ~_EVAL_46;
  assign _EVAL_98 = ~_EVAL_79;
  assign _EVAL_14 = ~_EVAL_35;
  assign _EVAL_83 = _EVAL_11 & _EVAL_168;
  assign _EVAL_124 = _EVAL_186 ? _EVAL_30 : 8'h0;
  assign _EVAL_72 = _EVAL_136 & _EVAL_158;
  assign _EVAL_173 = {1'b0,$signed(_EVAL_145)};
  assign _EVAL_119 = _EVAL_124[4:0];
  assign _EVAL_126 = _EVAL_0 & _EVAL_53;
  assign _EVAL_184 = _EVAL_70[31:0];
  assign _EVAL_17 = _EVAL_84 | _EVAL_58;
  assign _EVAL_109 = _EVAL_16 - 1'h1;
  assign _EVAL_154 = ~_EVAL_80;
  assign _EVAL_160 = _EVAL_11 & _EVAL_86;
  assign _EVAL_92 = 2'h1 << _EVAL_118;
  assign _EVAL_26 = _EVAL_147 - 1'h1;
  assign _EVAL_137 = _EVAL_1 != 3'h0;
  assign _EVAL_163 = $signed(_EVAL_63) == 16'sh0;
  assign _EVAL_27 = _EVAL_8 == 3'h1;
  assign _EVAL_182 = _EVAL <= 3'h4;
  assign _EVAL_30 = 8'h1 << _EVAL;
  assign _EVAL_133 = _EVAL_111 & _EVAL_35;
  assign _EVAL_78 = ~_EVAL_182;
  assign _EVAL_57 = _EVAL_8 <= 3'h6;
  assign _EVAL_183 = _EVAL_136 & _EVAL_191;
  assign _EVAL_74 = _EVAL_0 & _EVAL_51;
  assign _EVAL_50 = _EVAL_117 == 4'h0;
  assign _EVAL_134 = _EVAL_0 & _EVAL_93;
  assign _EVAL_165 = ~_EVAL_50;
  assign _EVAL_47 = ~_EVAL_172;
  assign _EVAL_15 = _EVAL_12 == 3'h3;
  assign _EVAL_202 = _EVAL_1 == 3'h0;
  assign _EVAL_171 = _EVAL_11 & _EVAL_105;
  assign _EVAL_75 = _EVAL_10 & _EVAL_0;
  assign _EVAL_70 = _EVAL_143 + 32'h1;
  assign _EVAL_104 = _EVAL_0 & _EVAL_123;
  assign _EVAL_77 = _EVAL_187 & _EVAL_35;
  assign _EVAL_24 = _EVAL_38[0];
  assign _EVAL_23 = ~_EVAL_181;
  assign _EVAL_164 = _EVAL_9 >= 2'h2;
  assign _EVAL_200 = ~_EVAL_202;
  assign _EVAL_41 = ~_EVAL_204;
  assign _EVAL_203 = {_EVAL_71,_EVAL_196,_EVAL_201,_EVAL_32};
  assign _EVAL_172 = _EVAL_3 == _EVAL_127;
  assign _EVAL_168 = _EVAL_12 == 3'h4;
  assign _EVAL_187 = ~_EVAL_111;
  assign _EVAL_96 = ~_EVAL_61;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_16 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_22 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_29 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_36 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_39 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_46 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_73 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_84 = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_107 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_127 = _RAND_9[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_138 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_143 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_147 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_195 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_5) begin
    if (_EVAL_141) begin
      if (_EVAL_113) begin
        _EVAL_16 <= 1'h0;
      end else begin
        _EVAL_16 <= _EVAL_62;
      end
    end
    if (_EVAL_153) begin
      _EVAL_22 <= _EVAL_12;
    end
    if (_EVAL_153) begin
      _EVAL_29 <= _EVAL_1;
    end
    if (_EVAL_75) begin
      if (_EVAL_55) begin
        _EVAL_36 <= 1'h0;
      end else begin
        _EVAL_36 <= _EVAL_21;
      end
    end
    if (_EVAL_125) begin
      _EVAL_39 <= _EVAL_8;
    end
    if (_EVAL_141) begin
      if (_EVAL_108) begin
        _EVAL_46 <= 1'h0;
      end else begin
        _EVAL_46 <= _EVAL_66;
      end
    end
    if (_EVAL_125) begin
      _EVAL_73 <= _EVAL;
    end
    _EVAL_84 <= _EVAL_17 & _EVAL_142;
    if (_EVAL_153) begin
      _EVAL_107 <= _EVAL_9;
    end
    if (_EVAL_153) begin
      _EVAL_127 <= _EVAL_3;
    end
    if (_EVAL_153) begin
      _EVAL_138 <= _EVAL_2;
    end
    if (_EVAL_69) begin
      _EVAL_143 <= 32'h0;
    end else begin
      _EVAL_143 <= _EVAL_184;
    end
    if (_EVAL_75) begin
      if (_EVAL_49) begin
        _EVAL_147 <= 1'h0;
      end else begin
        _EVAL_147 <= _EVAL_82;
      end
    end
    if (_EVAL_125) begin
      _EVAL_195 <= _EVAL_7;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(288f7fe0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26ba438d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(209fe8e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78e6c073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1df7baef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df275cb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f723c44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4d3bbf0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abbdbe1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50b3dba2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(616a730b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fa40640)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(588ee2fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1be3f668)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(531165f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b3e5b7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b04a078a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_15) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(151db744)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27ffe693)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7e138bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a88941c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(832a2f23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2f1b03f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_15) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e98919b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25cd420f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7f38a3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d75f6d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea510d66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef72ccf1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78aaf8e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa4ecc49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef800dd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb37614c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e66a53d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(781a99a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae542bd9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f153b933)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8a85551)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(809a9c60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c661c3ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28121978)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d4d2e22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d97fde5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1a4c508)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f00fc8dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bd11c33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc494ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a735556)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(928493d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84d0092a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9f56510)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48b8e9df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(161a701e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fded497)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62eed0c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b50cd0a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2604eba2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6a7b77a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8597974)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9432dfc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e797217)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24bbc2e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92cef5d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e54899f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9113b407)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61ff4225)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea9e0e51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(503bd64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d70a4bf0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d296070e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dcbc300)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31c50a9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a307cb1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
