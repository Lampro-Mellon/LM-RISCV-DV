//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_100_assert(
  input         _EVAL,
  input  [1:0]  _EVAL_0,
  input         _EVAL_1,
  input  [3:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  input  [14:0] _EVAL_12,
  input         _EVAL_13,
  input  [1:0]  _EVAL_14
);
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire [3:0] _EVAL_22;
  wire [4:0] _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire [1:0] _EVAL_29;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  reg  _EVAL_35;
  reg [31:0] _RAND_0;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  reg [1:0] _EVAL_40;
  reg [31:0] _RAND_1;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire [14:0] _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire [14:0] _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire [4:0] _EVAL_60;
  wire  _EVAL_61;
  wire [7:0] _EVAL_62;
  wire [1:0] _EVAL_63;
  wire  _EVAL_64;
  reg [31:0] _EVAL_65;
  reg [31:0] _RAND_2;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire [1:0] _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire [1:0] _EVAL_74;
  wire  _EVAL_75;
  wire [14:0] _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  reg [1:0] _EVAL_79;
  reg [31:0] _RAND_3;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire [7:0] _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire [15:0] _EVAL_86;
  wire  _EVAL_87;
  wire [4:0] _EVAL_88;
  wire [4:0] _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire [4:0] _EVAL_94;
  wire  _EVAL_95;
  reg [2:0] _EVAL_96;
  reg [31:0] _RAND_4;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire [15:0] _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  reg  _EVAL_107;
  reg [31:0] _RAND_5;
  wire  _EVAL_109;
  wire [1:0] _EVAL_110;
  wire  _EVAL_111;
  wire [3:0] _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire [7:0] _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  reg [14:0] _EVAL_125;
  reg [31:0] _RAND_6;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire [4:0] _EVAL_129;
  wire  _EVAL_131;
  wire [1:0] _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_136;
  wire [1:0] _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire [7:0] _EVAL_140;
  reg [2:0] _EVAL_142;
  reg [31:0] _RAND_7;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire [4:0] _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire [1:0] _EVAL_152;
  wire [3:0] _EVAL_153;
  wire [31:0] _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  reg  _EVAL_160;
  reg [31:0] _RAND_8;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire [4:0] _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire [15:0] _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [1:0] _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  reg  _EVAL_180;
  reg [31:0] _RAND_9;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire [4:0] _EVAL_191;
  reg [2:0] _EVAL_192;
  reg [31:0] _RAND_10;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  reg [4:0] _EVAL_198;
  reg [31:0] _RAND_11;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  reg [2:0] _EVAL_206;
  reg [31:0] _RAND_12;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire [3:0] _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire [1:0] _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire [32:0] _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  reg [2:0] _EVAL_249;
  reg [31:0] _RAND_13;
  wire  _EVAL_250;
  wire  _EVAL_251;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_48 = _EVAL_106 | _EVAL_1;
  assign _EVAL_15 = ~_EVAL_193;
  assign _EVAL_44 = _EVAL_3 == _EVAL_249;
  assign _EVAL_196 = _EVAL_90 & _EVAL_85;
  assign _EVAL_185 = _EVAL_65 < plusarg_reader_out;
  assign _EVAL_161 = _EVAL_225 | _EVAL_1;
  assign _EVAL_175 = _EVAL_231 | _EVAL_181;
  assign _EVAL_123 = _EVAL_7 == 3'h4;
  assign _EVAL_131 = _EVAL_101 & _EVAL_150;
  assign _EVAL_57 = _EVAL_174 == 2'h0;
  assign _EVAL_208 = _EVAL_173 | _EVAL_1;
  assign _EVAL_218 = _EVAL_13 & _EVAL_121;
  assign _EVAL_138 = ~_EVAL_150;
  assign _EVAL_216 = _EVAL_191 != _EVAL_60;
  assign _EVAL_238 = ~_EVAL_28;
  assign _EVAL_190 = _EVAL_13 & _EVAL_26;
  assign _EVAL_201 = ~_EVAL_146;
  assign _EVAL_151 = _EVAL_6 <= 3'h1;
  assign _EVAL_227 = _EVAL_163[0];
  assign _EVAL_225 = _EVAL_158 & _EVAL_156;
  assign _EVAL_231 = _EVAL_14 >= 2'h2;
  assign _EVAL_85 = _EVAL_12[1];
  assign _EVAL_122 = 8'h1 << _EVAL_11;
  assign _EVAL_222 = _EVAL_2 & _EVAL_112;
  assign _EVAL_116 = ~_EVAL_115;
  assign _EVAL_46 = _EVAL_220 | _EVAL_1;
  assign _EVAL_211 = _EVAL_50 | _EVAL_186;
  assign _EVAL_100 = _EVAL_246 | _EVAL_95;
  assign _EVAL_195 = ~_EVAL_77;
  assign _EVAL_152 = _EVAL_180 - 1'h1;
  assign _EVAL_226 = _EVAL_101 & _EVAL_138;
  assign _EVAL_128 = _EVAL_118 | _EVAL_1;
  assign _EVAL_83 = 8'h1 << _EVAL_5;
  assign _EVAL_129 = ~_EVAL_60;
  assign _EVAL_17 = _EVAL_175 | _EVAL_205;
  assign _EVAL_159 = ~_EVAL_194;
  assign _EVAL_69 = _EVAL_3 == 3'h1;
  assign _EVAL_248 = _EVAL_3 == 3'h2;
  assign _EVAL_165 = _EVAL_68[0];
  assign _EVAL_93 = ~_EVAL_52;
  assign _EVAL_214 = _EVAL_95 & _EVAL_73;
  assign _EVAL_59 = _EVAL_13 & _EVAL_114;
  assign _EVAL_233 = _EVAL_198 != 5'h0;
  assign _EVAL_97 = ~_EVAL_18;
  assign _EVAL_219 = ~_EVAL_236;
  assign _EVAL_207 = _EVAL_182 | _EVAL_57;
  assign _EVAL_243 = _EVAL_61 & _EVAL_145;
  assign _EVAL_49 = ~_EVAL_1;
  assign _EVAL_140 = _EVAL_133 ? _EVAL_83 : 8'h0;
  assign _EVAL_189 = ~_EVAL_208;
  assign _EVAL_209 = ~_EVAL_105;
  assign _EVAL_164 = ~_EVAL_37;
  assign _EVAL_204 = ~_EVAL_197;
  assign _EVAL_110 = _EVAL_11[2:1];
  assign _EVAL_244 = ~_EVAL_136;
  assign _EVAL_18 = _EVAL_23[0];
  assign _EVAL_153 = ~_EVAL_2;
  assign _EVAL_186 = plusarg_reader_out == 32'h0;
  assign _EVAL_39 = _EVAL_95 & _EVAL_247;
  assign _EVAL_156 = $signed(_EVAL_99) == 16'sh0;
  assign _EVAL_61 = _EVAL_137[0];
  assign _EVAL_38 = _EVAL_111 | _EVAL_1;
  assign _EVAL_167 = _EVAL_3 == 3'h5;
  assign _EVAL_197 = _EVAL_70 | _EVAL_1;
  assign _EVAL_42 = ~_EVAL_178;
  assign _EVAL_84 = ~_EVAL_247;
  assign _EVAL_126 = _EVAL_203 | _EVAL_1;
  assign _EVAL_136 = _EVAL_213 | _EVAL_1;
  assign _EVAL_75 = _EVAL_13 & _EVAL_80;
  assign _EVAL_134 = _EVAL_237 | _EVAL_1;
  assign _EVAL_26 = _EVAL_7 == 3'h5;
  assign _EVAL_246 = _EVAL_10 & _EVAL_9;
  assign _EVAL_31 = ~_EVAL_33;
  assign _EVAL_21 = _EVAL_239 | _EVAL_81;
  assign _EVAL_202 = _EVAL_211 | _EVAL_185;
  assign _EVAL_149 = _EVAL_191 | _EVAL_198;
  assign _EVAL_16 = _EVAL_3 == 3'h0;
  assign _EVAL_113 = _EVAL_29[0];
  assign _EVAL_117 = _EVAL_85 & _EVAL_138;
  assign _EVAL_239 = _EVAL_231 | _EVAL_196;
  assign _EVAL_34 = ~_EVAL_80;
  assign _EVAL_102 = _EVAL_162 | _EVAL_242;
  assign _EVAL_23 = _EVAL_198 >> _EVAL_5;
  assign _EVAL_166 = _EVAL_3 == 3'h7;
  assign _EVAL_106 = _EVAL_5 == _EVAL_206;
  assign _EVAL_162 = _EVAL_187 | _EVAL_124;
  assign _EVAL_28 = _EVAL_212 | _EVAL_1;
  assign _EVAL_99 = _EVAL_171;
  assign _EVAL_154 = _EVAL_245[31:0];
  assign _EVAL_111 = _EVAL_6 <= 3'h4;
  assign _EVAL_251 = _EVAL_5 == 3'h4;
  assign _EVAL_169 = _EVAL_152[0];
  assign _EVAL_163 = _EVAL_149 >> _EVAL_11;
  assign _EVAL_95 = _EVAL_8 & _EVAL_13;
  assign _EVAL_235 = ~_EVAL_103;
  assign _EVAL_76 = {{13'd0}, _EVAL_63};
  assign _EVAL_78 = ~_EVAL_134;
  assign _EVAL_87 = _EVAL_214 & _EVAL_34;
  assign _EVAL_232 = _EVAL_94[1:0];
  assign _EVAL_212 = _EVAL_2 == _EVAL_22;
  assign _EVAL_92 = ~_EVAL_35;
  assign _EVAL_114 = _EVAL_7 == 3'h1;
  assign _EVAL_217 = ~_EVAL_221;
  assign _EVAL_70 = _EVAL_216 | _EVAL_217;
  assign _EVAL_170 = _EVAL_9 & _EVAL_179;
  assign _EVAL_230 = ~_EVAL_128;
  assign _EVAL_224 = _EVAL_246 & _EVAL_92;
  assign _EVAL_228 = ~_EVAL_46;
  assign _EVAL_146 = _EVAL_202 | _EVAL_1;
  assign _EVAL_24 = _EVAL_9 & _EVAL_166;
  assign _EVAL_20 = _EVAL_9 & _EVAL_248;
  assign _EVAL_155 = _EVAL_12 == _EVAL_125;
  assign _EVAL_41 = ~_EVAL_48;
  assign _EVAL_80 = _EVAL_7 == 3'h6;
  assign _EVAL_179 = ~_EVAL_92;
  assign _EVAL_74 = 2'h1 << _EVAL_54;
  assign _EVAL_171 = $signed(_EVAL_86) & -16'sh1000;
  assign _EVAL_104 = ~_EVAL_51;
  assign _EVAL_77 = _EVAL_102 | _EVAL_1;
  assign _EVAL_72 = _EVAL_222 == 4'h0;
  assign _EVAL_199 = _EVAL_7 == 3'h2;
  assign _EVAL_29 = _EVAL_107 - 1'h1;
  assign _EVAL_52 = _EVAL_155 | _EVAL_1;
  assign _EVAL_229 = _EVAL_9 & _EVAL_167;
  assign _EVAL_89 = _EVAL_88 & _EVAL_129;
  assign _EVAL_205 = _EVAL_61 & _EVAL_131;
  assign _EVAL_86 = {1'b0,$signed(_EVAL_45)};
  assign _EVAL_127 = _EVAL_239 | _EVAL_243;
  assign _EVAL_68 = _EVAL_35 - 1'h1;
  assign _EVAL_32 = _EVAL_6 <= 3'h3;
  assign _EVAL_64 = _EVAL_6 == 3'h0;
  assign _EVAL_56 = _EVAL_72 | _EVAL_1;
  assign _EVAL_50 = ~_EVAL_233;
  assign _EVAL_150 = _EVAL_12[0];
  assign _EVAL_90 = _EVAL_137[1];
  assign _EVAL_135 = _EVAL_13 & _EVAL_123;
  assign _EVAL_245 = _EVAL_65 + 32'h1;
  assign _EVAL_67 = ~_EVAL_25;
  assign _EVAL_145 = _EVAL_85 & _EVAL_150;
  assign _EVAL_81 = _EVAL_61 & _EVAL_117;
  assign _EVAL_91 = _EVAL_168 | _EVAL_1;
  assign _EVAL_144 = _EVAL_153 == 4'h0;
  assign _EVAL_237 = _EVAL_7 == _EVAL_192;
  assign _EVAL_36 = _EVAL_97 | _EVAL_1;
  assign _EVAL_183 = _EVAL_9 & _EVAL_177;
  assign _EVAL_236 = _EVAL_172 | _EVAL_1;
  assign _EVAL_168 = _EVAL_0 >= 2'h2;
  assign _EVAL_181 = _EVAL_90 & _EVAL_101;
  assign _EVAL_241 = _EVAL_7 <= 3'h6;
  assign _EVAL_82 = _EVAL_13 & _EVAL_199;
  assign _EVAL_174 = _EVAL_5[2:1];
  assign _EVAL_173 = _EVAL_53 == 15'h0;
  assign _EVAL_242 = _EVAL_11 == 3'h4;
  assign _EVAL_221 = _EVAL_191 != 5'h0;
  assign _EVAL_177 = _EVAL_3 == 3'h6;
  assign _EVAL_66 = _EVAL_13 & _EVAL_84;
  assign _EVAL_54 = _EVAL_14[0];
  assign _EVAL_53 = _EVAL_12 & _EVAL_76;
  assign _EVAL_132 = _EVAL_160 - 1'h1;
  assign _EVAL_43 = _EVAL_132[0];
  assign _EVAL_62 = _EVAL_87 ? _EVAL_122 : 8'h0;
  assign _EVAL_98 = ~_EVAL_36;
  assign _EVAL_158 = _EVAL_14 <= 2'h2;
  assign _EVAL_47 = ~_EVAL_223;
  assign _EVAL_203 = _EVAL_0 == _EVAL_79;
  assign _EVAL_200 = _EVAL_61 & _EVAL_226;
  assign _EVAL_25 = _EVAL_44 | _EVAL_1;
  assign _EVAL_240 = ~_EVAL_56;
  assign _EVAL_101 = ~_EVAL_85;
  assign _EVAL_58 = _EVAL_9 & _EVAL_19;
  assign _EVAL_73 = ~_EVAL_107;
  assign _EVAL_182 = _EVAL_174 == 2'h1;
  assign _EVAL_220 = _EVAL_207 | _EVAL_251;
  assign _EVAL_137 = _EVAL_74 | 2'h1;
  assign _EVAL_139 = _EVAL_9 & _EVAL_69;
  assign _EVAL_118 = _EVAL_6 != 3'h0;
  assign _EVAL_105 = _EVAL_148 | _EVAL_1;
  assign _EVAL_124 = _EVAL_110 == 2'h0;
  assign _EVAL_27 = _EVAL_9 & _EVAL_109;
  assign _EVAL_37 = _EVAL_144 | _EVAL_1;
  assign _EVAL_119 = _EVAL_175 | _EVAL_200;
  assign _EVAL_143 = ~_EVAL_91;
  assign _EVAL_247 = ~_EVAL_180;
  assign _EVAL_109 = _EVAL_3 == 3'h3;
  assign _EVAL_193 = _EVAL_234 | _EVAL_1;
  assign _EVAL_184 = ~_EVAL_161;
  assign _EVAL_33 = _EVAL_64 | _EVAL_1;
  assign _EVAL_223 = _EVAL_227 | _EVAL_1;
  assign _EVAL_213 = _EVAL_14 == _EVAL_40;
  assign _EVAL_133 = _EVAL_246 & _EVAL_120;
  assign _EVAL_22 = {_EVAL_127,_EVAL_21,_EVAL_17,_EVAL_119};
  assign _EVAL_103 = _EVAL_241 | _EVAL_1;
  assign _EVAL_60 = _EVAL_62[4:0];
  assign _EVAL_112 = ~_EVAL_22;
  assign _EVAL_121 = _EVAL_7 == 3'h0;
  assign _EVAL_234 = _EVAL_6 == _EVAL_96;
  assign _EVAL_191 = _EVAL_140[4:0];
  assign _EVAL_88 = _EVAL_198 | _EVAL_191;
  assign _EVAL_194 = _EVAL_231 | _EVAL_1;
  assign _EVAL_45 = _EVAL_12 ^ 15'h4000;
  assign _EVAL_172 = ~_EVAL;
  assign _EVAL_147 = ~_EVAL_38;
  assign _EVAL_51 = _EVAL_151 | _EVAL_1;
  assign _EVAL_120 = ~_EVAL_160;
  assign _EVAL_178 = _EVAL_215 | _EVAL_1;
  assign _EVAL_187 = _EVAL_110 == 2'h1;
  assign _EVAL_94 = 5'h3 << _EVAL_14;
  assign _EVAL_63 = ~_EVAL_232;
  assign _EVAL_148 = _EVAL_11 == _EVAL_142;
  assign _EVAL_19 = _EVAL_3 == 3'h4;
  assign _EVAL_157 = ~_EVAL_126;
  assign _EVAL_115 = _EVAL_32 | _EVAL_1;
  assign _EVAL_250 = _EVAL_9 & _EVAL_16;
  assign _EVAL_215 = _EVAL_6 <= 3'h2;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_35 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_40 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_65 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_79 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_96 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_107 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_125 = _RAND_6[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_142 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_160 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_180 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_192 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_198 = _RAND_11[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_206 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_249 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_4) begin
    if (_EVAL_1) begin
      _EVAL_35 <= 1'h0;
    end else if (_EVAL_246) begin
      if (_EVAL_92) begin
        _EVAL_35 <= 1'h0;
      end else begin
        _EVAL_35 <= _EVAL_165;
      end
    end
    if (_EVAL_224) begin
      _EVAL_40 <= _EVAL_14;
    end
    if (_EVAL_1) begin
      _EVAL_65 <= 32'h0;
    end else if (_EVAL_100) begin
      _EVAL_65 <= 32'h0;
    end else begin
      _EVAL_65 <= _EVAL_154;
    end
    if (_EVAL_39) begin
      _EVAL_79 <= _EVAL_0;
    end
    if (_EVAL_224) begin
      _EVAL_96 <= _EVAL_6;
    end
    if (_EVAL_1) begin
      _EVAL_107 <= 1'h0;
    end else if (_EVAL_95) begin
      if (_EVAL_73) begin
        _EVAL_107 <= 1'h0;
      end else begin
        _EVAL_107 <= _EVAL_113;
      end
    end
    if (_EVAL_224) begin
      _EVAL_125 <= _EVAL_12;
    end
    if (_EVAL_39) begin
      _EVAL_142 <= _EVAL_11;
    end
    if (_EVAL_1) begin
      _EVAL_160 <= 1'h0;
    end else if (_EVAL_246) begin
      if (_EVAL_120) begin
        _EVAL_160 <= 1'h0;
      end else begin
        _EVAL_160 <= _EVAL_43;
      end
    end
    if (_EVAL_1) begin
      _EVAL_180 <= 1'h0;
    end else if (_EVAL_95) begin
      if (_EVAL_247) begin
        _EVAL_180 <= 1'h0;
      end else begin
        _EVAL_180 <= _EVAL_169;
      end
    end
    if (_EVAL_39) begin
      _EVAL_192 <= _EVAL_7;
    end
    if (_EVAL_1) begin
      _EVAL_198 <= 5'h0;
    end else begin
      _EVAL_198 <= _EVAL_89;
    end
    if (_EVAL_224) begin
      _EVAL_206 <= _EVAL_5;
    end
    if (_EVAL_224) begin
      _EVAL_249 <= _EVAL_3;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9356bc2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_31) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(757f155c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b4fee1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e300bdb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64aae1ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0fc3b6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7a11a07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb069a2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(194ed0d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a636e42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72165444)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac9c69ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e14230a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f82e3cc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cf76e6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(289149f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d2b36dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(738209ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8d75ac0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62ea902b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(caa5bab8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58c21f09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79452b41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d60ef20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccdd6f9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3cefdb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c53029d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92a34d8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70514dc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c94407e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9541a3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2a1ee35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc62aa3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ff3f45e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_31) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12f9d1d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61de9097)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_15) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(397ed70f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7f08a76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ca04690)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16f3ee8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14a41ec2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_31) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b63e85f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d500ede)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bda6277)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca3441b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f5863b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(882804f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a2c315)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22e8c74b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78532197)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d30563)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5e090b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e51ca1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6bcb29c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40a7a57f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9a84122)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73b33913)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4be6f6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bbba453)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a83fce0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b983b296)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b9f0454)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1bcb1e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_31) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7119e099)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_31) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae2f21ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69fce9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29551457)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_15) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf00dc2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d63c4e2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61a97c6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41e91bca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_31) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f900532)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cadf2d00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
