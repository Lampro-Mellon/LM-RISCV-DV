//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_51(
  input  [2:0]  _EVAL,
  output        _EVAL_0,
  input  [31:0] _EVAL_1,
  output        _EVAL_2,
  output [2:0]  _EVAL_3,
  output        _EVAL_4,
  output        _EVAL_5,
  input         _EVAL_6,
  output        _EVAL_7,
  input         _EVAL_8,
  output        _EVAL_9,
  output        _EVAL_10,
  output        _EVAL_11,
  output        _EVAL_12,
  output        _EVAL_13,
  input  [31:0] _EVAL_14,
  output [3:0]  _EVAL_15,
  input  [3:0]  _EVAL_16,
  input  [1:0]  _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19,
  input         _EVAL_20,
  input  [3:0]  _EVAL_21,
  input         _EVAL_22,
  output [31:0] _EVAL_23,
  input         _EVAL_24,
  output [3:0]  _EVAL_25,
  output [2:0]  _EVAL_26,
  input  [1:0]  _EVAL_27,
  output [31:0] _EVAL_28,
  output [31:0] _EVAL_29,
  input         _EVAL_30,
  input  [31:0] _EVAL_31,
  input  [2:0]  _EVAL_32,
  output        _EVAL_33,
  output        _EVAL_34,
  input  [2:0]  _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  input         _EVAL_38
);
  wire [2:0] fixer__EVAL;
  wire  fixer__EVAL_0;
  wire  fixer__EVAL_1;
  wire [31:0] fixer__EVAL_2;
  wire  fixer__EVAL_3;
  wire  fixer__EVAL_4;
  wire [2:0] fixer__EVAL_5;
  wire  fixer__EVAL_6;
  wire [31:0] fixer__EVAL_7;
  wire [3:0] fixer__EVAL_8;
  wire  fixer__EVAL_9;
  wire  fixer__EVAL_10;
  wire  fixer__EVAL_11;
  wire  fixer__EVAL_12;
  wire  fixer__EVAL_13;
  wire [31:0] fixer__EVAL_14;
  wire  fixer__EVAL_15;
  wire  fixer__EVAL_16;
  wire  fixer__EVAL_17;
  wire  fixer__EVAL_18;
  wire  fixer__EVAL_19;
  wire  fixer__EVAL_20;
  wire  fixer__EVAL_21;
  wire  fixer__EVAL_22;
  wire  fixer__EVAL_23;
  wire  fixer__EVAL_24;
  wire  fixer__EVAL_25;
  wire [3:0] fixer__EVAL_26;
  wire  fixer__EVAL_27;
  wire  fixer__EVAL_28;
  wire [31:0] fixer__EVAL_29;
  wire  fixer__EVAL_30;
  wire [2:0] fixer__EVAL_31;
  wire [2:0] fixer__EVAL_32;
  wire [1:0] fixer__EVAL_33;
  wire  fixer__EVAL_34;
  wire  fixer__EVAL_35;
  wire [3:0] fixer__EVAL_36;
  wire [1:0] fixer__EVAL_37;
  wire  fixer__EVAL_38;
  wire [3:0] fixer__EVAL_39;
  wire  fixer__EVAL_40;
  wire [31:0] fixer__EVAL_41;
  wire  fixer__EVAL_42;
  wire  fixer__EVAL_43;
  wire [3:0] fixer__EVAL_44;
  wire [3:0] fixer__EVAL_45;
  wire [31:0] fixer__EVAL_46;
  wire  buffer__EVAL;
  wire  buffer__EVAL_0;
  wire [2:0] buffer__EVAL_1;
  wire  buffer__EVAL_2;
  wire  buffer__EVAL_3;
  wire  buffer__EVAL_4;
  wire  buffer__EVAL_5;
  wire  buffer__EVAL_6;
  wire [31:0] buffer__EVAL_7;
  wire  buffer__EVAL_8;
  wire  buffer__EVAL_9;
  wire [3:0] buffer__EVAL_10;
  wire  buffer__EVAL_11;
  wire [31:0] buffer__EVAL_12;
  wire [31:0] buffer__EVAL_13;
  wire  buffer__EVAL_14;
  wire  buffer__EVAL_15;
  wire  buffer__EVAL_16;
  wire  buffer__EVAL_17;
  wire [31:0] buffer__EVAL_18;
  wire  buffer__EVAL_19;
  wire [3:0] buffer__EVAL_20;
  wire  buffer__EVAL_21;
  wire  buffer__EVAL_22;
  wire [31:0] buffer__EVAL_23;
  wire  buffer__EVAL_24;
  wire [3:0] buffer__EVAL_25;
  wire  buffer__EVAL_26;
  wire  buffer__EVAL_27;
  wire  buffer__EVAL_28;
  wire  buffer__EVAL_29;
  wire [31:0] buffer__EVAL_30;
  wire [1:0] buffer__EVAL_31;
  wire [3:0] buffer__EVAL_32;
  wire  buffer__EVAL_33;
  wire [2:0] buffer__EVAL_34;
  wire [3:0] buffer__EVAL_35;
  wire [3:0] buffer__EVAL_36;
  wire  buffer__EVAL_37;
  wire [2:0] buffer__EVAL_38;
  wire [2:0] buffer__EVAL_39;
  wire  buffer__EVAL_40;
  wire [2:0] buffer__EVAL_41;
  wire  buffer__EVAL_42;
  wire  buffer__EVAL_43;
  wire  buffer__EVAL_44;
  wire  buffer__EVAL_45;
  wire [1:0] buffer__EVAL_46;
  wire  buffer__EVAL_47;
  wire  buffer__EVAL_48;
  wire  buffer__EVAL_49;
  wire  ahb2tl__EVAL;
  wire  ahb2tl__EVAL_0;
  wire  ahb2tl__EVAL_1;
  wire  ahb2tl__EVAL_2;
  wire  ahb2tl__EVAL_3;
  wire [1:0] ahb2tl__EVAL_4;
  wire [31:0] ahb2tl__EVAL_5;
  wire [2:0] ahb2tl__EVAL_6;
  wire  ahb2tl__EVAL_7;
  wire [3:0] ahb2tl__EVAL_8;
  wire  ahb2tl__EVAL_9;
  wire [2:0] ahb2tl__EVAL_10;
  wire [31:0] ahb2tl__EVAL_11;
  wire  ahb2tl__EVAL_12;
  wire  ahb2tl__EVAL_13;
  wire  ahb2tl__EVAL_14;
  wire  ahb2tl__EVAL_15;
  wire  ahb2tl__EVAL_16;
  wire  ahb2tl__EVAL_17;
  wire [31:0] ahb2tl__EVAL_18;
  wire [31:0] ahb2tl__EVAL_19;
  wire  ahb2tl__EVAL_20;
  wire [2:0] ahb2tl__EVAL_21;
  wire  ahb2tl__EVAL_22;
  wire  ahb2tl__EVAL_23;
  wire [3:0] ahb2tl__EVAL_24;
  wire  ahb2tl__EVAL_25;
  wire  ahb2tl__EVAL_26;
  wire [3:0] ahb2tl__EVAL_27;
  wire [31:0] ahb2tl__EVAL_28;
  wire [31:0] ahb2tl__EVAL_29;
  wire  ahb2tl__EVAL_30;
  wire  widget__EVAL;
  wire  widget__EVAL_0;
  wire  widget__EVAL_1;
  wire [31:0] widget__EVAL_2;
  wire [31:0] widget__EVAL_3;
  wire  widget__EVAL_4;
  wire [3:0] widget__EVAL_5;
  wire  widget__EVAL_6;
  wire  widget__EVAL_7;
  wire  widget__EVAL_8;
  wire [1:0] widget__EVAL_9;
  wire  widget__EVAL_10;
  wire [2:0] widget__EVAL_11;
  wire [3:0] widget__EVAL_12;
  wire [2:0] widget__EVAL_13;
  wire  widget__EVAL_14;
  wire  widget__EVAL_15;
  wire  widget__EVAL_16;
  wire  widget__EVAL_17;
  wire [31:0] widget__EVAL_18;
  wire [31:0] widget__EVAL_19;
  wire  widget__EVAL_20;
  wire  widget__EVAL_21;
  wire  widget__EVAL_22;
  wire  widget__EVAL_23;
  wire  widget__EVAL_24;
  wire  widget__EVAL_25;
  wire [31:0] widget__EVAL_26;
  wire  widget__EVAL_27;
  wire  widget__EVAL_28;
  wire [3:0] widget__EVAL_29;
  wire  widget__EVAL_30;
  wire  widget__EVAL_31;
  wire  widget__EVAL_32;
  wire  widget__EVAL_33;
  wire  widget__EVAL_34;
  wire  widget__EVAL_35;
  wire [3:0] widget__EVAL_36;
  wire [2:0] widget__EVAL_37;
  wire  widget__EVAL_38;
  wire [3:0] widget__EVAL_39;
  wire  widget__EVAL_40;
  wire [31:0] widget__EVAL_41;
  _EVAL_47 fixer (
    ._EVAL(fixer__EVAL),
    ._EVAL_0(fixer__EVAL_0),
    ._EVAL_1(fixer__EVAL_1),
    ._EVAL_2(fixer__EVAL_2),
    ._EVAL_3(fixer__EVAL_3),
    ._EVAL_4(fixer__EVAL_4),
    ._EVAL_5(fixer__EVAL_5),
    ._EVAL_6(fixer__EVAL_6),
    ._EVAL_7(fixer__EVAL_7),
    ._EVAL_8(fixer__EVAL_8),
    ._EVAL_9(fixer__EVAL_9),
    ._EVAL_10(fixer__EVAL_10),
    ._EVAL_11(fixer__EVAL_11),
    ._EVAL_12(fixer__EVAL_12),
    ._EVAL_13(fixer__EVAL_13),
    ._EVAL_14(fixer__EVAL_14),
    ._EVAL_15(fixer__EVAL_15),
    ._EVAL_16(fixer__EVAL_16),
    ._EVAL_17(fixer__EVAL_17),
    ._EVAL_18(fixer__EVAL_18),
    ._EVAL_19(fixer__EVAL_19),
    ._EVAL_20(fixer__EVAL_20),
    ._EVAL_21(fixer__EVAL_21),
    ._EVAL_22(fixer__EVAL_22),
    ._EVAL_23(fixer__EVAL_23),
    ._EVAL_24(fixer__EVAL_24),
    ._EVAL_25(fixer__EVAL_25),
    ._EVAL_26(fixer__EVAL_26),
    ._EVAL_27(fixer__EVAL_27),
    ._EVAL_28(fixer__EVAL_28),
    ._EVAL_29(fixer__EVAL_29),
    ._EVAL_30(fixer__EVAL_30),
    ._EVAL_31(fixer__EVAL_31),
    ._EVAL_32(fixer__EVAL_32),
    ._EVAL_33(fixer__EVAL_33),
    ._EVAL_34(fixer__EVAL_34),
    ._EVAL_35(fixer__EVAL_35),
    ._EVAL_36(fixer__EVAL_36),
    ._EVAL_37(fixer__EVAL_37),
    ._EVAL_38(fixer__EVAL_38),
    ._EVAL_39(fixer__EVAL_39),
    ._EVAL_40(fixer__EVAL_40),
    ._EVAL_41(fixer__EVAL_41),
    ._EVAL_42(fixer__EVAL_42),
    ._EVAL_43(fixer__EVAL_43),
    ._EVAL_44(fixer__EVAL_44),
    ._EVAL_45(fixer__EVAL_45),
    ._EVAL_46(fixer__EVAL_46)
  );
  _EVAL_45 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32),
    ._EVAL_33(buffer__EVAL_33),
    ._EVAL_34(buffer__EVAL_34),
    ._EVAL_35(buffer__EVAL_35),
    ._EVAL_36(buffer__EVAL_36),
    ._EVAL_37(buffer__EVAL_37),
    ._EVAL_38(buffer__EVAL_38),
    ._EVAL_39(buffer__EVAL_39),
    ._EVAL_40(buffer__EVAL_40),
    ._EVAL_41(buffer__EVAL_41),
    ._EVAL_42(buffer__EVAL_42),
    ._EVAL_43(buffer__EVAL_43),
    ._EVAL_44(buffer__EVAL_44),
    ._EVAL_45(buffer__EVAL_45),
    ._EVAL_46(buffer__EVAL_46),
    ._EVAL_47(buffer__EVAL_47),
    ._EVAL_48(buffer__EVAL_48),
    ._EVAL_49(buffer__EVAL_49)
  );
  _EVAL_50 ahb2tl (
    ._EVAL(ahb2tl__EVAL),
    ._EVAL_0(ahb2tl__EVAL_0),
    ._EVAL_1(ahb2tl__EVAL_1),
    ._EVAL_2(ahb2tl__EVAL_2),
    ._EVAL_3(ahb2tl__EVAL_3),
    ._EVAL_4(ahb2tl__EVAL_4),
    ._EVAL_5(ahb2tl__EVAL_5),
    ._EVAL_6(ahb2tl__EVAL_6),
    ._EVAL_7(ahb2tl__EVAL_7),
    ._EVAL_8(ahb2tl__EVAL_8),
    ._EVAL_9(ahb2tl__EVAL_9),
    ._EVAL_10(ahb2tl__EVAL_10),
    ._EVAL_11(ahb2tl__EVAL_11),
    ._EVAL_12(ahb2tl__EVAL_12),
    ._EVAL_13(ahb2tl__EVAL_13),
    ._EVAL_14(ahb2tl__EVAL_14),
    ._EVAL_15(ahb2tl__EVAL_15),
    ._EVAL_16(ahb2tl__EVAL_16),
    ._EVAL_17(ahb2tl__EVAL_17),
    ._EVAL_18(ahb2tl__EVAL_18),
    ._EVAL_19(ahb2tl__EVAL_19),
    ._EVAL_20(ahb2tl__EVAL_20),
    ._EVAL_21(ahb2tl__EVAL_21),
    ._EVAL_22(ahb2tl__EVAL_22),
    ._EVAL_23(ahb2tl__EVAL_23),
    ._EVAL_24(ahb2tl__EVAL_24),
    ._EVAL_25(ahb2tl__EVAL_25),
    ._EVAL_26(ahb2tl__EVAL_26),
    ._EVAL_27(ahb2tl__EVAL_27),
    ._EVAL_28(ahb2tl__EVAL_28),
    ._EVAL_29(ahb2tl__EVAL_29),
    ._EVAL_30(ahb2tl__EVAL_30)
  );
  _EVAL_49 widget (
    ._EVAL(widget__EVAL),
    ._EVAL_0(widget__EVAL_0),
    ._EVAL_1(widget__EVAL_1),
    ._EVAL_2(widget__EVAL_2),
    ._EVAL_3(widget__EVAL_3),
    ._EVAL_4(widget__EVAL_4),
    ._EVAL_5(widget__EVAL_5),
    ._EVAL_6(widget__EVAL_6),
    ._EVAL_7(widget__EVAL_7),
    ._EVAL_8(widget__EVAL_8),
    ._EVAL_9(widget__EVAL_9),
    ._EVAL_10(widget__EVAL_10),
    ._EVAL_11(widget__EVAL_11),
    ._EVAL_12(widget__EVAL_12),
    ._EVAL_13(widget__EVAL_13),
    ._EVAL_14(widget__EVAL_14),
    ._EVAL_15(widget__EVAL_15),
    ._EVAL_16(widget__EVAL_16),
    ._EVAL_17(widget__EVAL_17),
    ._EVAL_18(widget__EVAL_18),
    ._EVAL_19(widget__EVAL_19),
    ._EVAL_20(widget__EVAL_20),
    ._EVAL_21(widget__EVAL_21),
    ._EVAL_22(widget__EVAL_22),
    ._EVAL_23(widget__EVAL_23),
    ._EVAL_24(widget__EVAL_24),
    ._EVAL_25(widget__EVAL_25),
    ._EVAL_26(widget__EVAL_26),
    ._EVAL_27(widget__EVAL_27),
    ._EVAL_28(widget__EVAL_28),
    ._EVAL_29(widget__EVAL_29),
    ._EVAL_30(widget__EVAL_30),
    ._EVAL_31(widget__EVAL_31),
    ._EVAL_32(widget__EVAL_32),
    ._EVAL_33(widget__EVAL_33),
    ._EVAL_34(widget__EVAL_34),
    ._EVAL_35(widget__EVAL_35),
    ._EVAL_36(widget__EVAL_36),
    ._EVAL_37(widget__EVAL_37),
    ._EVAL_38(widget__EVAL_38),
    ._EVAL_39(widget__EVAL_39),
    ._EVAL_40(widget__EVAL_40),
    ._EVAL_41(widget__EVAL_41)
  );
  assign _EVAL_4 = ahb2tl__EVAL_7;
  assign ahb2tl__EVAL_21 = _EVAL;
  assign fixer__EVAL_11 = widget__EVAL_28;
  assign widget__EVAL_32 = ahb2tl__EVAL_23;
  assign widget__EVAL_21 = fixer__EVAL_10;
  assign buffer__EVAL_36 = _EVAL_16;
  assign ahb2tl__EVAL_27 = _EVAL_21;
  assign widget__EVAL_2 = ahb2tl__EVAL_11;
  assign fixer__EVAL_0 = buffer__EVAL_19;
  assign _EVAL_29 = ahb2tl__EVAL_29;
  assign _EVAL_23 = buffer__EVAL_13;
  assign fixer__EVAL_22 = widget__EVAL_7;
  assign buffer__EVAL_38 = fixer__EVAL_31;
  assign _EVAL_13 = buffer__EVAL_37;
  assign fixer__EVAL_19 = widget__EVAL_35;
  assign widget__EVAL_11 = ahb2tl__EVAL_6;
  assign widget__EVAL_34 = _EVAL_36;
  assign buffer__EVAL_46 = _EVAL_27;
  assign _EVAL_26 = buffer__EVAL_1;
  assign widget__EVAL_3 = ahb2tl__EVAL_18;
  assign fixer__EVAL_25 = buffer__EVAL_5;
  assign widget__EVAL_10 = ahb2tl__EVAL_13;
  assign _EVAL_18 = buffer__EVAL_4;
  assign buffer__EVAL_34 = _EVAL_32;
  assign widget__EVAL_33 = ahb2tl__EVAL_14;
  assign _EVAL_12 = buffer__EVAL_45;
  assign _EVAL_28 = buffer__EVAL_30;
  assign widget__EVAL_12 = fixer__EVAL_44;
  assign fixer__EVAL_17 = widget__EVAL_14;
  assign buffer__EVAL_6 = _EVAL_30;
  assign fixer__EVAL_32 = buffer__EVAL_41;
  assign buffer__EVAL_18 = fixer__EVAL_2;
  assign _EVAL_5 = buffer__EVAL_49;
  assign widget__EVAL_0 = ahb2tl__EVAL_17;
  assign fixer__EVAL_6 = buffer__EVAL_11;
  assign ahb2tl__EVAL_5 = _EVAL_14;
  assign fixer__EVAL_41 = buffer__EVAL_7;
  assign ahb2tl__EVAL_20 = _EVAL_37;
  assign buffer__EVAL_15 = _EVAL_36;
  assign buffer__EVAL_17 = _EVAL_24;
  assign fixer__EVAL_39 = widget__EVAL_5;
  assign widget__EVAL_6 = fixer__EVAL_4;
  assign _EVAL_9 = buffer__EVAL_29;
  assign _EVAL_33 = buffer__EVAL_42;
  assign fixer__EVAL_8 = widget__EVAL_36;
  assign widget__EVAL_29 = ahb2tl__EVAL_24;
  assign _EVAL_2 = ahb2tl__EVAL_22;
  assign widget__EVAL_15 = fixer__EVAL_21;
  assign ahb2tl__EVAL_3 = _EVAL_6;
  assign _EVAL_34 = buffer__EVAL_40;
  assign ahb2tl__EVAL_10 = _EVAL_35;
  assign widget__EVAL = ahb2tl__EVAL_2;
  assign fixer__EVAL_12 = _EVAL_20;
  assign buffer__EVAL_2 = fixer__EVAL_24;
  assign fixer__EVAL_37 = buffer__EVAL_31;
  assign buffer__EVAL_24 = fixer__EVAL_20;
  assign buffer__EVAL_0 = fixer__EVAL_30;
  assign fixer__EVAL_29 = widget__EVAL_18;
  assign ahb2tl__EVAL_4 = _EVAL_17;
  assign fixer__EVAL_15 = buffer__EVAL_21;
  assign widget__EVAL_13 = fixer__EVAL;
  assign ahb2tl__EVAL_1 = _EVAL_20;
  assign fixer__EVAL_18 = widget__EVAL_25;
  assign fixer__EVAL_36 = buffer__EVAL_35;
  assign fixer__EVAL_34 = _EVAL_36;
  assign widget__EVAL_22 = fixer__EVAL_3;
  assign _EVAL_15 = buffer__EVAL_25;
  assign widget__EVAL_24 = ahb2tl__EVAL_15;
  assign buffer__EVAL_14 = _EVAL_8;
  assign buffer__EVAL_32 = fixer__EVAL_26;
  assign _EVAL_11 = buffer__EVAL_44;
  assign _EVAL_0 = buffer__EVAL_22;
  assign widget__EVAL_1 = _EVAL_20;
  assign buffer__EVAL_47 = fixer__EVAL_43;
  assign buffer__EVAL_26 = fixer__EVAL_13;
  assign ahb2tl__EVAL_9 = widget__EVAL_16;
  assign fixer__EVAL_42 = widget__EVAL_27;
  assign buffer__EVAL_27 = fixer__EVAL_1;
  assign fixer__EVAL_5 = widget__EVAL_37;
  assign ahb2tl__EVAL_19 = _EVAL_31;
  assign buffer__EVAL_8 = _EVAL_38;
  assign buffer__EVAL_48 = fixer__EVAL_28;
  assign ahb2tl__EVAL_0 = widget__EVAL_30;
  assign fixer__EVAL_38 = widget__EVAL_17;
  assign fixer__EVAL_40 = widget__EVAL_8;
  assign widget__EVAL_19 = fixer__EVAL_7;
  assign widget__EVAL_38 = fixer__EVAL_9;
  assign widget__EVAL_31 = ahb2tl__EVAL_25;
  assign fixer__EVAL_23 = buffer__EVAL_33;
  assign ahb2tl__EVAL = _EVAL_19;
  assign buffer__EVAL_12 = fixer__EVAL_46;
  assign buffer__EVAL_3 = _EVAL_22;
  assign ahb2tl__EVAL_30 = widget__EVAL_4;
  assign fixer__EVAL_35 = buffer__EVAL_28;
  assign buffer__EVAL_43 = fixer__EVAL_16;
  assign _EVAL_3 = buffer__EVAL_39;
  assign _EVAL_7 = buffer__EVAL_9;
  assign buffer__EVAL_16 = _EVAL_20;
  assign widget__EVAL_9 = fixer__EVAL_33;
  assign ahb2tl__EVAL_16 = _EVAL_36;
  assign _EVAL_10 = buffer__EVAL;
  assign buffer__EVAL_23 = _EVAL_1;
  assign _EVAL_25 = buffer__EVAL_20;
  assign widget__EVAL_20 = fixer__EVAL_27;
  assign widget__EVAL_23 = ahb2tl__EVAL_26;
  assign buffer__EVAL_10 = fixer__EVAL_45;
  assign ahb2tl__EVAL_12 = widget__EVAL_40;
  assign fixer__EVAL_14 = widget__EVAL_26;
  assign ahb2tl__EVAL_28 = widget__EVAL_41;
  assign widget__EVAL_39 = ahb2tl__EVAL_8;
endmodule
