//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_41(
  input         _EVAL,
  output        _EVAL_0,
  output        _EVAL_1,
  input  [3:0]  _EVAL_2,
  output [1:0]  _EVAL_3,
  output        _EVAL_4,
  output        _EVAL_5,
  input         _EVAL_6,
  output        _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  output        _EVAL_10,
  output [2:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [1:0]  _EVAL_14,
  output [2:0]  _EVAL_15,
  input  [31:0] _EVAL_16,
  output        _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19,
  output        _EVAL_20,
  output        _EVAL_21,
  output        _EVAL_22,
  output        _EVAL_23,
  output        _EVAL_24,
  input  [31:0] _EVAL_25,
  output [3:0]  _EVAL_26,
  output        _EVAL_27,
  output [31:0] _EVAL_28,
  input  [3:0]  _EVAL_29,
  output [2:0]  _EVAL_30,
  input  [31:0] _EVAL_31,
  input         _EVAL_32,
  output [3:0]  _EVAL_33,
  input         _EVAL_34,
  output        _EVAL_35,
  output [31:0] _EVAL_36,
  input         _EVAL_37,
  input         _EVAL_38,
  output        _EVAL_39,
  input         _EVAL_40,
  input  [3:0]  _EVAL_41,
  output [3:0]  _EVAL_42,
  input         _EVAL_43,
  input         _EVAL_44,
  input  [2:0]  _EVAL_45,
  input  [2:0]  _EVAL_46,
  input         _EVAL_47,
  input         _EVAL_48,
  input         _EVAL_49,
  input         _EVAL_50,
  input         _EVAL_51,
  output [31:0] _EVAL_52
);
  assign _EVAL_11 = _EVAL_46;
  assign _EVAL_0 = _EVAL_13;
  assign _EVAL_10 = _EVAL_44;
  assign _EVAL_26 = _EVAL_2;
  assign _EVAL_23 = _EVAL_47;
  assign _EVAL_30 = _EVAL_9;
  assign _EVAL_7 = _EVAL_51;
  assign _EVAL_27 = _EVAL_6;
  assign _EVAL_52 = _EVAL_31;
  assign _EVAL_17 = _EVAL_43;
  assign _EVAL_36 = _EVAL_16;
  assign _EVAL_28 = _EVAL_25;
  assign _EVAL_42 = _EVAL_41;
  assign _EVAL_33 = _EVAL_29;
  assign _EVAL_39 = _EVAL;
  assign _EVAL_5 = _EVAL_50;
  assign _EVAL_20 = _EVAL_37;
  assign _EVAL_22 = _EVAL_38;
  assign _EVAL_4 = _EVAL_32;
  assign _EVAL_35 = _EVAL_19;
  assign _EVAL_1 = _EVAL_48;
  assign _EVAL_18 = _EVAL_49;
  assign _EVAL_15 = _EVAL_45;
  assign _EVAL_3 = _EVAL_14;
  assign _EVAL_24 = _EVAL_8;
  assign _EVAL_21 = _EVAL_40;
endmodule
