//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_123_assert(
  input        _EVAL,
  input        _EVAL_0,
  input        _EVAL_1,
  input        _EVAL_2,
  input        _EVAL_3,
  input        _EVAL_4,
  input        _EVAL_5,
  input  [1:0] _EVAL_6,
  input  [2:0] _EVAL_7,
  input        _EVAL_8,
  input  [1:0] _EVAL_9,
  input        _EVAL_10,
  input        _EVAL_11,
  input  [3:0] _EVAL_12,
  input  [2:0] _EVAL_13,
  input  [8:0] _EVAL_14
);
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  reg [1:0] _EVAL_21;
  reg [31:0] _RAND_0;
  wire  _EVAL_22;
  wire [9:0] _EVAL_23;
  reg [31:0] _EVAL_24;
  reg [31:0] _RAND_1;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire [8:0] _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire [9:0] _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire [9:0] _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  reg [1:0] _EVAL_44;
  reg [31:0] _RAND_2;
  wire  _EVAL_45;
  wire [8:0] _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  reg  _EVAL_53;
  reg [31:0] _RAND_3;
  reg [8:0] _EVAL_54;
  reg [31:0] _RAND_4;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire [1:0] _EVAL_65;
  wire [1:0] _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire [9:0] _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire [1:0] _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire [9:0] _EVAL_79;
  wire  _EVAL_80;
  wire [32:0] _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  reg  _EVAL_89;
  reg [31:0] _RAND_5;
  wire [9:0] _EVAL_90;
  wire  _EVAL_91;
  wire [8:0] _EVAL_92;
  wire  _EVAL_93;
  reg  _EVAL_94;
  reg [31:0] _RAND_6;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire [9:0] _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  reg  _EVAL_102;
  reg [31:0] _RAND_7;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  reg  _EVAL_107;
  reg [31:0] _RAND_8;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire [8:0] _EVAL_117;
  wire  _EVAL_118;
  wire [9:0] _EVAL_119;
  wire [1:0] _EVAL_120;
  wire  _EVAL_121;
  wire [9:0] _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire [9:0] _EVAL_130;
  wire [9:0] _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire [3:0] _EVAL_137;
  reg [2:0] _EVAL_138;
  reg [31:0] _RAND_9;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire [9:0] _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire [9:0] _EVAL_156;
  wire  _EVAL_157;
  wire [1:0] _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire [9:0] _EVAL_163;
  wire [9:0] _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire [9:0] _EVAL_175;
  wire  _EVAL_177;
  wire [8:0] _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  reg [2:0] _EVAL_181;
  reg [31:0] _RAND_10;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire [1:0] _EVAL_184;
  wire  _EVAL_185;
  wire [1:0] _EVAL_186;
  wire  _EVAL_187;
  reg  _EVAL_188;
  reg [31:0] _RAND_11;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire [8:0] _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  reg  _EVAL_201;
  reg [31:0] _RAND_12;
  wire  _EVAL_202;
  wire [9:0] _EVAL_203;
  reg  _EVAL_204;
  reg [31:0] _RAND_13;
  wire [31:0] _EVAL_205;
  wire [9:0] _EVAL_206;
  wire  _EVAL_207;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_25 = _EVAL_9 == _EVAL_21;
  assign _EVAL_158 = _EVAL_204 - 1'h1;
  assign _EVAL_47 = _EVAL_115 | _EVAL_141;
  assign _EVAL_23 = $signed(_EVAL_130) & -10'sh20;
  assign _EVAL_169 = ~_EVAL_199;
  assign _EVAL_154 = _EVAL_13 == 3'h4;
  assign _EVAL_127 = _EVAL_147 | _EVAL_70;
  assign _EVAL_190 = _EVAL_51 | _EVAL_70;
  assign _EVAL_28 = _EVAL_207 | _EVAL_70;
  assign _EVAL_40 = _EVAL_50 | _EVAL_70;
  assign _EVAL_142 = _EVAL_4 & _EVAL_32;
  assign _EVAL_131 = {1'b0,$signed(_EVAL_46)};
  assign _EVAL_133 = _EVAL_120[0];
  assign _EVAL_88 = _EVAL_150 & _EVAL_68;
  assign _EVAL_39 = ~_EVAL_15;
  assign _EVAL_81 = _EVAL_24 + 32'h1;
  assign _EVAL_67 = _EVAL_123 | _EVAL_70;
  assign _EVAL_71 = $signed(_EVAL_97) & -10'sh80;
  assign _EVAL_119 = $signed(_EVAL_164) & -10'sh40;
  assign _EVAL_145 = _EVAL_1 & _EVAL_75;
  assign _EVAL_35 = $signed(_EVAL_131) & -10'sh4;
  assign _EVAL_182 = ~_EVAL_192;
  assign _EVAL_153 = $signed(_EVAL_163) == 10'sh0;
  assign _EVAL_26 = $signed(_EVAL_175) == 10'sh0;
  assign _EVAL_174 = ~_EVAL_67;
  assign _EVAL_120 = _EVAL_107 - 1'h1;
  assign _EVAL_121 = _EVAL_196 | _EVAL_70;
  assign _EVAL_22 = _EVAL_1 & _EVAL_139;
  assign _EVAL_159 = ~_EVAL_135;
  assign _EVAL_96 = ~_EVAL_31;
  assign _EVAL_78 = _EVAL_43 | _EVAL_70;
  assign _EVAL_69 = _EVAL_171 | _EVAL_70;
  assign _EVAL_61 = _EVAL_4 & _EVAL_60;
  assign _EVAL_74 = ~_EVAL_148;
  assign _EVAL_65 = _EVAL_91 ? 2'h1 : 2'h0;
  assign _EVAL_90 = _EVAL_23;
  assign _EVAL_27 = _EVAL_14 ^ 9'h60;
  assign _EVAL_139 = _EVAL_13 == 3'h0;
  assign _EVAL_29 = _EVAL_7 <= 3'h6;
  assign _EVAL_198 = ~_EVAL_127;
  assign _EVAL_196 = _EVAL_50 | _EVAL_0;
  assign _EVAL_203 = $signed(_EVAL_144) & -10'sh18;
  assign _EVAL_178 = _EVAL_14 ^ 9'h48;
  assign _EVAL_197 = _EVAL_14 & 9'h3;
  assign _EVAL_117 = _EVAL_14 ^ 9'h100;
  assign _EVAL_103 = ~_EVAL_183;
  assign _EVAL_114 = ~_EVAL_190;
  assign _EVAL_134 = _EVAL_1 & _EVAL_20;
  assign _EVAL_57 = ~_EVAL_172;
  assign _EVAL_186 = 2'h1 << _EVAL_2;
  assign _EVAL_34 = _EVAL_157 | _EVAL_194;
  assign _EVAL_52 = _EVAL & _EVAL_4;
  assign _EVAL_163 = _EVAL_35;
  assign _EVAL_143 = _EVAL_13 == 3'h1;
  assign _EVAL_195 = ~_EVAL_68;
  assign _EVAL_165 = $signed(_EVAL_90) == 10'sh0;
  assign _EVAL_98 = _EVAL_7 == 3'h0;
  assign _EVAL_42 = _EVAL_184[0];
  assign _EVAL_16 = $signed(_EVAL_41) == 10'sh0;
  assign _EVAL_184 = _EVAL_53 - 1'h1;
  assign _EVAL_101 = ~_EVAL_58;
  assign _EVAL_49 = ~_EVAL_40;
  assign _EVAL_51 = _EVAL_12 == 4'hf;
  assign _EVAL_141 = $signed(_EVAL_156) == 10'sh0;
  assign _EVAL_43 = _EVAL_14 == _EVAL_54;
  assign _EVAL_83 = _EVAL_137 == 4'h0;
  assign _EVAL_189 = ~_EVAL_121;
  assign _EVAL_173 = _EVAL_86 | _EVAL_70;
  assign _EVAL_126 = _EVAL_197 == 9'h0;
  assign _EVAL_147 = _EVAL_170 >> _EVAL_2;
  assign _EVAL_193 = ~_EVAL_102;
  assign _EVAL_68 = ~_EVAL_204;
  assign _EVAL_77 = ~_EVAL_200;
  assign _EVAL_192 = _EVAL_136 | _EVAL_70;
  assign _EVAL_112 = _EVAL_106 | _EVAL_70;
  assign _EVAL_125 = _EVAL_4 & _EVAL_30;
  assign _EVAL_124 = _EVAL_65[0];
  assign _EVAL_109 = _EVAL_1 & _EVAL_80;
  assign _EVAL_177 = ~_EVAL_69;
  assign _EVAL_38 = ~_EVAL_70;
  assign _EVAL_150 = _EVAL_10 & _EVAL_1;
  assign _EVAL_137 = ~_EVAL_12;
  assign _EVAL_136 = _EVAL_9 >= 2'h2;
  assign _EVAL_63 = _EVAL_7 == 3'h4;
  assign _EVAL_31 = _EVAL_47 | _EVAL_70;
  assign _EVAL_19 = _EVAL_150 | _EVAL_52;
  assign _EVAL_129 = _EVAL_161 | _EVAL_70;
  assign _EVAL_123 = _EVAL_6 == _EVAL_44;
  assign _EVAL_37 = ~_EVAL_53;
  assign _EVAL_166 = ~_EVAL_107;
  assign _EVAL_105 = _EVAL_29 | _EVAL_70;
  assign _EVAL_161 = ~_EVAL_0;
  assign _EVAL_172 = _EVAL_25 | _EVAL_70;
  assign _EVAL_18 = _EVAL_13 == 3'h5;
  assign _EVAL_194 = $signed(_EVAL_79) == 10'sh0;
  assign _EVAL_84 = ~_EVAL_99;
  assign _EVAL_55 = _EVAL_1 & _EVAL_195;
  assign _EVAL_140 = _EVAL_2 == _EVAL_94;
  assign _EVAL_59 = ~_EVAL_78;
  assign _EVAL_200 = _EVAL_149 | _EVAL_70;
  assign _EVAL_108 = _EVAL_1 & _EVAL_72;
  assign _EVAL_151 = _EVAL_6 == 2'h0;
  assign _EVAL_93 = plusarg_reader_out == 32'h0;
  assign _EVAL_70 = _EVAL_8;
  assign _EVAL_86 = ~_EVAL_2;
  assign _EVAL_62 = _EVAL_24 < plusarg_reader_out;
  assign _EVAL_157 = _EVAL_16 | _EVAL_153;
  assign _EVAL_15 = _EVAL_36 | _EVAL_70;
  assign _EVAL_156 = _EVAL_122;
  assign _EVAL_72 = _EVAL_13 == 3'h7;
  assign _EVAL_17 = _EVAL_4 & _EVAL_100;
  assign _EVAL_106 = _EVAL_7 == _EVAL_181;
  assign _EVAL_115 = _EVAL_167 | _EVAL_26;
  assign _EVAL_99 = _EVAL_126 | _EVAL_70;
  assign _EVAL_48 = _EVAL_132 | _EVAL_93;
  assign _EVAL_175 = _EVAL_71;
  assign _EVAL_36 = _EVAL_6 != 2'h2;
  assign _EVAL_183 = _EVAL_83 | _EVAL_70;
  assign _EVAL_128 = ~_EVAL_112;
  assign _EVAL_58 = _EVAL_66[0];
  assign _EVAL_202 = ~_EVAL_129;
  assign _EVAL_144 = {1'b0,$signed(_EVAL_178)};
  assign _EVAL_180 = _EVAL_188 | _EVAL_124;
  assign _EVAL_91 = _EVAL_150 & _EVAL_166;
  assign _EVAL_41 = _EVAL_119;
  assign _EVAL_168 = _EVAL_52 & _EVAL_37;
  assign _EVAL_80 = _EVAL_13 == 3'h2;
  assign _EVAL_46 = _EVAL_14 ^ 9'h44;
  assign _EVAL_162 = _EVAL_7 == 3'h1;
  assign _EVAL_187 = _EVAL_4 & _EVAL_63;
  assign _EVAL_199 = _EVAL_140 | _EVAL_70;
  assign _EVAL_104 = _EVAL_158[0];
  assign _EVAL_100 = _EVAL_7 == 3'h6;
  assign _EVAL_20 = _EVAL_13 == 3'h6;
  assign _EVAL_207 = _EVAL_48 | _EVAL_62;
  assign _EVAL_148 = _EVAL_132 | _EVAL_70;
  assign _EVAL_76 = _EVAL_102 - 1'h1;
  assign _EVAL_132 = ~_EVAL_188;
  assign _EVAL_118 = _EVAL_1 & _EVAL_143;
  assign _EVAL_97 = {1'b0,$signed(_EVAL_92)};
  assign _EVAL_92 = _EVAL_14 ^ 9'h80;
  assign _EVAL_130 = {1'b0,$signed(_EVAL_27)};
  assign _EVAL_205 = _EVAL_81[31:0];
  assign _EVAL_170 = _EVAL_124 | _EVAL_188;
  assign _EVAL_30 = _EVAL_7 == 3'h2;
  assign _EVAL_56 = ~_EVAL_100;
  assign _EVAL_75 = _EVAL_13 == 3'h3;
  assign _EVAL_33 = _EVAL_52 & _EVAL_193;
  assign _EVAL_66 = _EVAL_191 ? _EVAL_186 : 2'h0;
  assign _EVAL_122 = $signed(_EVAL_206) & -10'sh100;
  assign _EVAL_45 = _EVAL_179 | _EVAL_70;
  assign _EVAL_206 = {1'b0,$signed(_EVAL_117)};
  assign _EVAL_185 = ~_EVAL_105;
  assign _EVAL_155 = ~_EVAL_45;
  assign _EVAL_95 = ~_EVAL_173;
  assign _EVAL_191 = _EVAL_33 & _EVAL_56;
  assign _EVAL_149 = _EVAL_13 == _EVAL_138;
  assign _EVAL_60 = _EVAL_7 == 3'h5;
  assign _EVAL_164 = {1'b0,$signed(_EVAL_14)};
  assign _EVAL_73 = _EVAL_1 & _EVAL_154;
  assign _EVAL_167 = _EVAL_34 | _EVAL_165;
  assign _EVAL_110 = ~_EVAL_111;
  assign _EVAL_152 = _EVAL_1 & _EVAL_18;
  assign _EVAL_32 = ~_EVAL_37;
  assign _EVAL_135 = _EVAL_82 | _EVAL_70;
  assign _EVAL_50 = ~_EVAL_3;
  assign _EVAL_79 = _EVAL_203;
  assign _EVAL_179 = _EVAL_6 <= 2'h2;
  assign _EVAL_111 = _EVAL_151 | _EVAL_70;
  assign _EVAL_82 = _EVAL_3 == _EVAL_201;
  assign _EVAL_146 = _EVAL_76[0];
  assign _EVAL_85 = ~_EVAL_28;
  assign _EVAL_116 = _EVAL_4 & _EVAL_162;
  assign _EVAL_171 = _EVAL_11 == _EVAL_89;
  assign _EVAL_87 = _EVAL_4 & _EVAL_98;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_21 = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_24 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_44 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_53 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_54 = _RAND_4[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_89 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_94 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_102 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_107 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_138 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_181 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_188 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_201 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_204 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  if (_EVAL_8) begin
    _EVAL_24 = 32'h0;
  end
  if (_EVAL_8) begin
    _EVAL_53 = 1'h0;
  end
  if (_EVAL_8) begin
    _EVAL_102 = 1'h0;
  end
  if (_EVAL_8) begin
    _EVAL_107 = 1'h0;
  end
  if (_EVAL_8) begin
    _EVAL_188 = 1'h0;
  end
  if (_EVAL_8) begin
    _EVAL_204 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_5) begin
    if (_EVAL_168) begin
      _EVAL_21 <= _EVAL_9;
    end
    if (_EVAL_168) begin
      _EVAL_44 <= _EVAL_6;
    end
    if (_EVAL_88) begin
      _EVAL_54 <= _EVAL_14;
    end
    if (_EVAL_168) begin
      _EVAL_89 <= _EVAL_11;
    end
    if (_EVAL_168) begin
      _EVAL_94 <= _EVAL_2;
    end
    if (_EVAL_88) begin
      _EVAL_138 <= _EVAL_13;
    end
    if (_EVAL_168) begin
      _EVAL_181 <= _EVAL_7;
    end
    if (_EVAL_168) begin
      _EVAL_201 <= _EVAL_3;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5577e3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ea9e816)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(682dd615)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5cd13bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7ce340f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6264572)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d36ec8a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27f25775)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(868940fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e9a1d72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ecb0fb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e2f01f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b96f81b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19512b5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cffd24d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(254e24d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4b63298)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ef2feb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55f7620b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad6d1899)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9824f50d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e23f8298)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fb866c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9ef29e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46841f21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc3bbddb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cc37fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7e4fc26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba557f94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be997427)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee7bb1fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11952299)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a17eb4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6a9b46f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d89391e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(857e00ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb074361)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4c627cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb147ec3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff35720e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(270eb1de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75d00cc4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2332c1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1475e58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98e021df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(492f71c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2376447d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(370b8c91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cae3e3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bef6ae21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9582863)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75228d64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5ecdde1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2711a9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a739353)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38e64b79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac929197)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62a97ebd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c057339)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b590f093)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1d2cd03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84c2ab2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d03ea8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69395e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge _EVAL_5 or posedge _EVAL_8) begin
    if (_EVAL_8) begin
      _EVAL_24 <= 32'h0;
    end else if (_EVAL_19) begin
      _EVAL_24 <= 32'h0;
    end else begin
      _EVAL_24 <= _EVAL_205;
    end
  end
  always @(posedge _EVAL_5 or posedge _EVAL_8) begin
    if (_EVAL_8) begin
      _EVAL_53 <= 1'h0;
    end else if (_EVAL_52) begin
      if (_EVAL_37) begin
        _EVAL_53 <= 1'h0;
      end else begin
        _EVAL_53 <= _EVAL_42;
      end
    end
  end
  always @(posedge _EVAL_5 or posedge _EVAL_8) begin
    if (_EVAL_8) begin
      _EVAL_102 <= 1'h0;
    end else if (_EVAL_52) begin
      if (_EVAL_193) begin
        _EVAL_102 <= 1'h0;
      end else begin
        _EVAL_102 <= _EVAL_146;
      end
    end
  end
  always @(posedge _EVAL_5 or posedge _EVAL_8) begin
    if (_EVAL_8) begin
      _EVAL_107 <= 1'h0;
    end else if (_EVAL_150) begin
      if (_EVAL_166) begin
        _EVAL_107 <= 1'h0;
      end else begin
        _EVAL_107 <= _EVAL_133;
      end
    end
  end
  always @(posedge _EVAL_5 or posedge _EVAL_8) begin
    if (_EVAL_8) begin
      _EVAL_188 <= 1'h0;
    end else begin
      _EVAL_188 <= _EVAL_180 & _EVAL_101;
    end
  end
  always @(posedge _EVAL_5 or posedge _EVAL_8) begin
    if (_EVAL_8) begin
      _EVAL_204 <= 1'h0;
    end else if (_EVAL_150) begin
      if (_EVAL_68) begin
        _EVAL_204 <= 1'h0;
      end else begin
        _EVAL_204 <= _EVAL_104;
      end
    end
  end

endmodule
