//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_3_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input  [31:0] _EVAL_4,
  input         _EVAL_5,
  input  [1:0]  _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input  [3:0]  _EVAL_9,
  input  [3:0]  _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [3:0]  _EVAL_17
);
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire [1:0] _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire [5:0] _EVAL_41;
  reg [5:0] _EVAL_42;
  reg [31:0] _RAND_0;
  wire [32:0] _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  reg [1:0] _EVAL_49;
  reg [31:0] _RAND_1;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire [7:0] _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire [32:0] _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  reg [2:0] _EVAL_71;
  reg [31:0] _RAND_2;
  wire  _EVAL_72;
  reg [5:0] _EVAL_73;
  reg [31:0] _RAND_3;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire [31:0] _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire [32:0] _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire [32:0] _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire [6:0] _EVAL_94;
  wire [7:0] _EVAL_95;
  wire  _EVAL_96;
  reg [3:0] _EVAL_97;
  reg [31:0] _RAND_4;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire [6:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire [1:0] _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire [7:0] _EVAL_112;
  wire  _EVAL_113;
  wire [31:0] _EVAL_114;
  wire  _EVAL_115;
  wire [32:0] _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire [3:0] _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire [32:0] _EVAL_126;
  wire [31:0] _EVAL_127;
  wire  _EVAL_128;
  wire [32:0] _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  reg  _EVAL_137;
  reg [31:0] _RAND_5;
  wire [32:0] _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [6:0] _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire [3:0] _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire [32:0] _EVAL_154;
  wire  _EVAL_155;
  wire [32:0] _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire [1:0] _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_162;
  wire [22:0] _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  reg [2:0] _EVAL_171;
  reg [31:0] _RAND_6;
  wire  _EVAL_172;
  wire [32:0] _EVAL_173;
  wire  _EVAL_174;
  wire [5:0] _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire [3:0] _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire [32:0] _EVAL_186;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  reg [31:0] _EVAL_191;
  reg [31:0] _RAND_7;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  reg [31:0] _EVAL_199;
  reg [31:0] _RAND_8;
  wire  _EVAL_200;
  wire [3:0] _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire [32:0] _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  reg  _EVAL_211;
  reg [31:0] _RAND_9;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire [32:0] _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  reg  _EVAL_217;
  reg [31:0] _RAND_10;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire [6:0] _EVAL_220;
  wire  _EVAL_221;
  wire [31:0] _EVAL_222;
  wire [32:0] _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire [5:0] _EVAL_226;
  wire [31:0] _EVAL_227;
  wire  _EVAL_228;
  wire [31:0] _EVAL_229;
  reg [2:0] _EVAL_230;
  reg [31:0] _RAND_11;
  wire  _EVAL_231;
  wire [5:0] _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire [22:0] _EVAL_237;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  reg  _EVAL_249;
  reg [31:0] _RAND_12;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire [5:0] _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire [5:0] _EVAL_269;
  wire [1:0] _EVAL_270;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire [31:0] _EVAL_275;
  wire [32:0] _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire [1:0] _EVAL_280;
  wire  _EVAL_281;
  wire [7:0] _EVAL_283;
  wire  _EVAL_284;
  reg [5:0] _EVAL_285;
  reg [31:0] _RAND_13;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire [32:0] _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  reg [3:0] _EVAL_297;
  reg [31:0] _RAND_14;
  wire [32:0] _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire [32:0] _EVAL_305;
  wire  _EVAL_306;
  wire [31:0] _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  reg [5:0] _EVAL_316;
  reg [31:0] _RAND_15;
  wire  _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_278 = _EVAL_15 & _EVAL_281;
  assign _EVAL_31 = _EVAL_277 ? _EVAL_270 : 2'h0;
  assign _EVAL_129 = _EVAL_186;
  assign _EVAL_29 = _EVAL_10 >= 4'h2;
  assign _EVAL_146 = ~_EVAL_1;
  assign _EVAL_179 = ~_EVAL_13;
  assign _EVAL_173 = _EVAL_85;
  assign _EVAL_138 = {1'b0,$signed(_EVAL_229)};
  assign _EVAL_233 = ~_EVAL_263;
  assign _EVAL_33 = _EVAL_152 & _EVAL_91;
  assign _EVAL_69 = _EVAL_96 | _EVAL_189;
  assign _EVAL_39 = _EVAL_306 | _EVAL_216;
  assign _EVAL_260 = _EVAL & _EVAL_14;
  assign _EVAL_64 = ~_EVAL_87;
  assign _EVAL_18 = _EVAL_114 == 32'h0;
  assign _EVAL_43 = _EVAL_208;
  assign _EVAL_95 = _EVAL_237[7:0];
  assign _EVAL_279 = _EVAL_217 | _EVAL_259;
  assign _EVAL_183 = ~_EVAL_36;
  assign _EVAL_244 = ~_EVAL_122;
  assign _EVAL_89 = _EVAL_179 | _EVAL_3;
  assign _EVAL_84 = _EVAL_7 == 3'h5;
  assign _EVAL_206 = _EVAL_4 == _EVAL_199;
  assign _EVAL_308 = _EVAL_17 == _EVAL_181;
  assign _EVAL_276 = $signed(_EVAL_223) & -33'sh2000;
  assign _EVAL_298 = $signed(_EVAL_214) & -33'sh5000;
  assign _EVAL_292 = ~_EVAL_234;
  assign _EVAL_267 = _EVAL_14 & _EVAL_200;
  assign _EVAL_116 = _EVAL_156;
  assign _EVAL_81 = _EVAL_316 == 6'h0;
  assign _EVAL_151 = _EVAL_197 | _EVAL_8;
  assign _EVAL_140 = ~_EVAL_219;
  assign _EVAL_272 = _EVAL_147 | _EVAL_296;
  assign _EVAL_117 = ~_EVAL_106;
  assign _EVAL_126 = {1'b0,$signed(_EVAL_78)};
  assign _EVAL_273 = _EVAL_248 & _EVAL_74;
  assign _EVAL_124 = _EVAL_302 & _EVAL_53;
  assign _EVAL_170 = _EVAL_14 & _EVAL_210;
  assign _EVAL_190 = ~_EVAL_65;
  assign _EVAL_218 = _EVAL_13 == _EVAL_211;
  assign _EVAL_65 = _EVAL_225 | _EVAL_8;
  assign _EVAL_142 = _EVAL_4[1];
  assign _EVAL_96 = _EVAL_74 | _EVAL_32;
  assign _EVAL_305 = _EVAL_276;
  assign _EVAL_309 = ~_EVAL_182;
  assign _EVAL_51 = _EVAL_111 | _EVAL_8;
  assign _EVAL_74 = $signed(_EVAL_43) == 33'sh0;
  assign _EVAL_36 = _EVAL_83 | _EVAL_8;
  assign _EVAL_236 = _EVAL_272 | _EVAL_33;
  assign _EVAL_155 = _EVAL_145 | _EVAL_8;
  assign _EVAL_112 = ~_EVAL_283;
  assign _EVAL_83 = _EVAL_2 <= 3'h6;
  assign _EVAL_290 = ~_EVAL_121;
  assign _EVAL_270 = 2'h1 << _EVAL_1;
  assign _EVAL_289 = $signed(_EVAL_173) == 33'sh0;
  assign _EVAL_216 = _EVAL_224 & _EVAL_115;
  assign _EVAL_56 = _EVAL_14 & _EVAL_105;
  assign _EVAL_130 = ~_EVAL_187;
  assign _EVAL_109 = ~_EVAL_204;
  assign _EVAL_106 = _EVAL_2 == 3'h6;
  assign _EVAL_115 = $signed(_EVAL_305) == 33'sh0;
  assign _EVAL_21 = ~_EVAL_98;
  assign _EVAL_22 = _EVAL_15 & _EVAL_86;
  assign _EVAL_162 = _EVAL_9[0];
  assign _EVAL_72 = ~_EVAL_128;
  assign _EVAL_258 = _EVAL_12 == _EVAL_230;
  assign _EVAL_28 = _EVAL_120 | _EVAL_8;
  assign _EVAL_182 = _EVAL_29 | _EVAL_8;
  assign _EVAL_104 = _EVAL_141 | _EVAL_203;
  assign _EVAL_255 = _EVAL_279 & _EVAL_110;
  assign _EVAL_234 = _EVAL_7[2];
  assign _EVAL_159 = 2'h1 << _EVAL_162;
  assign _EVAL_98 = _EVAL_146 | _EVAL_8;
  assign _EVAL_103 = _EVAL_73 - 6'h1;
  assign _EVAL_77 = _EVAL_311 | _EVAL_8;
  assign _EVAL_38 = ~_EVAL_51;
  assign _EVAL_61 = _EVAL_205 | _EVAL_8;
  assign _EVAL_123 = ~_EVAL_17;
  assign _EVAL_275 = _EVAL_68[31:0];
  assign _EVAL_187 = _EVAL_19 | _EVAL_8;
  assign _EVAL_62 = _EVAL_218 | _EVAL_8;
  assign _EVAL_256 = _EVAL_288 & _EVAL_302;
  assign _EVAL_79 = ~_EVAL_119;
  assign _EVAL_136 = _EVAL_149 | _EVAL_8;
  assign _EVAL_19 = _EVAL_148 == 4'h0;
  assign _EVAL_283 = _EVAL_164[7:0];
  assign _EVAL_30 = ~_EVAL_151;
  assign _EVAL_160 = _EVAL_241 | _EVAL_8;
  assign _EVAL_143 = _EVAL_285 - 6'h1;
  assign _EVAL_168 = _EVAL_69 | _EVAL_115;
  assign _EVAL_107 = _EVAL_14 & _EVAL_106;
  assign _EVAL_164 = 23'hff << _EVAL_9;
  assign _EVAL_118 = _EVAL_246 | _EVAL_8;
  assign _EVAL_210 = _EVAL_2 == 3'h0;
  assign _EVAL_55 = ~_EVAL_95;
  assign _EVAL_82 = _EVAL_9 <= 4'h6;
  assign _EVAL_87 = _EVAL_157 | _EVAL_8;
  assign _EVAL_319 = ~_EVAL_184;
  assign _EVAL_254 = ~_EVAL_301;
  assign _EVAL_240 = _EVAL_80 & _EVAL_117;
  assign _EVAL_311 = _EVAL_259 | _EVAL_217;
  assign _EVAL_223 = {1'b0,$signed(_EVAL_127)};
  assign _EVAL_312 = ~_EVAL_195;
  assign _EVAL_196 = _EVAL_308 | _EVAL_8;
  assign _EVAL_262 = _EVAL_224 & _EVAL_228;
  assign _EVAL_314 = _EVAL_18 | _EVAL_8;
  assign _EVAL_204 = _EVAL_213 | _EVAL_8;
  assign _EVAL_113 = _EVAL_280[0];
  assign _EVAL_229 = _EVAL_4 ^ 32'h40000000;
  assign _EVAL_193 = _EVAL_15 & _EVAL_185;
  assign _EVAL_299 = _EVAL_152 & _EVAL_192;
  assign _EVAL_205 = _EVAL_12 != 3'h0;
  assign _EVAL_105 = _EVAL_2 == 3'h5;
  assign _EVAL_266 = _EVAL_103[5:0];
  assign _EVAL_78 = _EVAL_4 ^ 32'h2000000;
  assign _EVAL_153 = _EVAL_251 | _EVAL_8;
  assign _EVAL_235 = _EVAL_2[0];
  assign _EVAL_148 = _EVAL_17 & _EVAL_201;
  assign _EVAL_50 = _EVAL_15 & _EVAL_176;
  assign _EVAL_304 = _EVAL_88 | _EVAL_8;
  assign _EVAL_248 = _EVAL_9 <= 4'h8;
  assign _EVAL_253 = _EVAL_152 & _EVAL_124;
  assign _EVAL_133 = _EVAL_7 == _EVAL_71;
  assign _EVAL_188 = ~_EVAL_62;
  assign _EVAL_157 = _EVAL_12 == 3'h0;
  assign _EVAL_184 = _EVAL_265 | _EVAL_8;
  assign _EVAL_288 = _EVAL_108[1];
  assign _EVAL_277 = _EVAL_144 & _EVAL_81;
  assign _EVAL_68 = _EVAL_191 + 32'h1;
  assign _EVAL_135 = _EVAL_152 & _EVAL_131;
  assign _EVAL_195 = _EVAL_76 | _EVAL_8;
  assign _EVAL_192 = _EVAL_302 & _EVAL_231;
  assign _EVAL_175 = _EVAL_143[5:0];
  assign _EVAL_34 = _EVAL_180 | _EVAL_189;
  assign _EVAL_134 = ~_EVAL_28;
  assign _EVAL_166 = _EVAL_42 == 6'h0;
  assign _EVAL_90 = {1'b0,$signed(_EVAL_227)};
  assign _EVAL_201 = ~_EVAL_181;
  assign _EVAL_75 = _EVAL_191 < plusarg_reader_out;
  assign _EVAL_94 = _EVAL_316 - 6'h1;
  assign _EVAL_177 = ~_EVAL_25;
  assign _EVAL_295 = _EVAL_70 | _EVAL_8;
  assign _EVAL_176 = _EVAL_7 == 3'h3;
  assign _EVAL_317 = _EVAL_147 | _EVAL_256;
  assign _EVAL_144 = _EVAL_16 & _EVAL_15;
  assign _EVAL_228 = _EVAL_34 | _EVAL_115;
  assign _EVAL_198 = _EVAL_7 == 3'h6;
  assign _EVAL_286 = ~_EVAL_47;
  assign _EVAL_46 = _EVAL_14 & _EVAL_284;
  assign _EVAL_200 = _EVAL_2 == 3'h2;
  assign _EVAL_32 = $signed(_EVAL_116) == 33'sh0;
  assign _EVAL_52 = ~_EVAL_318;
  assign _EVAL_91 = _EVAL_142 & _EVAL_231;
  assign _EVAL_44 = _EVAL_207 | _EVAL_8;
  assign _EVAL_232 = _EVAL_94[5:0];
  assign _EVAL_214 = {1'b0,$signed(_EVAL_4)};
  assign _EVAL_25 = _EVAL_179 | _EVAL_8;
  assign _EVAL_145 = _EVAL_104 | _EVAL_75;
  assign _EVAL_167 = ~_EVAL_77;
  assign _EVAL_88 = _EVAL_6 == 2'h0;
  assign _EVAL_149 = _EVAL_12 <= 3'h4;
  assign _EVAL_131 = _EVAL_142 & _EVAL_53;
  assign _EVAL_180 = _EVAL_264 | _EVAL_32;
  assign _EVAL_203 = plusarg_reader_out == 32'h0;
  assign _EVAL_224 = _EVAL_9 <= 4'h2;
  assign _EVAL_80 = _EVAL_260 & _EVAL_26;
  assign _EVAL_139 = _EVAL_260 & _EVAL_166;
  assign _EVAL_99 = _EVAL_259 != _EVAL_113;
  assign _EVAL_66 = ~_EVAL_118;
  assign _EVAL_222 = {{24'd0}, _EVAL_112};
  assign _EVAL_263 = _EVAL_147 | _EVAL_8;
  assign _EVAL_287 = _EVAL_245 | _EVAL_273;
  assign _EVAL_247 = _EVAL_252 | _EVAL_8;
  assign _EVAL_318 = _EVAL_89 | _EVAL_8;
  assign _EVAL_252 = _EVAL_12 <= 3'h1;
  assign _EVAL_197 = _EVAL_1 == _EVAL_137;
  assign _EVAL_293 = {1'b0,$signed(_EVAL_307)};
  assign _EVAL_231 = _EVAL_4[0];
  assign _EVAL_53 = ~_EVAL_231;
  assign _EVAL_280 = _EVAL_240 ? 2'h1 : 2'h0;
  assign _EVAL_132 = ~_EVAL_48;
  assign _EVAL_284 = ~_EVAL_166;
  assign _EVAL_122 = _EVAL_303 | _EVAL_8;
  assign _EVAL_45 = ~_EVAL_44;
  assign _EVAL_296 = _EVAL_288 & _EVAL_142;
  assign _EVAL_237 = 23'hff << _EVAL_10;
  assign _EVAL_307 = _EVAL_4 ^ 32'h80000000;
  assign _EVAL_57 = _EVAL_15 & _EVAL_286;
  assign _EVAL_215 = _EVAL_7 == 3'h7;
  assign _EVAL_208 = $signed(_EVAL_90) & -33'sh1000;
  assign _EVAL_111 = _EVAL_12 <= 3'h2;
  assign _EVAL_306 = _EVAL_100 | _EVAL_273;
  assign _EVAL_141 = ~_EVAL_217;
  assign _EVAL_154 = _EVAL_298;
  assign _EVAL_54 = _EVAL_15 & _EVAL_84;
  assign _EVAL_264 = $signed(_EVAL_129) == 33'sh0;
  assign _EVAL_158 = ~_EVAL_136;
  assign _EVAL_257 = ~_EVAL_5;
  assign _EVAL_27 = _EVAL_6 == _EVAL_49;
  assign _EVAL_120 = _EVAL_9 == _EVAL_297;
  assign _EVAL_181 = {_EVAL_236,_EVAL_221,_EVAL_172,_EVAL_212};
  assign _EVAL_259 = _EVAL_31[0];
  assign _EVAL_265 = _EVAL_11 == _EVAL_249;
  assign _EVAL_147 = _EVAL_9 >= 4'h2;
  assign _EVAL_85 = $signed(_EVAL_138) & -33'sh2000;
  assign _EVAL_300 = _EVAL_144 & _EVAL_47;
  assign _EVAL_207 = _EVAL_2 == _EVAL_171;
  assign _EVAL_186 = $signed(_EVAL_293) & -33'shc000;
  assign _EVAL_226 = _EVAL_55[7:2];
  assign _EVAL_268 = ~_EVAL_295;
  assign _EVAL_313 = _EVAL_14 & _EVAL_202;
  assign _EVAL_241 = _EVAL_6 != 2'h2;
  assign _EVAL_76 = _EVAL_165 | _EVAL_273;
  assign _EVAL_37 = ~_EVAL_314;
  assign _EVAL_165 = _EVAL_224 & _EVAL_34;
  assign _EVAL_63 = _EVAL_217 >> _EVAL_1;
  assign _EVAL_119 = _EVAL_206 | _EVAL_8;
  assign _EVAL_108 = _EVAL_159 | 2'h1;
  assign _EVAL_221 = _EVAL_272 | _EVAL_135;
  assign _EVAL_127 = _EVAL_4 ^ 32'h20000000;
  assign _EVAL_213 = ~_EVAL_3;
  assign _EVAL_315 = ~_EVAL_196;
  assign _EVAL_178 = ~_EVAL_261;
  assign _EVAL_48 = _EVAL_27 | _EVAL_8;
  assign _EVAL_58 = _EVAL_123 == 4'h0;
  assign _EVAL_219 = _EVAL_194 | _EVAL_8;
  assign _EVAL_60 = ~_EVAL_174;
  assign _EVAL_110 = ~_EVAL_113;
  assign _EVAL_172 = _EVAL_317 | _EVAL_299;
  assign _EVAL_24 = ~_EVAL_259;
  assign _EVAL_100 = _EVAL_82 & _EVAL_289;
  assign _EVAL_114 = _EVAL_4 & _EVAL_222;
  assign _EVAL_245 = _EVAL_262 | _EVAL_100;
  assign _EVAL_261 = _EVAL_133 | _EVAL_8;
  assign _EVAL_121 = _EVAL_258 | _EVAL_8;
  assign _EVAL_291 = _EVAL_144 | _EVAL_260;
  assign _EVAL_128 = _EVAL_39 | _EVAL_8;
  assign _EVAL_227 = _EVAL_4 ^ 32'h3000;
  assign _EVAL_251 = _EVAL_10 == _EVAL_97;
  assign _EVAL_194 = _EVAL_12 <= 3'h3;
  assign _EVAL_250 = ~_EVAL_61;
  assign _EVAL_41 = _EVAL_220[5:0];
  assign _EVAL_150 = _EVAL_7 == 3'h4;
  assign _EVAL_93 = _EVAL_287 | _EVAL_8;
  assign _EVAL_301 = _EVAL_58 | _EVAL_8;
  assign _EVAL_269 = _EVAL_112[7:2];
  assign _EVAL_67 = ~_EVAL_155;
  assign _EVAL_125 = _EVAL_14 & _EVAL_294;
  assign _EVAL_246 = _EVAL_99 | _EVAL_24;
  assign _EVAL_101 = ~_EVAL_160;
  assign _EVAL_220 = _EVAL_42 - 6'h1;
  assign _EVAL_152 = _EVAL_108[0];
  assign _EVAL_92 = ~_EVAL_93;
  assign _EVAL_281 = _EVAL_7 == 3'h0;
  assign _EVAL_310 = _EVAL_15 & _EVAL_215;
  assign _EVAL_294 = _EVAL_2 == 3'h1;
  assign _EVAL_209 = ~_EVAL_8;
  assign _EVAL_59 = ~_EVAL_153;
  assign _EVAL_212 = _EVAL_317 | _EVAL_253;
  assign _EVAL_274 = _EVAL_15 & _EVAL_198;
  assign _EVAL_202 = _EVAL_2 == 3'h4;
  assign _EVAL_189 = $signed(_EVAL_154) == 33'sh0;
  assign _EVAL_174 = _EVAL_257 | _EVAL_8;
  assign _EVAL_23 = ~_EVAL_247;
  assign _EVAL_185 = _EVAL_7 == 3'h1;
  assign _EVAL_302 = ~_EVAL_142;
  assign _EVAL_225 = _EVAL_6 <= 2'h2;
  assign _EVAL_70 = _EVAL_224 & _EVAL_168;
  assign _EVAL_169 = _EVAL_15 & _EVAL_150;
  assign _EVAL_20 = ~_EVAL_304;
  assign _EVAL_303 = ~_EVAL_63;
  assign _EVAL_156 = $signed(_EVAL_126) & -33'sh1000000;
  assign _EVAL_47 = _EVAL_285 == 6'h0;
  assign _EVAL_26 = _EVAL_73 == 6'h0;
  assign _EVAL_86 = _EVAL_7 == 3'h2;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_42 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_49 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_71 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_73 = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_97 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_137 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_171 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_191 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_199 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_211 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_217 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_230 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_249 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_285 = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_297 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_316 = _RAND_15[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_0) begin
    if (_EVAL_8) begin
      _EVAL_42 <= 6'h0;
    end else if (_EVAL_260) begin
      if (_EVAL_166) begin
        if (_EVAL_235) begin
          _EVAL_42 <= _EVAL_226;
        end else begin
          _EVAL_42 <= 6'h0;
        end
      end else begin
        _EVAL_42 <= _EVAL_41;
      end
    end
    if (_EVAL_139) begin
      _EVAL_49 <= _EVAL_6;
    end
    if (_EVAL_300) begin
      _EVAL_71 <= _EVAL_7;
    end
    if (_EVAL_8) begin
      _EVAL_73 <= 6'h0;
    end else if (_EVAL_260) begin
      if (_EVAL_26) begin
        if (_EVAL_235) begin
          _EVAL_73 <= _EVAL_226;
        end else begin
          _EVAL_73 <= 6'h0;
        end
      end else begin
        _EVAL_73 <= _EVAL_266;
      end
    end
    if (_EVAL_139) begin
      _EVAL_97 <= _EVAL_10;
    end
    if (_EVAL_300) begin
      _EVAL_137 <= _EVAL_1;
    end
    if (_EVAL_139) begin
      _EVAL_171 <= _EVAL_2;
    end
    if (_EVAL_8) begin
      _EVAL_191 <= 32'h0;
    end else if (_EVAL_291) begin
      _EVAL_191 <= 32'h0;
    end else begin
      _EVAL_191 <= _EVAL_275;
    end
    if (_EVAL_300) begin
      _EVAL_199 <= _EVAL_4;
    end
    if (_EVAL_139) begin
      _EVAL_211 <= _EVAL_13;
    end
    if (_EVAL_8) begin
      _EVAL_217 <= 1'h0;
    end else begin
      _EVAL_217 <= _EVAL_255;
    end
    if (_EVAL_300) begin
      _EVAL_230 <= _EVAL_12;
    end
    if (_EVAL_139) begin
      _EVAL_249 <= _EVAL_11;
    end
    if (_EVAL_8) begin
      _EVAL_285 <= 6'h0;
    end else if (_EVAL_144) begin
      if (_EVAL_47) begin
        if (_EVAL_292) begin
          _EVAL_285 <= _EVAL_269;
        end else begin
          _EVAL_285 <= 6'h0;
        end
      end else begin
        _EVAL_285 <= _EVAL_175;
      end
    end
    if (_EVAL_300) begin
      _EVAL_297 <= _EVAL_9;
    end
    if (_EVAL_8) begin
      _EVAL_316 <= 6'h0;
    end else if (_EVAL_144) begin
      if (_EVAL_81) begin
        if (_EVAL_292) begin
          _EVAL_316 <= _EVAL_269;
        end else begin
          _EVAL_316 <= 6'h0;
        end
      end else begin
        _EVAL_316 <= _EVAL_232;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(973d3d27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b7e2cac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cc9430e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_315) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75a7bb37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfc1e5e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_319) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3077870c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87c34980)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7948daa4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4e3b221)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c094666d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_315) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62e42b01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b5539e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45020510)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3eaf366)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb676072)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f03cefcd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_315) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e18949fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c4d8f9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9501695)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9160c6cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c11b9cdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(159644f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45ef046c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7703fe8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(404f295b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(126f11b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe1a54e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3b3550b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57675fe7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acc4a14e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_315) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28e080c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95bcd848)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2374d12d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1eccbe17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f235c2f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bcf3968)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4f4f5b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba03a61b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e667d8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ecb7afa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(896fab16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d7a156)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c30990e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f14de05b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6de631c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(375bbfd9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a41a0eeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(100314c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b0bd75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78f12382)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27ab42c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34c54d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb149846)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8d1200a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecde388b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(497409d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_319) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3303b7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf0d49c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3de62cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14a1d723)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5823fdee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7f13ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_315) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_315) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87dd874c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d7d8eed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dba0e9fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_315) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6998087)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b367ae7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_315) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed999f5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(255330cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d10e8b63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d9c690a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3333342)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b648c4b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f868aba1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5f7fbff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b8b7769)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a9556a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3eaeb681)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c001ef10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_315) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32c875c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(201427d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_315) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13fa6ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd25b46c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb5087ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
