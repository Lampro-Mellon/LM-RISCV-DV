//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
bind _EVAL_4 _EVAL_4_assert _EVAL_4_assert_0 (.*);
bind _EVAL_6 _EVAL_6_assert _EVAL_6_assert_0 (.*);
bind _EVAL_8 _EVAL_8_assert _EVAL_8_assert_0 (.*);
bind _EVAL_11 _EVAL_11_assert _EVAL_11_assert_0 (.*);
bind _EVAL_13 _EVAL_13_assert _EVAL_13_assert_0 (.*);
bind _EVAL_16 _EVAL_16_assert _EVAL_16_assert_0 (.*);
bind _EVAL_18 _EVAL_18_assert _EVAL_18_assert_0 (.*);
bind _EVAL_22 _EVAL_22_assert _EVAL_22_assert_0 (.*);
bind _EVAL_24 _EVAL_24_assert _EVAL_24_assert_0 (.*);
bind _EVAL_26 _EVAL_26_assert _EVAL_26_assert_0 (.*);
bind _EVAL_28 _EVAL_28_assert _EVAL_28_assert_0 (.*);
bind _EVAL_32 _EVAL_32_assert _EVAL_32_assert_0 (.*);
bind _EVAL_35 _EVAL_35_assert _EVAL_35_assert_0 (.*);
bind _EVAL_41 _EVAL_41_assert _EVAL_41_assert_0 (.*);
bind _EVAL_45 _EVAL_45_assert _EVAL_45_assert_0 (.*);
bind _EVAL_47 _EVAL_47_assert _EVAL_47_assert_0 (.*);
bind _EVAL_49 _EVAL_49_assert _EVAL_49_assert_0 (.*);
bind _EVAL_50 _EVAL_50_assert _EVAL_50_assert_0 (.*);
bind _EVAL_54 _EVAL_54_assert _EVAL_54_assert_0 (.*);
bind _EVAL_59 _EVAL_59_assert _EVAL_59_assert_0 (.*);
bind _EVAL_61 _EVAL_61_assert _EVAL_61_assert_0 (.*);
bind _EVAL_63 _EVAL_63_assert _EVAL_63_assert_0 (.*);
bind _EVAL_67 _EVAL_67_assert _EVAL_67_assert_0 (.*);
bind _EVAL_69 _EVAL_69_assert _EVAL_69_assert_0 (.*);
bind _EVAL_72 _EVAL_72_assert _EVAL_72_assert_0 (.*);
bind _EVAL_75 _EVAL_75_assert _EVAL_75_assert_0 (.*);
bind _EVAL_78 _EVAL_78_assert _EVAL_78_assert_0 (.*);
bind _EVAL_81 _EVAL_81_assert _EVAL_81_assert_0 (.*);
bind _EVAL_85 _EVAL_85_assert _EVAL_85_assert_0 (.*);
bind _EVAL_89 _EVAL_89_assert _EVAL_89_assert_0 (.*);
bind _EVAL_91 _EVAL_91_assert _EVAL_91_assert_0 (.*);
bind _EVAL_93 _EVAL_93_assert _EVAL_93_assert_0 (.*);
bind _EVAL_95 _EVAL_95_assert _EVAL_95_assert_0 (.*);
bind _EVAL_99 _EVAL_99_assert _EVAL_99_assert_0 (.*);
bind _EVAL_101 _EVAL_101_assert _EVAL_101_assert_0 (.*);
bind _EVAL_106 _EVAL_106_assert _EVAL_106_assert_0 (.*);
bind _EVAL_116 _EVAL_116_assert _EVAL_116_assert_0 (.*);
bind _EVAL_118 _EVAL_118_assert _EVAL_118_assert_0 (.*);
bind _EVAL_121 _EVAL_121_assert _EVAL_121_assert_0 (.*);
bind _EVAL_124 _EVAL_124_assert _EVAL_124_assert_0 (.*);
bind _EVAL_126 _EVAL_126_assert _EVAL_126_assert_0 (.*);
bind _EVAL_134 _EVAL_134_assert _EVAL_134_assert_0 (.*);
bind _EVAL_141 _EVAL_141_assert _EVAL_141_assert_0 (.*);
bind _EVAL_145 _EVAL_145_assert _EVAL_145_assert_0 (.*);
bind _EVAL_151 _EVAL_151_assert _EVAL_151_assert_0 (.*);
bind _EVAL_154 _EVAL_154_assert _EVAL_154_assert_0 (.*);
bind _EVAL_156 _EVAL_156_assert _EVAL_156_assert_0 (.*);
bind _EVAL_158 _EVAL_158_assert _EVAL_158_assert_0 (.*);
bind _EVAL_160 _EVAL_160_assert _EVAL_160_assert_0 (.*);
bind _EVAL_162 _EVAL_162_assert _EVAL_162_assert_0 (.*);
bind _EVAL_164 _EVAL_164_assert _EVAL_164_assert_0 (.*);
bind _EVAL_165 _EVAL_165_assert _EVAL_165_assert_0 (.*);
bind _EVAL_167 _EVAL_167_assert _EVAL_167_assert_0 (.*);
bind _EVAL_169 _EVAL_169_assert _EVAL_169_assert_0 (.*);
bind _EVAL_172 _EVAL_172_assert _EVAL_172_assert_0 (.*);
bind _EVAL_174 _EVAL_174_assert _EVAL_174_assert_0 (.*);
bind _EVAL_177 _EVAL_177_assert _EVAL_177_assert_0 (.*);
bind SiFive_TLTestIndicator SiFive_TLTestIndicator_assert SiFive_TLTestIndicator_assert_0 (.*);
bind _EVAL_180 _EVAL_180_assert _EVAL_180_assert_0 (.*);
bind _EVAL_181 _EVAL_181_assert _EVAL_181_assert_0 (.*);
bind _EVAL_182 _EVAL_182_assert _EVAL_182_assert_0 (.*);
bind _EVAL_183 _EVAL_183_assert _EVAL_183_assert_0 (.*);
bind _EVAL_184 _EVAL_184_assert _EVAL_184_assert_0 (.*);
bind _EVAL_186 _EVAL_186_assert _EVAL_186_assert_0 (.*);
bind _EVAL_187 _EVAL_187_assert _EVAL_187_assert_0 (.*);