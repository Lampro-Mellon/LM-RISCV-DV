//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_12_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input  [1:0]  _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  input  [3:0]  _EVAL_6,
  input         _EVAL_7,
  input  [31:0] _EVAL_8,
  input         _EVAL_9,
  input  [1:0]  _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [2:0]  _EVAL_13,
  input         _EVAL_14
);
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  reg [2:0] _EVAL_19;
  reg [31:0] _RAND_0;
  wire  _EVAL_20;
  wire [1:0] _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  reg [2:0] _EVAL_24;
  reg [31:0] _RAND_1;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire [32:0] _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire [4:0] _EVAL_33;
  wire  _EVAL_34;
  wire [1:0] _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire [7:0] _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire [7:0] _EVAL_48;
  wire  _EVAL_49;
  reg [1:0] _EVAL_50;
  reg [31:0] _RAND_2;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire [1:0] _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire [4:0] _EVAL_62;
  wire [4:0] _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  reg [2:0] _EVAL_80;
  reg [31:0] _RAND_3;
  wire  _EVAL_81;
  reg  _EVAL_82;
  reg [31:0] _RAND_4;
  wire [32:0] _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire [1:0] _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire [1:0] _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_113;
  wire [31:0] plusarg_reader_out;
  reg [1:0] _EVAL_114;
  reg [31:0] _RAND_5;
  wire [4:0] _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire [3:0] _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire [4:0] _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire [3:0] _EVAL_126;
  wire  _EVAL_127;
  wire [4:0] _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire [31:0] _EVAL_135;
  wire  _EVAL_136;
  reg  _EVAL_137;
  reg [31:0] _RAND_6;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire [4:0] _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  reg [2:0] _EVAL_149;
  reg [31:0] _RAND_7;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire [3:0] _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  reg [4:0] _EVAL_155;
  reg [31:0] _RAND_8;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire [1:0] _EVAL_160;
  wire [32:0] _EVAL_162;
  wire [1:0] _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire [31:0] _EVAL_166;
  wire [1:0] _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  reg [31:0] _EVAL_173;
  reg [31:0] _RAND_9;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire [3:0] _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire [1:0] _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire [4:0] _EVAL_200;
  reg [2:0] _EVAL_201;
  reg [31:0] _RAND_10;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  reg  _EVAL_215;
  reg [31:0] _RAND_11;
  wire [7:0] _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire [4:0] _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire [31:0] _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire [1:0] _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  reg  _EVAL_238;
  reg [31:0] _RAND_12;
  wire  _EVAL_239;
  wire [7:0] _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire [31:0] _EVAL_244;
  reg [31:0] _EVAL_245;
  reg [31:0] _RAND_13;
  wire [32:0] _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_31 = _EVAL_9 & _EVAL_38;
  assign _EVAL_196 = ~_EVAL_146;
  assign _EVAL_110 = ~_EVAL_158;
  assign _EVAL_158 = _EVAL_208 | _EVAL;
  assign _EVAL_96 = _EVAL_119 == 4'h0;
  assign _EVAL_169 = _EVAL_47 & _EVAL_214;
  assign _EVAL_234 = ~_EVAL_214;
  assign _EVAL_81 = _EVAL_232 | _EVAL;
  assign _EVAL_194 = _EVAL_4 == _EVAL_19;
  assign _EVAL_108 = ~_EVAL_183;
  assign _EVAL_93 = _EVAL_8 == _EVAL_245;
  assign _EVAL_243 = _EVAL_12 <= 3'h1;
  assign _EVAL_116 = ~_EVAL;
  assign _EVAL_144 = _EVAL_25 | _EVAL;
  assign _EVAL_205 = _EVAL_7 & _EVAL_177;
  assign _EVAL_35 = _EVAL_33[1:0];
  assign _EVAL_242 = _EVAL_4 <= 3'h6;
  assign _EVAL_247 = _EVAL_168 == 2'h0;
  assign _EVAL_191 = _EVAL_7 & _EVAL_140;
  assign _EVAL_125 = _EVAL_7 & _EVAL_94;
  assign _EVAL_246 = {1'b0,$signed(_EVAL_228)};
  assign _EVAL_54 = ~_EVAL_120;
  assign _EVAL_59 = _EVAL_0[2:1];
  assign _EVAL_126 = _EVAL_6 & _EVAL_179;
  assign _EVAL_228 = _EVAL_8 ^ 32'h80000000;
  assign _EVAL_244 = _EVAL_8 & _EVAL_135;
  assign _EVAL_75 = _EVAL_26 | _EVAL_207;
  assign _EVAL_189 = _EVAL_197 | _EVAL_133;
  assign _EVAL_166 = _EVAL_83[31:0];
  assign _EVAL_28 = _EVAL_10 == _EVAL_114;
  assign _EVAL_179 = ~_EVAL_152;
  assign _EVAL_97 = _EVAL_235 | _EVAL;
  assign _EVAL_208 = _EVAL_111 | _EVAL_250;
  assign _EVAL_199 = ~_EVAL_225;
  assign _EVAL_227 = _EVAL_212 & _EVAL_43;
  assign _EVAL_121 = ~_EVAL_79;
  assign _EVAL_207 = _EVAL_173 < plusarg_reader_out;
  assign _EVAL_63 = _EVAL_123 >> _EVAL_5;
  assign _EVAL_79 = _EVAL_53 | _EVAL;
  assign _EVAL_43 = ~_EVAL_82;
  assign _EVAL_68 = _EVAL_109 | _EVAL_154;
  assign _EVAL_102 = _EVAL_59 == 2'h1;
  assign _EVAL_240 = _EVAL_69 ? _EVAL_39 : 8'h0;
  assign _EVAL_233 = ~_EVAL_238;
  assign _EVAL_130 = _EVAL_155 | _EVAL_220;
  assign _EVAL_159 = ~_EVAL_32;
  assign _EVAL_176 = _EVAL_16 | _EVAL;
  assign _EVAL_213 = ~_EVAL_215;
  assign _EVAL_115 = _EVAL_130 & _EVAL_62;
  assign _EVAL_188 = _EVAL_101 | 2'h1;
  assign _EVAL_232 = _EVAL_2 == _EVAL_50;
  assign _EVAL_51 = ~_EVAL_176;
  assign _EVAL_142 = _EVAL_96 | _EVAL;
  assign _EVAL_181 = _EVAL_9 & _EVAL_41;
  assign _EVAL_32 = _EVAL_103 | _EVAL;
  assign _EVAL_170 = ~_EVAL_157;
  assign _EVAL_39 = 8'h1 << _EVAL_5;
  assign _EVAL_49 = _EVAL_65 | _EVAL;
  assign _EVAL_235 = _EVAL_5 == _EVAL_201;
  assign _EVAL_225 = _EVAL_93 | _EVAL;
  assign _EVAL_251 = _EVAL_231[0];
  assign _EVAL_64 = _EVAL_105[0];
  assign _EVAL_77 = $signed(_EVAL_162) == 33'sh0;
  assign _EVAL_83 = _EVAL_173 + 32'h1;
  assign _EVAL_84 = _EVAL_188[1];
  assign _EVAL_29 = $signed(_EVAL_246) & -33'sh4000;
  assign _EVAL_134 = ~_EVAL_202;
  assign _EVAL_60 = _EVAL_212 & _EVAL_213;
  assign _EVAL_132 = _EVAL_7 & _EVAL_156;
  assign _EVAL_221 = _EVAL_61 & _EVAL_234;
  assign _EVAL_124 = _EVAL_13 == 3'h3;
  assign _EVAL_193 = _EVAL_7 & _EVAL_73;
  assign _EVAL_214 = _EVAL_8[0];
  assign _EVAL_217 = _EVAL_6 == _EVAL_152;
  assign _EVAL_30 = plusarg_reader_out == 32'h0;
  assign _EVAL_15 = _EVAL_63[0];
  assign _EVAL_90 = _EVAL_46 | _EVAL_98;
  assign _EVAL_27 = _EVAL_9 & _EVAL_183;
  assign _EVAL_183 = _EVAL_4 == 3'h6;
  assign _EVAL_198 = ~_EVAL_1;
  assign _EVAL_241 = ~_EVAL_81;
  assign _EVAL_26 = _EVAL_138 | _EVAL_30;
  assign _EVAL_101 = 2'h1 << _EVAL_104;
  assign _EVAL_136 = _EVAL_242 | _EVAL;
  assign _EVAL_122 = _EVAL_4 == 3'h1;
  assign _EVAL_41 = _EVAL_4 == 3'h5;
  assign _EVAL_203 = _EVAL_184 | _EVAL_107;
  assign _EVAL_151 = _EVAL_212 | _EVAL_44;
  assign _EVAL_76 = ~_EVAL_22;
  assign _EVAL_160 = _EVAL_238 - 1'h1;
  assign _EVAL_58 = _EVAL_175 | _EVAL;
  assign _EVAL_248 = _EVAL_84 & _EVAL_61;
  assign _EVAL_120 = _EVAL_127 | _EVAL;
  assign _EVAL_70 = _EVAL_13 == _EVAL_80;
  assign _EVAL_141 = _EVAL_240[4:0];
  assign _EVAL_168 = _EVAL_5[2:1];
  assign _EVAL_103 = _EVAL_12 <= 3'h2;
  assign _EVAL_220 = _EVAL_48[4:0];
  assign _EVAL_74 = _EVAL_165 | _EVAL;
  assign _EVAL_55 = _EVAL_218 & _EVAL_222;
  assign _EVAL_223 = _EVAL_12 == 3'h0;
  assign _EVAL_92 = _EVAL_4 == 3'h2;
  assign _EVAL_162 = _EVAL_29;
  assign _EVAL_38 = ~_EVAL_233;
  assign _EVAL_61 = _EVAL_8[1];
  assign _EVAL_52 = _EVAL_189 | _EVAL;
  assign _EVAL_71 = _EVAL_84 & _EVAL_47;
  assign _EVAL_150 = _EVAL_44 & _EVAL_233;
  assign _EVAL_69 = _EVAL_249 & _EVAL_108;
  assign _EVAL_104 = _EVAL_10[0];
  assign _EVAL_73 = _EVAL_13 == 3'h6;
  assign _EVAL_18 = ~_EVAL_43;
  assign _EVAL_36 = _EVAL_61 & _EVAL_214;
  assign _EVAL_218 = _EVAL_188[0];
  assign _EVAL_119 = ~_EVAL_6;
  assign _EVAL_135 = {{30'd0}, _EVAL_21};
  assign _EVAL_236 = ~_EVAL_178;
  assign _EVAL_226 = _EVAL_160[0];
  assign _EVAL_195 = ~_EVAL_136;
  assign _EVAL_143 = ~_EVAL_85;
  assign _EVAL_45 = _EVAL_217 | _EVAL;
  assign _EVAL_131 = ~_EVAL_52;
  assign _EVAL_46 = _EVAL_40 | _EVAL_71;
  assign _EVAL_113 = _EVAL_9 & _EVAL_122;
  assign _EVAL_48 = _EVAL_60 ? _EVAL_216 : 8'h0;
  assign _EVAL_56 = _EVAL_46 | _EVAL_55;
  assign _EVAL_40 = _EVAL_10 >= 2'h2;
  assign _EVAL_172 = ~_EVAL_237;
  assign _EVAL_86 = _EVAL_200[0];
  assign _EVAL_200 = _EVAL_155 >> _EVAL_0;
  assign _EVAL_180 = _EVAL_203 | _EVAL;
  assign _EVAL_16 = _EVAL_12 != 3'h0;
  assign _EVAL_216 = 8'h1 << _EVAL_0;
  assign _EVAL_85 = _EVAL_40 | _EVAL;
  assign _EVAL_202 = _EVAL_243 | _EVAL;
  assign _EVAL_171 = _EVAL_244 == 32'h0;
  assign _EVAL_192 = _EVAL_4 == 3'h4;
  assign _EVAL_204 = _EVAL_198 | _EVAL;
  assign _EVAL_57 = ~_EVAL_137;
  assign _EVAL_209 = _EVAL_9 & _EVAL_23;
  assign _EVAL_88 = _EVAL_9 & _EVAL_192;
  assign _EVAL_25 = _EVAL_2 >= 2'h2;
  assign _EVAL_178 = _EVAL_75 | _EVAL;
  assign _EVAL_72 = _EVAL_28 | _EVAL;
  assign _EVAL_190 = _EVAL_10 <= 2'h2;
  assign _EVAL_164 = _EVAL_9 & _EVAL_92;
  assign _EVAL_123 = _EVAL_220 | _EVAL_155;
  assign _EVAL_230 = _EVAL_12 == _EVAL_149;
  assign _EVAL_37 = _EVAL_7 & _EVAL_124;
  assign _EVAL_157 = _EVAL_171 | _EVAL;
  assign _EVAL_148 = ~_EVAL_72;
  assign _EVAL_185 = ~_EVAL_180;
  assign _EVAL_186 = ~_EVAL_144;
  assign _EVAL_153 = _EVAL_7 & _EVAL_224;
  assign _EVAL_250 = _EVAL_0 == 3'h4;
  assign _EVAL_21 = ~_EVAL_35;
  assign _EVAL_34 = _EVAL_59 == 2'h0;
  assign _EVAL_239 = ~_EVAL_204;
  assign _EVAL_105 = _EVAL_215 - 1'h1;
  assign _EVAL_117 = _EVAL_15 | _EVAL;
  assign _EVAL_211 = _EVAL_126 == 4'h0;
  assign _EVAL_152 = {_EVAL_68,_EVAL_89,_EVAL_90,_EVAL_56};
  assign _EVAL_229 = ~_EVAL_142;
  assign _EVAL_184 = _EVAL_220 != _EVAL_141;
  assign _EVAL_62 = ~_EVAL_141;
  assign _EVAL_182 = _EVAL_211 | _EVAL;
  assign _EVAL_22 = _EVAL_230 | _EVAL;
  assign _EVAL_133 = _EVAL_5 == 3'h4;
  assign _EVAL_65 = _EVAL_12 <= 3'h3;
  assign _EVAL_89 = _EVAL_109 | _EVAL_174;
  assign _EVAL_163 = _EVAL_137 - 1'h1;
  assign _EVAL_156 = _EVAL_13 == 3'h5;
  assign _EVAL_100 = ~_EVAL_45;
  assign _EVAL_231 = _EVAL_82 - 1'h1;
  assign _EVAL_78 = _EVAL_163[0];
  assign _EVAL_197 = _EVAL_99 | _EVAL_247;
  assign _EVAL_165 = _EVAL_190 & _EVAL_77;
  assign _EVAL_87 = ~_EVAL_97;
  assign _EVAL_44 = _EVAL_14 & _EVAL_9;
  assign _EVAL_127 = ~_EVAL_86;
  assign _EVAL_53 = _EVAL_12 <= 3'h4;
  assign _EVAL_147 = ~_EVAL_118;
  assign _EVAL_154 = _EVAL_218 & _EVAL_36;
  assign _EVAL_33 = 5'h3 << _EVAL_10;
  assign _EVAL_219 = ~_EVAL_49;
  assign _EVAL_175 = _EVAL_0 == _EVAL_24;
  assign _EVAL_140 = _EVAL_13 == 3'h0;
  assign _EVAL_91 = ~_EVAL_117;
  assign _EVAL_107 = ~_EVAL_206;
  assign _EVAL_138 = ~_EVAL_42;
  assign _EVAL_47 = ~_EVAL_61;
  assign _EVAL_20 = ~_EVAL_74;
  assign _EVAL_224 = _EVAL_13 == 3'h7;
  assign _EVAL_17 = _EVAL_13 == 3'h2;
  assign _EVAL_94 = _EVAL_13 == 3'h1;
  assign _EVAL_212 = _EVAL_11 & _EVAL_7;
  assign _EVAL_95 = ~_EVAL_182;
  assign _EVAL_222 = _EVAL_47 & _EVAL_234;
  assign _EVAL_106 = _EVAL_7 & _EVAL_18;
  assign _EVAL_98 = _EVAL_218 & _EVAL_169;
  assign _EVAL_206 = _EVAL_220 != 5'h0;
  assign _EVAL_139 = ~_EVAL_58;
  assign _EVAL_249 = _EVAL_44 & _EVAL_57;
  assign _EVAL_66 = _EVAL_7 & _EVAL_17;
  assign _EVAL_146 = _EVAL_223 | _EVAL;
  assign _EVAL_237 = _EVAL_194 | _EVAL;
  assign _EVAL_174 = _EVAL_218 & _EVAL_221;
  assign _EVAL_118 = _EVAL_70 | _EVAL;
  assign _EVAL_109 = _EVAL_40 | _EVAL_248;
  assign _EVAL_23 = _EVAL_4 == 3'h0;
  assign _EVAL_111 = _EVAL_102 | _EVAL_34;
  assign _EVAL_99 = _EVAL_168 == 2'h1;
  assign _EVAL_177 = _EVAL_13 == 3'h4;
  assign _EVAL_42 = _EVAL_155 != 5'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_19 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_24 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_50 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_80 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_82 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_114 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_137 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_149 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_155 = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_173 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_201 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_215 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_238 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_245 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_3) begin
    if (_EVAL_150) begin
      _EVAL_19 <= _EVAL_4;
    end
    if (_EVAL_227) begin
      _EVAL_24 <= _EVAL_0;
    end
    if (_EVAL_150) begin
      _EVAL_50 <= _EVAL_2;
    end
    if (_EVAL_227) begin
      _EVAL_80 <= _EVAL_13;
    end
    if (_EVAL) begin
      _EVAL_82 <= 1'h0;
    end else if (_EVAL_212) begin
      if (_EVAL_43) begin
        _EVAL_82 <= 1'h0;
      end else begin
        _EVAL_82 <= _EVAL_251;
      end
    end
    if (_EVAL_227) begin
      _EVAL_114 <= _EVAL_10;
    end
    if (_EVAL) begin
      _EVAL_137 <= 1'h0;
    end else if (_EVAL_44) begin
      if (_EVAL_57) begin
        _EVAL_137 <= 1'h0;
      end else begin
        _EVAL_137 <= _EVAL_78;
      end
    end
    if (_EVAL_227) begin
      _EVAL_149 <= _EVAL_12;
    end
    if (_EVAL) begin
      _EVAL_155 <= 5'h0;
    end else begin
      _EVAL_155 <= _EVAL_115;
    end
    if (_EVAL) begin
      _EVAL_173 <= 32'h0;
    end else if (_EVAL_151) begin
      _EVAL_173 <= 32'h0;
    end else begin
      _EVAL_173 <= _EVAL_166;
    end
    if (_EVAL_150) begin
      _EVAL_201 <= _EVAL_5;
    end
    if (_EVAL) begin
      _EVAL_215 <= 1'h0;
    end else if (_EVAL_212) begin
      if (_EVAL_213) begin
        _EVAL_215 <= 1'h0;
      end else begin
        _EVAL_215 <= _EVAL_64;
      end
    end
    if (_EVAL) begin
      _EVAL_238 <= 1'h0;
    end else if (_EVAL_44) begin
      if (_EVAL_233) begin
        _EVAL_238 <= 1'h0;
      end else begin
        _EVAL_238 <= _EVAL_226;
      end
    end
    if (_EVAL_227) begin
      _EVAL_245 <= _EVAL_8;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25531acb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b68f5572)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91fe0ff3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(874c249b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cd7a948)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa07a1db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7bff0e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47c62ed1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f839033)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fc6f4a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(426609ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e1d76bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d142cdb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e3ededa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d13b3668)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93c924bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9507db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca60b184)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a727e7ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2289fa49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac4f316d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac221499)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d538f979)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1285dbe7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f39f19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(629eca36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17fb72cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a363b48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a36ec6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc5241d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd0cedba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8f9bffb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db8ef96e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c7c0479)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53a42092)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dae8ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99800631)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e83a3f85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe378ad2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed15cdb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63f5f684)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be646378)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecb66f8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a67002d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f55abd0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e698479a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7bea7b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca0a9591)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93dbf033)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37945f82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43e16498)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2337e47f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59791d1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f51e3a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3409ccd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4079a7a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd3d0482)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0f736da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6e38063)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b27e69f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b6f8952)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7863406f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c512fb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa817192)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bf1268c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2e23a30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7601a13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7729445)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17ef0836)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4179e682)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fcdc29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f07af8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eab9bb4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
