//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_68_assert(
  input         _EVAL,
  input  [3:0]  _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input  [29:0] _EVAL_8,
  input  [1:0]  _EVAL_9,
  input         _EVAL_10,
  input  [3:0]  _EVAL_11,
  input         _EVAL_12,
  input  [3:0]  _EVAL_13,
  input  [2:0]  _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18
);
  wire  _EVAL_19;
  wire [3:0] _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire [7:0] _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire [7:0] _EVAL_30;
  wire  _EVAL_31;
  wire [29:0] _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire [30:0] _EVAL_35;
  wire  _EVAL_36;
  wire [1:0] _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire [6:0] _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire [30:0] _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_61;
  wire [30:0] _EVAL_63;
  wire  _EVAL_64;
  wire [7:0] _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire [30:0] _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  reg [2:0] _EVAL_78;
  reg [31:0] _RAND_0;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire [4:0] _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire [22:0] _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire [32:0] _EVAL_117;
  wire  _EVAL_118;
  reg [2:0] _EVAL_119;
  reg [31:0] _RAND_1;
  wire  _EVAL_120;
  wire [30:0] _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire [4:0] _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire [5:0] _EVAL_134;
  wire  _EVAL_135;
  reg [3:0] _EVAL_136;
  reg [31:0] _RAND_2;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire [4:0] _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire [31:0] _EVAL_146;
  wire [29:0] _EVAL_147;
  reg [2:0] _EVAL_148;
  reg [31:0] _RAND_3;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire [30:0] _EVAL_152;
  wire [29:0] _EVAL_153;
  wire  _EVAL_154;
  reg [31:0] _EVAL_155;
  reg [31:0] _RAND_4;
  wire [31:0] plusarg_reader_out;
  wire [5:0] _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  reg [5:0] _EVAL_162;
  reg [31:0] _RAND_5;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire [30:0] _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire [7:0] _EVAL_172;
  wire  _EVAL_173;
  reg [2:0] _EVAL_174;
  reg [31:0] _RAND_6;
  wire [22:0] _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  reg [29:0] _EVAL_179;
  reg [31:0] _RAND_7;
  wire  _EVAL_180;
  wire [5:0] _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  reg [5:0] _EVAL_193;
  reg [31:0] _RAND_8;
  reg [5:0] _EVAL_194;
  reg [31:0] _RAND_9;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  reg [1:0] _EVAL_202;
  reg [31:0] _RAND_10;
  wire  _EVAL_204;
  wire [4:0] _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire [30:0] _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire [5:0] _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire [1:0] _EVAL_217;
  wire [7:0] _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire [30:0] _EVAL_222;
  wire [4:0] _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire [7:0] _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire [3:0] _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire [29:0] _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire [4:0] _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire [5:0] _EVAL_248;
  wire  _EVAL_249;
  wire [6:0] _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire [6:0] _EVAL_254;
  wire [29:0] _EVAL_255;
  wire  _EVAL_256;
  wire [30:0] _EVAL_257;
  wire [1:0] _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  reg [3:0] _EVAL_262;
  reg [31:0] _RAND_11;
  wire  _EVAL_263;
  wire [1:0] _EVAL_264;
  reg [5:0] _EVAL_265;
  reg [31:0] _RAND_12;
  wire  _EVAL_266;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire [30:0] _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire [4:0] _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire [7:0] _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire [30:0] _EVAL_287;
  wire [3:0] _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire [7:0] _EVAL_296;
  wire [4:0] _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire [3:0] _EVAL_301;
  wire  _EVAL_302;
  reg [4:0] _EVAL_303;
  reg [31:0] _RAND_13;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire [6:0] _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire [5:0] _EVAL_312;
  wire  _EVAL_313;
  reg  _EVAL_314;
  reg [31:0] _RAND_14;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  reg [2:0] _EVAL_318;
  reg [31:0] _RAND_15;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire  _EVAL_321;
  reg  _EVAL_322;
  reg [31:0] _RAND_16;
  wire  _EVAL_323;
  wire  _EVAL_324;
  wire  _EVAL_325;
  wire  _EVAL_326;
  wire  _EVAL_327;
  wire  _EVAL_328;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_178 = _EVAL_76 | _EVAL_16;
  assign _EVAL_277 = _EVAL_212 & _EVAL_216;
  assign _EVAL_20 = _EVAL_13 & _EVAL_230;
  assign _EVAL_150 = _EVAL_5 == 3'h3;
  assign _EVAL_55 = _EVAL_19 | _EVAL_16;
  assign _EVAL_248 = _EVAL_250[5:0];
  assign _EVAL_118 = _EVAL_42 | _EVAL_277;
  assign _EVAL_327 = _EVAL_212 & _EVAL_204;
  assign _EVAL_292 = plusarg_reader_out == 32'h0;
  assign _EVAL_56 = _EVAL_165 | _EVAL_229;
  assign _EVAL_165 = _EVAL_201 | _EVAL_98;
  assign _EVAL_139 = ~_EVAL_79;
  assign _EVAL_93 = ~_EVAL_192;
  assign _EVAL_187 = ~_EVAL_286;
  assign _EVAL_167 = $signed(_EVAL_287) & -31'sh2000;
  assign _EVAL_210 = _EVAL_9 != 2'h2;
  assign _EVAL_296 = _EVAL_108 ? _EVAL_227 : 8'h0;
  assign _EVAL_182 = _EVAL_11 <= 4'h8;
  assign _EVAL_217 = _EVAL_1[2:1];
  assign _EVAL_57 = ~_EVAL_12;
  assign _EVAL_107 = ~_EVAL_249;
  assign _EVAL_44 = _EVAL_193 - 6'h1;
  assign _EVAL_309 = _EVAL_162 - 6'h1;
  assign _EVAL_306 = _EVAL_20 == 4'h0;
  assign _EVAL_85 = $signed(_EVAL_70) == 31'sh0;
  assign _EVAL_190 = ~_EVAL_48;
  assign _EVAL_195 = _EVAL_4 == 3'h0;
  assign _EVAL_245 = ~_EVAL_313;
  assign _EVAL_244 = _EVAL_242 | _EVAL_16;
  assign _EVAL_89 = _EVAL_265 == 6'h0;
  assign _EVAL_275 = _EVAL_223 & _EVAL_205;
  assign _EVAL_175 = 23'hff << _EVAL_11;
  assign _EVAL_168 = _EVAL_75 | _EVAL_16;
  assign _EVAL_288 = ~_EVAL_13;
  assign _EVAL_240 = _EVAL_54 | _EVAL_80;
  assign _EVAL_316 = _EVAL_59 & _EVAL_282;
  assign _EVAL_100 = _EVAL_2 & _EVAL_96;
  assign _EVAL_142 = _EVAL_81 | _EVAL_303;
  assign _EVAL_220 = _EVAL_32 == 30'h0;
  assign _EVAL_235 = _EVAL_283 | _EVAL_16;
  assign _EVAL_312 = _EVAL_23[7:2];
  assign _EVAL_180 = _EVAL_106 | _EVAL_12;
  assign _EVAL_238 = ~_EVAL_86;
  assign _EVAL_219 = ~_EVAL_69;
  assign _EVAL_177 = _EVAL_5 == 3'h4;
  assign _EVAL_124 = ~_EVAL_304;
  assign _EVAL_65 = _EVAL_120 ? _EVAL_218 : 8'h0;
  assign _EVAL_205 = ~_EVAL_126;
  assign _EVAL_84 = _EVAL_268 | _EVAL_239;
  assign _EVAL_67 = _EVAL_5 == 3'h6;
  assign _EVAL_72 = ~_EVAL_131;
  assign _EVAL_36 = _EVAL_206 & _EVAL_260;
  assign _EVAL_95 = ~_EVAL_320;
  assign _EVAL_29 = ~_EVAL_149;
  assign _EVAL_70 = _EVAL_63;
  assign _EVAL_200 = ~_EVAL_294;
  assign _EVAL_241 = _EVAL_142 >> _EVAL_1;
  assign _EVAL_50 = $signed(_EVAL_222) & -31'sh1000000;
  assign _EVAL_37 = _EVAL_3[2:1];
  assign _EVAL_161 = _EVAL_5 == 3'h7;
  assign _EVAL_117 = _EVAL_155 + 32'h1;
  assign _EVAL_176 = _EVAL_271 | _EVAL_88;
  assign _EVAL_52 = _EVAL_14 == 3'h0;
  assign _EVAL_130 = _EVAL_212 & _EVAL_138;
  assign _EVAL_221 = _EVAL_8[0];
  assign _EVAL_160 = _EVAL_144 | _EVAL_16;
  assign _EVAL_27 = ~_EVAL_231;
  assign _EVAL_259 = ~_EVAL_6;
  assign _EVAL_74 = _EVAL_5 == 3'h0;
  assign _EVAL_222 = {1'b0,$signed(_EVAL_147)};
  assign _EVAL_40 = _EVAL_2 & _EVAL_247;
  assign _EVAL_228 = _EVAL_9 == 2'h0;
  assign _EVAL_310 = ~_EVAL_61;
  assign _EVAL_104 = ~_EVAL_102;
  assign _EVAL_189 = _EVAL_37 == 2'h0;
  assign _EVAL_214 = _EVAL_217 == 2'h1;
  assign _EVAL_326 = ~_EVAL_235;
  assign _EVAL_311 = _EVAL_4 <= 3'h4;
  assign _EVAL_63 = $signed(_EVAL_270) & -31'sh5000;
  assign _EVAL_99 = _EVAL_264[1];
  assign _EVAL_35 = _EVAL_50;
  assign _EVAL_138 = _EVAL_125 | _EVAL_85;
  assign _EVAL_321 = _EVAL_272 | _EVAL_295;
  assign _EVAL_111 = ~_EVAL_55;
  assign _EVAL_42 = _EVAL_182 & _EVAL_269;
  assign _EVAL_204 = _EVAL_138 | _EVAL_216;
  assign _EVAL_283 = _EVAL_14 <= 3'h6;
  assign _EVAL_38 = _EVAL_116 | _EVAL_310;
  assign _EVAL_43 = _EVAL_1 == _EVAL_119;
  assign _EVAL_172 = ~_EVAL_280;
  assign _EVAL_225 = ~_EVAL_168;
  assign _EVAL_268 = _EVAL_289 | _EVAL_189;
  assign _EVAL_157 = _EVAL_254[5:0];
  assign _EVAL_307 = _EVAL_18 & _EVAL_31;
  assign _EVAL_302 = _EVAL_5[2];
  assign _EVAL_208 = _EVAL_165 | _EVAL_316;
  assign _EVAL_23 = ~_EVAL_30;
  assign _EVAL_164 = ~_EVAL_266;
  assign _EVAL_183 = _EVAL_18 & _EVAL_67;
  assign _EVAL_247 = ~_EVAL_260;
  assign _EVAL_252 = _EVAL_14 == 3'h5;
  assign _EVAL_256 = _EVAL_2 & _EVAL_300;
  assign _EVAL_125 = $signed(_EVAL_35) == 31'sh0;
  assign _EVAL_80 = _EVAL_1 == 3'h4;
  assign _EVAL_170 = _EVAL_18 & _EVAL_150;
  assign _EVAL_31 = ~_EVAL_196;
  assign _EVAL_58 = _EVAL_99 & _EVAL_45;
  assign _EVAL_21 = _EVAL_193 == 6'h0;
  assign _EVAL_243 = _EVAL_217 == 2'h0;
  assign _EVAL_171 = ~_EVAL_244;
  assign _EVAL_215 = _EVAL_18 & _EVAL_177;
  assign _EVAL_297 = _EVAL_303 >> _EVAL_3;
  assign _EVAL_264 = _EVAL_258 | 2'h1;
  assign _EVAL_258 = 2'h1 << _EVAL_25;
  assign _EVAL_293 = _EVAL_180 | _EVAL_16;
  assign _EVAL_131 = _EVAL_305 | _EVAL_16;
  assign _EVAL_46 = _EVAL_195 | _EVAL_16;
  assign _EVAL_260 = _EVAL_194 == 6'h0;
  assign _EVAL_276 = _EVAL_272 | _EVAL_191;
  assign _EVAL_216 = $signed(_EVAL_121) == 31'sh0;
  assign _EVAL_324 = _EVAL_154 | _EVAL_85;
  assign _EVAL_199 = _EVAL_151 | _EVAL_16;
  assign _EVAL_113 = ~_EVAL_185;
  assign _EVAL_48 = _EVAL_91 | _EVAL_16;
  assign _EVAL_33 = _EVAL_241[0];
  assign _EVAL_163 = _EVAL_297[0];
  assign _EVAL_280 = _EVAL_109[7:0];
  assign _EVAL_69 = _EVAL_220 | _EVAL_16;
  assign _EVAL_266 = _EVAL_166 | _EVAL_16;
  assign _EVAL_141 = ~_EVAL_188;
  assign _EVAL_305 = ~_EVAL_163;
  assign _EVAL_323 = _EVAL_18 & _EVAL_132;
  assign _EVAL_140 = ~_EVAL_207;
  assign _EVAL_191 = _EVAL_59 & _EVAL_273;
  assign _EVAL_92 = _EVAL_115 | _EVAL_16;
  assign _EVAL_273 = _EVAL_45 & _EVAL_145;
  assign _EVAL_246 = ~_EVAL_160;
  assign _EVAL_317 = _EVAL_274 & _EVAL_145;
  assign _EVAL_137 = ~_EVAL_129;
  assign _EVAL_66 = _EVAL_4 == _EVAL_148;
  assign _EVAL_281 = ~_EVAL_71;
  assign _EVAL_207 = _EVAL_303 != 5'h0;
  assign _EVAL_79 = _EVAL_328 | _EVAL_16;
  assign _EVAL_300 = _EVAL_14 == 3'h4;
  assign _EVAL_213 = _EVAL_44[5:0];
  assign _EVAL_284 = ~_EVAL_263;
  assign _EVAL_22 = _EVAL_236 | _EVAL_16;
  assign _EVAL_209 = {1'b0,$signed(_EVAL_233)};
  assign _EVAL_282 = _EVAL_274 & _EVAL_221;
  assign _EVAL_132 = _EVAL_5 == 3'h5;
  assign _EVAL_75 = _EVAL_5 == _EVAL_78;
  assign _EVAL_234 = _EVAL_18 & _EVAL_261;
  assign _EVAL_101 = ~_EVAL_278;
  assign _EVAL_301 = {_EVAL_321,_EVAL_276,_EVAL_208,_EVAL_56};
  assign _EVAL_298 = _EVAL_5 == 3'h1;
  assign _EVAL_86 = _EVAL_325 | _EVAL_16;
  assign _EVAL_242 = _EVAL_3 == _EVAL_174;
  assign _EVAL_227 = 8'h1 << _EVAL_1;
  assign _EVAL_53 = _EVAL_240 | _EVAL_16;
  assign _EVAL_291 = ~_EVAL_169;
  assign _EVAL_77 = ~_EVAL_143;
  assign _EVAL_255 = _EVAL_8 ^ 30'h20000000;
  assign _EVAL_278 = _EVAL_158 | _EVAL_16;
  assign _EVAL_263 = _EVAL_159 | _EVAL_16;
  assign _EVAL_120 = _EVAL_122 & _EVAL_21;
  assign _EVAL_24 = ~_EVAL_22;
  assign _EVAL_237 = ~_EVAL_112;
  assign _EVAL_133 = _EVAL_18 & _EVAL_161;
  assign _EVAL_146 = _EVAL_117[31:0];
  assign _EVAL_34 = _EVAL_2 & _EVAL_320;
  assign _EVAL_71 = _EVAL_118 | _EVAL_16;
  assign _EVAL_270 = {1'b0,$signed(_EVAL_8)};
  assign _EVAL_218 = 8'h1 << _EVAL_3;
  assign _EVAL_249 = _EVAL_311 | _EVAL_16;
  assign _EVAL_287 = {1'b0,$signed(_EVAL_255)};
  assign _EVAL_274 = ~_EVAL_45;
  assign _EVAL_295 = _EVAL_59 & _EVAL_232;
  assign _EVAL_290 = _EVAL_43 | _EVAL_16;
  assign _EVAL_106 = ~_EVAL;
  assign _EVAL_102 = _EVAL_197 | _EVAL_16;
  assign _EVAL_197 = _EVAL_4 <= 3'h1;
  assign _EVAL_250 = _EVAL_265 - 6'h1;
  assign _EVAL_271 = _EVAL_140 | _EVAL_292;
  assign _EVAL_328 = _EVAL_13 == _EVAL_301;
  assign _EVAL_299 = _EVAL_206 & _EVAL_89;
  assign _EVAL_87 = ~_EVAL_302;
  assign _EVAL_198 = _EVAL_2 & _EVAL_52;
  assign _EVAL_32 = _EVAL_8 & _EVAL_153;
  assign _EVAL_144 = _EVAL_288 == 4'h0;
  assign _EVAL_212 = _EVAL_11 <= 4'h2;
  assign _EVAL_233 = _EVAL_8 ^ 30'h3000;
  assign _EVAL_158 = _EVAL_11 == _EVAL_136;
  assign _EVAL_129 = _EVAL_210 | _EVAL_16;
  assign _EVAL_320 = _EVAL_14 == 3'h6;
  assign _EVAL_110 = _EVAL_14 == _EVAL_318;
  assign _EVAL_169 = _EVAL_39 | _EVAL_16;
  assign _EVAL_229 = _EVAL_59 & _EVAL_317;
  assign _EVAL_123 = ~_EVAL_82;
  assign _EVAL_152 = $signed(_EVAL_209) & -31'sh1000;
  assign _EVAL_185 = _EVAL_201 | _EVAL_16;
  assign _EVAL_109 = 23'hff << _EVAL_0;
  assign _EVAL_184 = _EVAL_2 & _EVAL_127;
  assign _EVAL_159 = _EVAL_17 == _EVAL_314;
  assign _EVAL_181 = _EVAL_172[7:2];
  assign _EVAL_76 = _EVAL_212 & _EVAL_28;
  assign _EVAL_153 = {{22'd0}, _EVAL_23};
  assign _EVAL_232 = _EVAL_45 & _EVAL_221;
  assign _EVAL_223 = _EVAL_303 | _EVAL_81;
  assign _EVAL_96 = _EVAL_14 == 3'h2;
  assign _EVAL_25 = _EVAL_11[0];
  assign _EVAL_143 = _EVAL_49 | _EVAL_16;
  assign _EVAL_192 = _EVAL_176 | _EVAL_16;
  assign _EVAL_230 = ~_EVAL_301;
  assign _EVAL_166 = _EVAL_4 != 3'h0;
  assign _EVAL_239 = _EVAL_3 == 3'h4;
  assign _EVAL_285 = _EVAL_122 | _EVAL_206;
  assign _EVAL_127 = _EVAL_14 == 3'h1;
  assign _EVAL_98 = _EVAL_99 & _EVAL_274;
  assign _EVAL_97 = _EVAL_14[0];
  assign _EVAL_114 = ~_EVAL_83;
  assign _EVAL_254 = _EVAL_194 - 6'h1;
  assign _EVAL_126 = _EVAL_296[4:0];
  assign _EVAL_19 = _EVAL_0 >= 4'h2;
  assign _EVAL_319 = ~_EVAL_199;
  assign _EVAL_294 = _EVAL_33 | _EVAL_16;
  assign _EVAL_196 = _EVAL_162 == 6'h0;
  assign _EVAL_186 = ~_EVAL_293;
  assign _EVAL_272 = _EVAL_201 | _EVAL_58;
  assign _EVAL_211 = _EVAL_106 | _EVAL_16;
  assign _EVAL_261 = _EVAL_5 == 3'h2;
  assign _EVAL_251 = _EVAL_18 & _EVAL_74;
  assign _EVAL_121 = _EVAL_167;
  assign _EVAL_28 = _EVAL_324 | _EVAL_216;
  assign _EVAL_49 = _EVAL == _EVAL_322;
  assign _EVAL_257 = _EVAL_152;
  assign _EVAL_41 = _EVAL_51 | _EVAL_16;
  assign _EVAL_88 = _EVAL_155 < plusarg_reader_out;
  assign _EVAL_45 = _EVAL_8[1];
  assign _EVAL_73 = _EVAL_2 & _EVAL_252;
  assign _EVAL_54 = _EVAL_214 | _EVAL_243;
  assign _EVAL_51 = _EVAL_4 <= 3'h3;
  assign _EVAL_154 = _EVAL_269 | _EVAL_125;
  assign _EVAL_115 = _EVAL_4 <= 3'h2;
  assign _EVAL_103 = ~_EVAL_46;
  assign _EVAL_188 = _EVAL_259 | _EVAL_16;
  assign _EVAL_147 = _EVAL_8 ^ 30'h2000000;
  assign _EVAL_134 = _EVAL_309[5:0];
  assign _EVAL_253 = _EVAL_122 & _EVAL_196;
  assign _EVAL_68 = ~_EVAL_211;
  assign _EVAL_39 = _EVAL_42 | _EVAL_130;
  assign _EVAL_122 = _EVAL_15 & _EVAL_18;
  assign _EVAL_286 = _EVAL_84 | _EVAL_16;
  assign _EVAL_149 = _EVAL_66 | _EVAL_16;
  assign _EVAL_201 = _EVAL_11 >= 4'h2;
  assign _EVAL_236 = _EVAL_9 <= 2'h2;
  assign _EVAL_90 = _EVAL_9 == _EVAL_202;
  assign _EVAL_313 = _EVAL_38 | _EVAL_16;
  assign _EVAL_289 = _EVAL_37 == 2'h1;
  assign _EVAL_226 = ~_EVAL_92;
  assign _EVAL_64 = _EVAL_18 & _EVAL_298;
  assign _EVAL_61 = _EVAL_81 != 5'h0;
  assign _EVAL_135 = ~_EVAL_16;
  assign _EVAL_116 = _EVAL_81 != _EVAL_126;
  assign _EVAL_112 = _EVAL_306 | _EVAL_16;
  assign _EVAL_224 = ~_EVAL_53;
  assign _EVAL_108 = _EVAL_299 & _EVAL_95;
  assign _EVAL_81 = _EVAL_65[4:0];
  assign _EVAL_128 = ~_EVAL_290;
  assign _EVAL_231 = _EVAL_228 | _EVAL_16;
  assign _EVAL_59 = _EVAL_264[0];
  assign _EVAL_30 = _EVAL_175[7:0];
  assign _EVAL_173 = ~_EVAL_178;
  assign _EVAL_206 = _EVAL_10 & _EVAL_2;
  assign _EVAL_269 = $signed(_EVAL_257) == 31'sh0;
  assign _EVAL_83 = _EVAL_110 | _EVAL_16;
  assign _EVAL_304 = _EVAL_90 | _EVAL_16;
  assign _EVAL_151 = _EVAL_0 == _EVAL_262;
  assign _EVAL_82 = _EVAL_57 | _EVAL_16;
  assign _EVAL_325 = _EVAL_42 | _EVAL_327;
  assign _EVAL_315 = ~_EVAL_41;
  assign _EVAL_91 = _EVAL_8 == _EVAL_179;
  assign _EVAL_145 = ~_EVAL_221;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_78 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_119 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_136 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_148 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_155 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_162 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_174 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_179 = _RAND_7[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_193 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_194 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_202 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_262 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_265 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_303 = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_314 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_318 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_322 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_7) begin
    if (_EVAL_253) begin
      _EVAL_78 <= _EVAL_5;
    end
    if (_EVAL_36) begin
      _EVAL_119 <= _EVAL_1;
    end
    if (_EVAL_253) begin
      _EVAL_136 <= _EVAL_11;
    end
    if (_EVAL_253) begin
      _EVAL_148 <= _EVAL_4;
    end
    if (_EVAL_16) begin
      _EVAL_155 <= 32'h0;
    end else if (_EVAL_285) begin
      _EVAL_155 <= 32'h0;
    end else begin
      _EVAL_155 <= _EVAL_146;
    end
    if (_EVAL_16) begin
      _EVAL_162 <= 6'h0;
    end else if (_EVAL_122) begin
      if (_EVAL_196) begin
        if (_EVAL_87) begin
          _EVAL_162 <= _EVAL_312;
        end else begin
          _EVAL_162 <= 6'h0;
        end
      end else begin
        _EVAL_162 <= _EVAL_134;
      end
    end
    if (_EVAL_253) begin
      _EVAL_174 <= _EVAL_3;
    end
    if (_EVAL_253) begin
      _EVAL_179 <= _EVAL_8;
    end
    if (_EVAL_16) begin
      _EVAL_193 <= 6'h0;
    end else if (_EVAL_122) begin
      if (_EVAL_21) begin
        if (_EVAL_87) begin
          _EVAL_193 <= _EVAL_312;
        end else begin
          _EVAL_193 <= 6'h0;
        end
      end else begin
        _EVAL_193 <= _EVAL_213;
      end
    end
    if (_EVAL_16) begin
      _EVAL_194 <= 6'h0;
    end else if (_EVAL_206) begin
      if (_EVAL_260) begin
        if (_EVAL_97) begin
          _EVAL_194 <= _EVAL_181;
        end else begin
          _EVAL_194 <= 6'h0;
        end
      end else begin
        _EVAL_194 <= _EVAL_157;
      end
    end
    if (_EVAL_36) begin
      _EVAL_202 <= _EVAL_9;
    end
    if (_EVAL_36) begin
      _EVAL_262 <= _EVAL_0;
    end
    if (_EVAL_16) begin
      _EVAL_265 <= 6'h0;
    end else if (_EVAL_206) begin
      if (_EVAL_89) begin
        if (_EVAL_97) begin
          _EVAL_265 <= _EVAL_181;
        end else begin
          _EVAL_265 <= 6'h0;
        end
      end else begin
        _EVAL_265 <= _EVAL_248;
      end
    end
    if (_EVAL_16) begin
      _EVAL_303 <= 5'h0;
    end else begin
      _EVAL_303 <= _EVAL_275;
    end
    if (_EVAL_36) begin
      _EVAL_314 <= _EVAL_17;
    end
    if (_EVAL_36) begin
      _EVAL_318 <= _EVAL_14;
    end
    if (_EVAL_36) begin
      _EVAL_322 <= _EVAL;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6f53541)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d978793)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3646731d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41eb4c4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90462bf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b23a1438)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6b61ffa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(313da8f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ffc4745)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_284) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33f76c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af68d4fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1f93038)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4680104e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(823f3ee5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_326) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a44f09b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fe79116)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aab94b5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(779f3049)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9e4b0d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e855e76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e611be7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cb82c46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9db7fb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74deb43d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edfbdf44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(444124fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69d3747d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ab0f300)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d571e0e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_315) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3398e15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e50ce45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c986fd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b9fd994)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12a28a27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24bcd191)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7dee780d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(707facad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8871216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f34b233)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77657903)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51f0d0e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51cc2e56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ec0b68f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_319) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4aa4adff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0804dcf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d6d5cbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5477e2b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0f794a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90add815)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb419481)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ab9fc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_326) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40bcc523)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3899a543)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7551a132)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_315) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27884d66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36deb12c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2759ebe1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e558afe6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e586387)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32fd271f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54e711d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a5a596)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad9538bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7dd5fd65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_284) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e7c054e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f0fbbff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e7935bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(706963ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0b44d58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69c64524)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cec438b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(975e6892)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf216331)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebf149db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3047b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_319) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3ff4a5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1cfd66c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3624f1bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cad08fb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d1b7c61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37f78014)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4034538)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dfe948f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0e30cb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95f4742a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67408174)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(711b348)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b05f66f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(563b975b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27992035)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e39e5cee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
