//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_120_assert(
  input        _EVAL,
  input        _EVAL_0,
  input  [3:0] _EVAL_1,
  input        _EVAL_2,
  input  [2:0] _EVAL_3,
  input  [6:0] _EVAL_4,
  input  [2:0] _EVAL_5,
  input        _EVAL_6,
  input        _EVAL_7,
  input        _EVAL_8
);
  wire  _EVAL_9;
  reg  _EVAL_10;
  reg [31:0] _RAND_0;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_11;
  wire  _EVAL_12;
  wire  _EVAL_13;
  wire  _EVAL_14;
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  reg [2:0] _EVAL_19;
  reg [31:0] _RAND_1;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire [1:0] _EVAL_24;
  wire [7:0] _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  reg [2:0] _EVAL_30;
  reg [31:0] _RAND_2;
  wire  _EVAL_31;
  reg [31:0] _EVAL_32;
  reg [31:0] _RAND_3;
  wire  _EVAL_33;
  wire  _EVAL_34;
  reg [6:0] _EVAL_35;
  reg [31:0] _RAND_4;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire [1:0] _EVAL_45;
  wire [6:0] _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire [7:0] _EVAL_53;
  wire [1:0] _EVAL_54;
  wire  _EVAL_55;
  wire [1:0] _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire [7:0] _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire [31:0] _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire [1:0] _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  reg  _EVAL_78;
  reg [31:0] _RAND_5;
  wire  _EVAL_79;
  reg  _EVAL_80;
  reg [31:0] _RAND_6;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire [7:0] _EVAL_83;
  wire  _EVAL_84;
  wire [7:0] _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  reg  _EVAL_90;
  reg [31:0] _RAND_7;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire [7:0] _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire [6:0] _EVAL_98;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire [6:0] _EVAL_103;
  wire [1:0] _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  reg  _EVAL_109;
  reg [31:0] _RAND_8;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire [32:0] _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire [3:0] _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_77 = ~_EVAL_49;
  assign _EVAL_28 = _EVAL_4 == _EVAL_35;
  assign _EVAL_75 = _EVAL_6;
  assign _EVAL_17 = _EVAL & _EVAL_7;
  assign _EVAL_94 = _EVAL_24[0];
  assign _EVAL_107 = $signed(_EVAL_53) == 8'sh0;
  assign _EVAL_49 = _EVAL_65 | _EVAL_75;
  assign _EVAL_21 = ~_EVAL_9;
  assign _EVAL_34 = _EVAL_54[0];
  assign _EVAL_70 = _EVAL_3 <= 3'h6;
  assign _EVAL_64 = _EVAL_17 & _EVAL_108;
  assign _EVAL_16 = plusarg_reader_out == 32'h0;
  assign _EVAL_102 = ~_EVAL_20;
  assign _EVAL_101 = _EVAL_7 & _EVAL_71;
  assign _EVAL_121 = _EVAL_7 & _EVAL_82;
  assign _EVAL_81 = _EVAL_5 == 3'h7;
  assign _EVAL_95 = $signed(_EVAL_62) & -8'sh14;
  assign _EVAL_13 = _EVAL_22 & _EVAL_21;
  assign _EVAL_108 = ~_EVAL_78;
  assign _EVAL_79 = ~_EVAL_106;
  assign _EVAL_39 = ~_EVAL_113;
  assign _EVAL_11 = _EVAL_120 | _EVAL_27;
  assign _EVAL_63 = _EVAL_0 & _EVAL_73;
  assign _EVAL_27 = _EVAL_32 < plusarg_reader_out;
  assign _EVAL_42 = ~_EVAL_75;
  assign _EVAL_52 = ~_EVAL_94;
  assign _EVAL_58 = _EVAL_7 & _EVAL_44;
  assign _EVAL_85 = _EVAL_95;
  assign _EVAL_67 = _EVAL_114[31:0];
  assign _EVAL_31 = _EVAL_2 & _EVAL_0;
  assign _EVAL_92 = _EVAL_5 == 3'h4;
  assign _EVAL_51 = _EVAL_5 == 3'h0;
  assign _EVAL_57 = ~_EVAL_23;
  assign _EVAL_43 = ~_EVAL_80;
  assign _EVAL_53 = _EVAL_83;
  assign _EVAL_123 = ~_EVAL_108;
  assign _EVAL_98 = _EVAL_4 & 7'h3;
  assign _EVAL_113 = _EVAL_74 | _EVAL_75;
  assign _EVAL_54 = _EVAL_80 - 1'h1;
  assign _EVAL_37 = ~_EVAL_10;
  assign _EVAL_46 = _EVAL_4 ^ 7'h40;
  assign _EVAL_25 = {1'b0,$signed(_EVAL_103)};
  assign _EVAL_12 = _EVAL_11 | _EVAL_75;
  assign _EVAL_36 = _EVAL_7 & _EVAL_40;
  assign _EVAL_115 = _EVAL_17 | _EVAL_31;
  assign _EVAL_87 = _EVAL_7 & _EVAL_81;
  assign _EVAL_103 = _EVAL_4 ^ 7'h54;
  assign _EVAL_45 = _EVAL_78 - 1'h1;
  assign _EVAL_125 = _EVAL_1 == 4'hf;
  assign _EVAL_124 = _EVAL_72[0];
  assign _EVAL_73 = ~_EVAL_37;
  assign _EVAL_89 = _EVAL_0 & _EVAL_84;
  assign _EVAL_71 = _EVAL_5 == 3'h6;
  assign _EVAL_62 = {1'b0,$signed(_EVAL_46)};
  assign _EVAL_84 = _EVAL_3 == 3'h5;
  assign _EVAL_23 = _EVAL_91 | _EVAL_75;
  assign _EVAL_100 = _EVAL_7 & _EVAL_119;
  assign _EVAL_120 = _EVAL_74 | _EVAL_16;
  assign _EVAL_104 = _EVAL_93 ? 2'h1 : 2'h0;
  assign _EVAL_91 = _EVAL_122 == 4'h0;
  assign _EVAL_9 = _EVAL_3 == 3'h6;
  assign _EVAL_26 = ~_EVAL_88;
  assign _EVAL_68 = _EVAL_28 | _EVAL_75;
  assign _EVAL_40 = _EVAL_5 == 3'h5;
  assign _EVAL_66 = ~_EVAL_38;
  assign _EVAL_119 = _EVAL_5 == 3'h3;
  assign _EVAL_33 = ~_EVAL_90;
  assign _EVAL_117 = ~_EVAL_76;
  assign _EVAL_97 = _EVAL_7 & _EVAL_51;
  assign _EVAL_122 = ~_EVAL_1;
  assign _EVAL_47 = ~_EVAL_14;
  assign _EVAL_86 = _EVAL_7 & _EVAL_92;
  assign _EVAL_111 = _EVAL_104[0];
  assign _EVAL_44 = _EVAL_5 == 3'h1;
  assign _EVAL_60 = _EVAL_0 & _EVAL_110;
  assign _EVAL_29 = ~_EVAL_68;
  assign _EVAL_59 = $signed(_EVAL_85) == 8'sh0;
  assign _EVAL_93 = _EVAL_17 & _EVAL_43;
  assign _EVAL_106 = _EVAL_105 | _EVAL_75;
  assign _EVAL_18 = _EVAL_56[0];
  assign _EVAL_72 = _EVAL_90 - 1'h1;
  assign _EVAL_116 = _EVAL_59 | _EVAL_107;
  assign _EVAL_114 = _EVAL_32 + 32'h1;
  assign _EVAL_55 = _EVAL_109 | _EVAL_111;
  assign _EVAL_76 = _EVAL_70 | _EVAL_75;
  assign _EVAL_20 = _EVAL_112 | _EVAL_75;
  assign _EVAL_56 = _EVAL_10 - 1'h1;
  assign _EVAL_38 = _EVAL_15 | _EVAL_75;
  assign _EVAL_96 = _EVAL_31 & _EVAL_37;
  assign _EVAL_74 = ~_EVAL_109;
  assign _EVAL_61 = _EVAL_45[0];
  assign _EVAL_15 = _EVAL_111 | _EVAL_109;
  assign _EVAL_82 = _EVAL_5 == 3'h2;
  assign _EVAL_112 = _EVAL_98 == 7'h0;
  assign _EVAL_50 = ~_EVAL_12;
  assign _EVAL_65 = _EVAL_3 == _EVAL_30;
  assign _EVAL_110 = _EVAL_3 == 3'h4;
  assign _EVAL_118 = _EVAL_7 & _EVAL_123;
  assign _EVAL_105 = _EVAL_5 == _EVAL_19;
  assign _EVAL_22 = _EVAL_31 & _EVAL_33;
  assign _EVAL_14 = _EVAL_116 | _EVAL_75;
  assign _EVAL_83 = $signed(_EVAL_25) & -8'sh4;
  assign _EVAL_24 = _EVAL_13 ? 2'h1 : 2'h0;
  assign _EVAL_88 = _EVAL_125 | _EVAL_75;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_10 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_19 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_30 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_32 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_35 = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_78 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_80 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_90 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_109 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  if (_EVAL_6) begin
    _EVAL_10 = 1'h0;
  end
  if (_EVAL_6) begin
    _EVAL_32 = 32'h0;
  end
  if (_EVAL_6) begin
    _EVAL_78 = 1'h0;
  end
  if (_EVAL_6) begin
    _EVAL_80 = 1'h0;
  end
  if (_EVAL_6) begin
    _EVAL_90 = 1'h0;
  end
  if (_EVAL_6) begin
    _EVAL_109 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_8) begin
    if (_EVAL_64) begin
      _EVAL_19 <= _EVAL_5;
    end
    if (_EVAL_96) begin
      _EVAL_30 <= _EVAL_3;
    end
    if (_EVAL_64) begin
      _EVAL_35 <= _EVAL_4;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f03c93db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f12c637b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e896bfd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(716e875f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9330054)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbded0c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0b5db0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(689826d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f35a4a67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dd3e621)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d3359)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7485c1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3faced2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cce52d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e664d71b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88a50af8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fcfe327)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca09b8e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb86bb3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2178fd8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29053e33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4611982e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8209ca7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48eb767f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9e328fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be2d9bae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_66) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff3b360c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49ce3bfc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65e5c2da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2ca9b17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b61d8023)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9902ab1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b598ee9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_66) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dbc1628)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b0987cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge _EVAL_8 or posedge _EVAL_6) begin
    if (_EVAL_6) begin
      _EVAL_10 <= 1'h0;
    end else if (_EVAL_31) begin
      if (_EVAL_37) begin
        _EVAL_10 <= 1'h0;
      end else begin
        _EVAL_10 <= _EVAL_18;
      end
    end
  end
  always @(posedge _EVAL_8 or posedge _EVAL_6) begin
    if (_EVAL_6) begin
      _EVAL_32 <= 32'h0;
    end else if (_EVAL_115) begin
      _EVAL_32 <= 32'h0;
    end else begin
      _EVAL_32 <= _EVAL_67;
    end
  end
  always @(posedge _EVAL_8 or posedge _EVAL_6) begin
    if (_EVAL_6) begin
      _EVAL_78 <= 1'h0;
    end else if (_EVAL_17) begin
      if (_EVAL_108) begin
        _EVAL_78 <= 1'h0;
      end else begin
        _EVAL_78 <= _EVAL_61;
      end
    end
  end
  always @(posedge _EVAL_8 or posedge _EVAL_6) begin
    if (_EVAL_6) begin
      _EVAL_80 <= 1'h0;
    end else if (_EVAL_17) begin
      if (_EVAL_43) begin
        _EVAL_80 <= 1'h0;
      end else begin
        _EVAL_80 <= _EVAL_34;
      end
    end
  end
  always @(posedge _EVAL_8 or posedge _EVAL_6) begin
    if (_EVAL_6) begin
      _EVAL_90 <= 1'h0;
    end else if (_EVAL_31) begin
      if (_EVAL_33) begin
        _EVAL_90 <= 1'h0;
      end else begin
        _EVAL_90 <= _EVAL_124;
      end
    end
  end
  always @(posedge _EVAL_8 or posedge _EVAL_6) begin
    if (_EVAL_6) begin
      _EVAL_109 <= 1'h0;
    end else begin
      _EVAL_109 <= _EVAL_55 & _EVAL_52;
    end
  end

endmodule
