//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_59(
  input  [31:0] _EVAL,
  input         _EVAL_0,
  output        _EVAL_1,
  output        _EVAL_2,
  input  [2:0]  _EVAL_3,
  output        _EVAL_4,
  output        _EVAL_5,
  input  [31:0] _EVAL_6,
  output [29:0] _EVAL_7,
  input  [2:0]  _EVAL_8,
  output        _EVAL_9,
  input         _EVAL_10,
  output [31:0] _EVAL_11,
  input         _EVAL_12,
  input  [3:0]  _EVAL_13,
  input         _EVAL_14,
  output        _EVAL_15,
  input  [29:0] _EVAL_16,
  output [3:0]  _EVAL_17,
  input         _EVAL_18,
  input  [3:0]  _EVAL_19,
  output [2:0]  _EVAL_20,
  output [3:0]  _EVAL_21,
  input  [2:0]  _EVAL_22,
  input         _EVAL_23,
  output [2:0]  _EVAL_24,
  output [1:0]  _EVAL_25,
  output        _EVAL_26,
  input  [2:0]  _EVAL_27,
  output [31:0] _EVAL_28,
  output        _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  input  [1:0]  _EVAL_33,
  output        _EVAL_34,
  output [3:0]  _EVAL_35,
  output        _EVAL_36,
  input         _EVAL_37,
  input  [3:0]  _EVAL_38,
  output [2:0]  _EVAL_39,
  input         _EVAL_40,
  input         _EVAL_41,
  input         _EVAL_42,
  output        _EVAL_43,
  input  [2:0]  _EVAL_44,
  output [2:0]  _EVAL_45,
  input         _EVAL_46,
  output        _EVAL_47,
  output [2:0]  _EVAL_48
);
  reg [2:0] _EVAL_49;
  reg [31:0] _RAND_0;
  wire [29:0] _EVAL_50;
  wire  _EVAL_52;
  wire [30:0] _EVAL_53;
  wire  _EVAL_55;
  wire [30:0] _EVAL_56;
  wire [22:0] _EVAL_61;
  wire [6:0] _EVAL_62;
  wire  _EVAL_66;
  wire [30:0] _EVAL_67;
  wire  _EVAL_68;
  reg  _EVAL_69;
  reg [31:0] _RAND_1;
  wire  _EVAL_72;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire [5:0] _EVAL_77;
  wire [29:0] _EVAL_79;
  wire [1:0] _EVAL_80;
  wire [30:0] _EVAL_81;
  wire  _EVAL_82;
  wire [1:0] _EVAL_83;
  wire  _EVAL_84;
  wire [7:0] _EVAL_85;
  wire [1:0] _EVAL_87;
  reg [5:0] _EVAL_89;
  reg [31:0] _RAND_2;
  wire [6:0] _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire [29:0] _EVAL_94;
  wire  _EVAL_96;
  wire [7:0] _EVAL_97;
  wire  _EVAL_100;
  wire [7:0] _EVAL_101;
  wire  _EVAL_102;
  wire [5:0] _EVAL_103;
  wire [30:0] _EVAL_105;
  wire [2:0] _EVAL_107;
  wire [5:0] _EVAL_110;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire [30:0] _EVAL_116;
  wire  _EVAL_118;
  wire [1:0] _EVAL_119;
  reg [5:0] _EVAL_120;
  reg [31:0] _RAND_3;
  wire [30:0] _EVAL_123;
  wire [7:0] _EVAL_124;
  wire [30:0] _EVAL_125;
  wire  _EVAL_127;
  wire [2:0] _EVAL_128;
  wire  _EVAL_129;
  wire [22:0] _EVAL_132;
  wire [30:0] _EVAL_134;
  wire [30:0] _EVAL_137;
  wire [1:0] _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire [30:0] _EVAL_141;
  wire  _EVAL_143;
  wire [2:0] _EVAL_145;
  wire [2:0] _EVAL_146;
  reg  _EVAL_148;
  reg [31:0] _RAND_4;
  wire [30:0] _EVAL_149;
  wire  _EVAL_151;
  wire [1:0] _EVAL_153;
  wire [30:0] _EVAL_154;
  wire [30:0] _EVAL_156;
  wire  _EVAL_157;
  wire [2:0] _EVAL_159;
  wire [5:0] _EVAL_160;
  wire [29:0] _EVAL_161;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire [30:0] _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  assign _EVAL_139 = _EVAL_3[2];
  assign _EVAL_129 = _EVAL_74 | _EVAL_143;
  assign _EVAL_110 = _EVAL_97[7:2];
  assign _EVAL_79 = _EVAL_16 ^ 30'h2000;
  assign _EVAL_157 = _EVAL_82 & _EVAL_129;
  assign _EVAL_163 = $signed(_EVAL_67) == 31'sh0;
  assign _EVAL_96 = _EVAL_75 & _EVAL_140;
  assign _EVAL_94 = _EVAL_16 ^ 30'h20000000;
  assign _EVAL_91 = _EVAL_120 - 6'h1;
  assign _EVAL_7 = _EVAL_16;
  assign _EVAL_93 = _EVAL_68 & _EVAL_75;
  assign _EVAL_35 = _EVAL_19;
  assign _EVAL_166 = {1'b0,$signed(_EVAL_50)};
  assign _EVAL_76 = _EVAL_115 | _EVAL_148;
  assign _EVAL_53 = $signed(_EVAL_137) & 31'sh22006000;
  assign _EVAL_159 = _EVAL_107 | _EVAL_128;
  assign _EVAL_62 = _EVAL_89 - 6'h1;
  assign _EVAL_83 = _EVAL_138 | _EVAL_87;
  assign _EVAL_107 = {{1'd0}, _EVAL_153};
  assign _EVAL_45 = _EVAL_44;
  assign _EVAL_102 = _EVAL_31 & _EVAL_40;
  assign _EVAL_20 = _EVAL_3;
  assign _EVAL_171 = 3'h0 == _EVAL_44;
  assign _EVAL_4 = _EVAL_32;
  assign _EVAL_56 = _EVAL_53;
  assign _EVAL_164 = _EVAL_72 & _EVAL_102;
  assign _EVAL_43 = _EVAL_0;
  assign _EVAL_85 = _EVAL_61[7:0];
  assign _EVAL_141 = {1'b0,$signed(_EVAL_161)};
  assign _EVAL_11 = _EVAL_6;
  assign _EVAL_105 = {1'b0,$signed(_EVAL_79)};
  assign _EVAL_61 = 23'hff << _EVAL_13;
  assign _EVAL_149 = _EVAL_156;
  assign _EVAL_132 = 23'hff << _EVAL_38;
  assign _EVAL_5 = _EVAL_14 & _EVAL_118;
  assign _EVAL_172 = $signed(_EVAL_149) == 31'sh0;
  assign _EVAL_75 = _EVAL_167 & _EVAL_30;
  assign _EVAL_74 = _EVAL_145 == 3'h0;
  assign _EVAL_167 = _EVAL_14 & _EVAL_118;
  assign _EVAL_100 = _EVAL_89 == 6'h0;
  assign _EVAL_145 = _EVAL_159 | _EVAL_146;
  assign _EVAL_55 = _EVAL_171 | _EVAL_69;
  assign _EVAL_127 = $signed(_EVAL_56) == 31'sh0;
  assign _EVAL_140 = _EVAL_80 == 2'h0;
  assign _EVAL_47 = _EVAL_10;
  assign _EVAL_173 = $signed(_EVAL_134) == 31'sh0;
  assign _EVAL_66 = _EVAL_8[0];
  assign _EVAL_21 = _EVAL_13;
  assign _EVAL_50 = _EVAL_16 ^ 30'h2000000;
  assign _EVAL_80 = _EVAL_44[2:1];
  assign _EVAL_67 = _EVAL_125;
  assign _EVAL_24 = _EVAL_22;
  assign _EVAL_2 = _EVAL_30 & _EVAL_118;
  assign _EVAL_116 = $signed(_EVAL_141) & 31'sh22006000;
  assign _EVAL_48 = _EVAL_8;
  assign _EVAL_29 = _EVAL_42;
  assign _EVAL_156 = $signed(_EVAL_105) & 31'sh22006000;
  assign _EVAL_17 = _EVAL_38;
  assign _EVAL_118 = ~_EVAL_157;
  assign _EVAL_146 = _EVAL_173 ? 3'h5 : 3'h0;
  assign _EVAL_115 = 3'h1 == _EVAL_44;
  assign _EVAL_87 = _EVAL_163 ? 2'h2 : 2'h0;
  assign _EVAL_77 = _EVAL_91[5:0];
  assign _EVAL_153 = _EVAL_83 | _EVAL_119;
  assign _EVAL_103 = _EVAL_101[7:2];
  assign _EVAL_151 = ~_EVAL_139;
  assign _EVAL_72 = _EVAL_100 & _EVAL_84;
  assign _EVAL_68 = _EVAL_120 == 6'h0;
  assign _EVAL_34 = _EVAL_41;
  assign _EVAL_143 = _EVAL_49 != _EVAL_145;
  assign _EVAL_123 = $signed(_EVAL_154) & 31'sh22006000;
  assign _EVAL_25 = _EVAL_33;
  assign _EVAL_52 = _EVAL_140 & _EVAL_68;
  assign _EVAL_119 = _EVAL_92 ? 2'h3 : 2'h0;
  assign _EVAL_28 = _EVAL;
  assign _EVAL_15 = _EVAL_31;
  assign _EVAL_97 = ~_EVAL_124;
  assign _EVAL_9 = _EVAL_40;
  assign _EVAL_124 = _EVAL_132[7:0];
  assign _EVAL_128 = _EVAL_127 ? 3'h4 : 3'h0;
  assign _EVAL_154 = {1'b0,$signed(_EVAL_16)};
  assign _EVAL_161 = _EVAL_16 ^ 30'h4000;
  assign _EVAL_81 = _EVAL_123;
  assign _EVAL_1 = _EVAL_46;
  assign _EVAL_137 = {1'b0,$signed(_EVAL_94)};
  assign _EVAL_39 = _EVAL_27;
  assign _EVAL_92 = $signed(_EVAL_81) == 31'sh0;
  assign _EVAL_82 = _EVAL_52 & _EVAL_114;
  assign _EVAL_84 = _EVAL_8 != 3'h6;
  assign _EVAL_26 = _EVAL_18;
  assign _EVAL_134 = _EVAL_116;
  assign _EVAL_160 = _EVAL_62[5:0];
  assign _EVAL_125 = $signed(_EVAL_166) & 31'sh22000000;
  assign _EVAL_114 = _EVAL_69 | _EVAL_148;
  assign _EVAL_138 = {{1'd0}, _EVAL_172};
  assign _EVAL_101 = ~_EVAL_85;
  assign _EVAL_36 = _EVAL_23;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_49 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_69 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_89 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_120 = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_148 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_12) begin
    if (_EVAL_96) begin
      _EVAL_49 <= _EVAL_145;
    end
    if (_EVAL_37) begin
      _EVAL_69 <= 1'h0;
    end else if (_EVAL_164) begin
      if (3'h0 == _EVAL_22) begin
        _EVAL_69 <= 1'h0;
      end else if (_EVAL_93) begin
        _EVAL_69 <= _EVAL_55;
      end
    end else if (_EVAL_93) begin
      _EVAL_69 <= _EVAL_55;
    end
    if (_EVAL_37) begin
      _EVAL_89 <= 6'h0;
    end else if (_EVAL_102) begin
      if (_EVAL_100) begin
        if (_EVAL_66) begin
          _EVAL_89 <= _EVAL_103;
        end else begin
          _EVAL_89 <= 6'h0;
        end
      end else begin
        _EVAL_89 <= _EVAL_160;
      end
    end
    if (_EVAL_37) begin
      _EVAL_120 <= 6'h0;
    end else if (_EVAL_75) begin
      if (_EVAL_68) begin
        if (_EVAL_151) begin
          _EVAL_120 <= _EVAL_110;
        end else begin
          _EVAL_120 <= 6'h0;
        end
      end else begin
        _EVAL_120 <= _EVAL_77;
      end
    end
    if (_EVAL_37) begin
      _EVAL_148 <= 1'h0;
    end else if (_EVAL_164) begin
      if (3'h1 == _EVAL_22) begin
        _EVAL_148 <= 1'h0;
      end else if (_EVAL_93) begin
        _EVAL_148 <= _EVAL_76;
      end
    end else if (_EVAL_93) begin
      _EVAL_148 <= _EVAL_76;
    end
  end
endmodule
