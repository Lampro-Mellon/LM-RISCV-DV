//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_15_assert(
  input  [3:0]  _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input  [1:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  input  [1:0]  _EVAL_11,
  input  [31:0] _EVAL_12,
  input  [2:0]  _EVAL_13,
  input         _EVAL_14
);
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire [31:0] _EVAL_26;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  reg [31:0] _EVAL_31;
  reg [31:0] _RAND_0;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire [4:0] _EVAL_36;
  wire  _EVAL_37;
  wire [1:0] _EVAL_38;
  wire [1:0] _EVAL_39;
  wire  _EVAL_40;
  wire [3:0] _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire [7:0] _EVAL_44;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire [3:0] _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire [32:0] _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  reg  _EVAL_66;
  reg [31:0] _RAND_1;
  wire  _EVAL_67;
  wire [32:0] _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_71;
  wire [32:0] _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire [7:0] _EVAL_77;
  wire [3:0] _EVAL_78;
  wire  _EVAL_79;
  wire [1:0] _EVAL_80;
  wire [4:0] _EVAL_81;
  reg [1:0] _EVAL_82;
  reg [31:0] _RAND_2;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire [4:0] _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  reg [2:0] _EVAL_99;
  reg [31:0] _RAND_3;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire [7:0] _EVAL_106;
  wire  _EVAL_107;
  wire [31:0] _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  reg  _EVAL_111;
  reg [31:0] _RAND_4;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire [1:0] _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire [4:0] _EVAL_129;
  wire  _EVAL_130;
  wire [1:0] _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire [1:0] _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire [4:0] _EVAL_148;
  wire  _EVAL_149;
  reg  _EVAL_150;
  reg [31:0] _RAND_5;
  wire [32:0] _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire [4:0] _EVAL_167;
  reg [2:0] _EVAL_168;
  reg [31:0] _RAND_6;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire [4:0] _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  reg [2:0] _EVAL_174;
  reg [31:0] _RAND_7;
  wire [4:0] _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  reg [1:0] _EVAL_179;
  reg [31:0] _RAND_8;
  wire [7:0] _EVAL_180;
  wire  _EVAL_181;
  wire [1:0] _EVAL_182;
  wire [1:0] _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire [4:0] _EVAL_186;
  wire  _EVAL_187;
  wire [3:0] _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  reg [2:0] _EVAL_195;
  reg [31:0] _RAND_9;
  wire [1:0] _EVAL_196;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  reg [4:0] _EVAL_205;
  reg [31:0] _RAND_10;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire [31:0] _EVAL_215;
  wire  _EVAL_216;
  reg  _EVAL_217;
  reg [31:0] _RAND_11;
  wire  _EVAL_218;
  wire [31:0] _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_222;
  wire [1:0] _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  reg [2:0] _EVAL_234;
  reg [31:0] _RAND_12;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  reg [31:0] _EVAL_246;
  reg [31:0] _RAND_13;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_98 = _EVAL_207 & _EVAL_209;
  assign _EVAL_186 = _EVAL_205 >> _EVAL_9;
  assign _EVAL_78 = _EVAL & _EVAL_51;
  assign _EVAL_149 = ~_EVAL_237;
  assign _EVAL_105 = ~_EVAL_18;
  assign _EVAL_250 = ~_EVAL_111;
  assign _EVAL_236 = _EVAL_42 | _EVAL_14;
  assign _EVAL_35 = ~_EVAL_136;
  assign _EVAL_144 = _EVAL_129[0];
  assign _EVAL_165 = _EVAL_102 | _EVAL_14;
  assign _EVAL_141 = _EVAL_187 | _EVAL_14;
  assign _EVAL_21 = _EVAL_157 | _EVAL_58;
  assign _EVAL_48 = _EVAL_144 | _EVAL_14;
  assign _EVAL_202 = _EVAL_1 != 3'h0;
  assign _EVAL_145 = _EVAL_113 | _EVAL_14;
  assign _EVAL_18 = _EVAL_133 | _EVAL_14;
  assign _EVAL_72 = _EVAL_246 + 32'h1;
  assign _EVAL_64 = ~_EVAL_66;
  assign _EVAL_97 = _EVAL_125 | _EVAL_225;
  assign _EVAL_79 = _EVAL_1 <= 3'h2;
  assign _EVAL_189 = _EVAL_13 == 3'h4;
  assign _EVAL_67 = _EVAL_43 & _EVAL_49;
  assign _EVAL_192 = _EVAL_87 | _EVAL_14;
  assign _EVAL_120 = _EVAL_86 != _EVAL_36;
  assign _EVAL_143 = _EVAL_118 | _EVAL_14;
  assign _EVAL_107 = _EVAL_223[0];
  assign _EVAL_183 = 2'h1 << _EVAL_238;
  assign _EVAL_54 = _EVAL_56 | _EVAL_14;
  assign _EVAL_170 = ~_EVAL_64;
  assign _EVAL_108 = {{30'd0}, _EVAL_196};
  assign _EVAL_244 = _EVAL_10 & _EVAL_247;
  assign _EVAL_228 = ~_EVAL_141;
  assign _EVAL_29 = _EVAL_10 & _EVAL_229;
  assign _EVAL_235 = _EVAL_2 == 3'h6;
  assign _EVAL_32 = ~_EVAL_150;
  assign _EVAL_51 = ~_EVAL_188;
  assign _EVAL_84 = ~_EVAL_242;
  assign _EVAL_215 = _EVAL_72[31:0];
  assign _EVAL_225 = _EVAL_207 & _EVAL_181;
  assign _EVAL_25 = _EVAL_11 <= 2'h2;
  assign _EVAL_172 = _EVAL_139 | _EVAL_14;
  assign _EVAL_241 = _EVAL_39[0];
  assign _EVAL_185 = _EVAL_202 | _EVAL_14;
  assign _EVAL_220 = _EVAL_13 == 3'h2;
  assign _EVAL_237 = _EVAL_12[1];
  assign _EVAL_94 = _EVAL_5 & _EVAL_6;
  assign _EVAL_34 = ~_EVAL_32;
  assign _EVAL_131 = _EVAL_4[2:1];
  assign _EVAL_60 = _EVAL_153 & _EVAL_149;
  assign _EVAL_198 = _EVAL_10 & _EVAL_189;
  assign _EVAL_53 = _EVAL_12 == _EVAL_31;
  assign _EVAL_47 = _EVAL_10 & _EVAL_100;
  assign _EVAL_223 = _EVAL_217 - 1'h1;
  assign _EVAL_122 = _EVAL_30 | _EVAL_134;
  assign _EVAL_188 = {_EVAL_138,_EVAL_243,_EVAL_224,_EVAL_97};
  assign _EVAL_57 = $signed(_EVAL_68) & -33'sh4000;
  assign _EVAL_91 = ~_EVAL_16;
  assign _EVAL_129 = _EVAL_81 >> _EVAL_4;
  assign _EVAL_134 = _EVAL_9 == 3'h4;
  assign _EVAL_151 = _EVAL_57;
  assign _EVAL_59 = _EVAL_201 | _EVAL_14;
  assign _EVAL_103 = ~_EVAL_83;
  assign _EVAL_136 = _EVAL_191 | _EVAL_14;
  assign _EVAL_227 = _EVAL_79 | _EVAL_14;
  assign _EVAL_104 = _EVAL_2 == 3'h2;
  assign _EVAL_22 = _EVAL_73 | _EVAL_14;
  assign _EVAL_87 = _EVAL_8 >= 2'h2;
  assign _EVAL_208 = _EVAL_131 == 2'h0;
  assign _EVAL_92 = _EVAL_13 == 3'h0;
  assign _EVAL_247 = _EVAL_13 == 3'h3;
  assign _EVAL_240 = _EVAL_4 == _EVAL_234;
  assign _EVAL_95 = ~_EVAL_192;
  assign _EVAL_155 = _EVAL_37 | _EVAL_69;
  assign _EVAL_52 = _EVAL_162 | _EVAL_14;
  assign _EVAL_68 = {1'b0,$signed(_EVAL_26)};
  assign _EVAL_238 = _EVAL_11[0];
  assign _EVAL_156 = _EVAL_12[0];
  assign _EVAL_102 = _EVAL_13 == _EVAL_99;
  assign _EVAL_137 = _EVAL_117 | _EVAL_14;
  assign _EVAL_114 = ~_EVAL_71;
  assign _EVAL_201 = ~_EVAL_3;
  assign _EVAL_177 = _EVAL_182 == 2'h0;
  assign _EVAL_222 = _EVAL_153 & _EVAL_237;
  assign _EVAL_138 = _EVAL_128 | _EVAL_50;
  assign _EVAL_39 = _EVAL_66 - 1'h1;
  assign _EVAL_26 = _EVAL_12 ^ 32'h80008000;
  assign _EVAL_173 = _EVAL_21 | _EVAL_14;
  assign _EVAL_133 = _EVAL_1 <= 3'h4;
  assign _EVAL_212 = ~_EVAL_173;
  assign _EVAL_46 = ~_EVAL_185;
  assign _EVAL_216 = _EVAL_1 == _EVAL_174;
  assign _EVAL_126 = _EVAL_155 | _EVAL_14;
  assign _EVAL_162 = _EVAL_78 == 4'h0;
  assign _EVAL_230 = ~_EVAL_248;
  assign _EVAL_243 = _EVAL_128 | _EVAL_98;
  assign _EVAL_153 = _EVAL_38[1];
  assign _EVAL_81 = _EVAL_86 | _EVAL_205;
  assign _EVAL_239 = ~_EVAL_14;
  assign _EVAL_83 = _EVAL_154 | _EVAL_14;
  assign _EVAL_164 = _EVAL_6 & _EVAL_55;
  assign _EVAL_37 = _EVAL_251 | _EVAL_33;
  assign _EVAL_17 = _EVAL_6 & _EVAL_235;
  assign _EVAL_16 = _EVAL_122 | _EVAL_14;
  assign _EVAL_203 = ~_EVAL_190;
  assign _EVAL_63 = _EVAL_123 | _EVAL_14;
  assign _EVAL_100 = _EVAL_13 == 3'h1;
  assign _EVAL_213 = _EVAL_6 & _EVAL_184;
  assign _EVAL_194 = _EVAL_10 & _EVAL_92;
  assign _EVAL_214 = ~_EVAL_63;
  assign _EVAL_36 = _EVAL_106[4:0];
  assign _EVAL_58 = _EVAL_4 == 3'h4;
  assign _EVAL_207 = _EVAL_38[0];
  assign _EVAL_210 = ~_EVAL_48;
  assign _EVAL_113 = _EVAL_41 == 4'h0;
  assign _EVAL_77 = 8'h1 << _EVAL_9;
  assign _EVAL_28 = _EVAL_193 & _EVAL_32;
  assign _EVAL_44 = 8'h1 << _EVAL_4;
  assign _EVAL_33 = plusarg_reader_out == 32'h0;
  assign _EVAL_132 = _EVAL_124[0];
  assign _EVAL_115 = _EVAL_13 == 3'h6;
  assign _EVAL_121 = _EVAL_76 | _EVAL_14;
  assign _EVAL_50 = _EVAL_207 & _EVAL_130;
  assign _EVAL_89 = _EVAL_6 & _EVAL_104;
  assign _EVAL_146 = ~_EVAL_137;
  assign _EVAL_148 = _EVAL_167 & _EVAL_175;
  assign _EVAL_181 = _EVAL_149 & _EVAL_218;
  assign _EVAL_211 = _EVAL_140[0];
  assign _EVAL_184 = _EVAL_2 == 3'h0;
  assign _EVAL_248 = _EVAL_88 | _EVAL_14;
  assign _EVAL_157 = _EVAL_200 | _EVAL_208;
  assign _EVAL_245 = ~_EVAL_145;
  assign _EVAL_55 = _EVAL_2 == 3'h5;
  assign _EVAL_231 = _EVAL_186[0];
  assign _EVAL_69 = _EVAL_246 < plusarg_reader_out;
  assign _EVAL_118 = _EVAL_1 == 3'h0;
  assign _EVAL_43 = _EVAL_94 & _EVAL_20;
  assign _EVAL_171 = 5'h3 << _EVAL_11;
  assign _EVAL_130 = _EVAL_237 & _EVAL_156;
  assign _EVAL_176 = _EVAL_10 & _EVAL_34;
  assign _EVAL_249 = ~_EVAL_121;
  assign _EVAL_147 = _EVAL_10 & _EVAL_220;
  assign _EVAL_233 = _EVAL_149 & _EVAL_156;
  assign _EVAL_242 = _EVAL_216 | _EVAL_14;
  assign _EVAL_200 = _EVAL_131 == 2'h1;
  assign _EVAL_154 = _EVAL_219 == 32'h0;
  assign _EVAL_251 = ~_EVAL_116;
  assign _EVAL_128 = _EVAL_73 | _EVAL_222;
  assign _EVAL_125 = _EVAL_73 | _EVAL_60;
  assign _EVAL_163 = _EVAL_86 != 5'h0;
  assign _EVAL_71 = _EVAL_53 | _EVAL_14;
  assign _EVAL_38 = _EVAL_183 | 2'h1;
  assign _EVAL_139 = _EVAL_1 <= 3'h1;
  assign _EVAL_40 = _EVAL_10 & _EVAL_115;
  assign _EVAL_187 = _EVAL_9 == _EVAL_195;
  assign _EVAL_61 = _EVAL_2 == 3'h1;
  assign _EVAL_49 = ~_EVAL_235;
  assign _EVAL_166 = ~_EVAL_172;
  assign _EVAL_191 = ~_EVAL_231;
  assign _EVAL_80 = _EVAL_171[1:0];
  assign _EVAL_119 = ~_EVAL_236;
  assign _EVAL_219 = _EVAL_12 & _EVAL_108;
  assign _EVAL_23 = ~_EVAL_22;
  assign _EVAL_62 = ~_EVAL_160;
  assign _EVAL_175 = ~_EVAL_36;
  assign _EVAL_209 = _EVAL_237 & _EVAL_218;
  assign _EVAL_199 = ~_EVAL_52;
  assign _EVAL_109 = ~_EVAL_163;
  assign _EVAL_224 = _EVAL_125 | _EVAL_161;
  assign _EVAL_93 = _EVAL_2 <= 3'h6;
  assign _EVAL_167 = _EVAL_205 | _EVAL_86;
  assign _EVAL_124 = _EVAL_111 - 1'h1;
  assign _EVAL_182 = _EVAL_9[2:1];
  assign _EVAL_85 = _EVAL_240 | _EVAL_14;
  assign _EVAL_135 = _EVAL_94 & _EVAL_64;
  assign _EVAL_232 = ~_EVAL_59;
  assign _EVAL_152 = _EVAL_1 <= 3'h3;
  assign _EVAL_75 = ~_EVAL_126;
  assign _EVAL_42 = _EVAL_11 == _EVAL_82;
  assign _EVAL_110 = _EVAL_6 & _EVAL_170;
  assign _EVAL_160 = _EVAL_152 | _EVAL_14;
  assign _EVAL_90 = ~_EVAL_54;
  assign _EVAL_101 = _EVAL_13 == 3'h7;
  assign _EVAL_117 = _EVAL_120 | _EVAL_109;
  assign _EVAL_229 = _EVAL_13 == 3'h5;
  assign _EVAL_73 = _EVAL_11 >= 2'h2;
  assign _EVAL_159 = ~_EVAL_165;
  assign _EVAL_30 = _EVAL_112 | _EVAL_177;
  assign _EVAL_193 = _EVAL_0 & _EVAL_10;
  assign _EVAL_106 = _EVAL_67 ? _EVAL_44 : 8'h0;
  assign _EVAL_196 = ~_EVAL_80;
  assign _EVAL_158 = _EVAL_2 == 3'h4;
  assign _EVAL_178 = ~_EVAL_227;
  assign _EVAL_169 = $signed(_EVAL_151) == 33'sh0;
  assign _EVAL_27 = ~_EVAL_85;
  assign _EVAL_96 = ~_EVAL_143;
  assign _EVAL_86 = _EVAL_180[4:0];
  assign _EVAL_20 = ~_EVAL_217;
  assign _EVAL_180 = _EVAL_19 ? _EVAL_77 : 8'h0;
  assign _EVAL_24 = _EVAL_10 & _EVAL_101;
  assign _EVAL_19 = _EVAL_193 & _EVAL_250;
  assign _EVAL_76 = _EVAL_25 & _EVAL_169;
  assign _EVAL_140 = _EVAL_150 - 1'h1;
  assign _EVAL_88 = _EVAL == _EVAL_188;
  assign _EVAL_123 = _EVAL_8 == _EVAL_179;
  assign _EVAL_218 = ~_EVAL_156;
  assign _EVAL_56 = _EVAL_2 == _EVAL_168;
  assign _EVAL_41 = ~_EVAL;
  assign _EVAL_74 = _EVAL_6 & _EVAL_61;
  assign _EVAL_142 = _EVAL_193 | _EVAL_94;
  assign _EVAL_161 = _EVAL_207 & _EVAL_233;
  assign _EVAL_190 = _EVAL_93 | _EVAL_14;
  assign _EVAL_112 = _EVAL_182 == 2'h1;
  assign _EVAL_127 = _EVAL_6 & _EVAL_158;
  assign _EVAL_116 = _EVAL_205 != 5'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_31 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_66 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_82 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_99 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_111 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_150 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_168 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_174 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_179 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_195 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_205 = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_217 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_234 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_246 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_7) begin
    if (_EVAL_28) begin
      _EVAL_31 <= _EVAL_12;
    end
    if (_EVAL_14) begin
      _EVAL_66 <= 1'h0;
    end else if (_EVAL_94) begin
      if (_EVAL_64) begin
        _EVAL_66 <= 1'h0;
      end else begin
        _EVAL_66 <= _EVAL_241;
      end
    end
    if (_EVAL_28) begin
      _EVAL_82 <= _EVAL_11;
    end
    if (_EVAL_28) begin
      _EVAL_99 <= _EVAL_13;
    end
    if (_EVAL_14) begin
      _EVAL_111 <= 1'h0;
    end else if (_EVAL_193) begin
      if (_EVAL_250) begin
        _EVAL_111 <= 1'h0;
      end else begin
        _EVAL_111 <= _EVAL_132;
      end
    end
    if (_EVAL_14) begin
      _EVAL_150 <= 1'h0;
    end else if (_EVAL_193) begin
      if (_EVAL_32) begin
        _EVAL_150 <= 1'h0;
      end else begin
        _EVAL_150 <= _EVAL_211;
      end
    end
    if (_EVAL_135) begin
      _EVAL_168 <= _EVAL_2;
    end
    if (_EVAL_28) begin
      _EVAL_174 <= _EVAL_1;
    end
    if (_EVAL_135) begin
      _EVAL_179 <= _EVAL_8;
    end
    if (_EVAL_28) begin
      _EVAL_195 <= _EVAL_9;
    end
    if (_EVAL_14) begin
      _EVAL_205 <= 5'h0;
    end else begin
      _EVAL_205 <= _EVAL_148;
    end
    if (_EVAL_14) begin
      _EVAL_217 <= 1'h0;
    end else if (_EVAL_94) begin
      if (_EVAL_20) begin
        _EVAL_217 <= 1'h0;
      end else begin
        _EVAL_217 <= _EVAL_107;
      end
    end
    if (_EVAL_135) begin
      _EVAL_234 <= _EVAL_4;
    end
    if (_EVAL_14) begin
      _EVAL_246 <= 32'h0;
    end else if (_EVAL_142) begin
      _EVAL_246 <= 32'h0;
    end else begin
      _EVAL_246 <= _EVAL_215;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d6912ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12cc085b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b5df1bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5da7ef03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(153b1d4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9ed589f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac9897ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9988054)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(681ced20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d932328)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(374eebc4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dae890)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b834302)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e81f766)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5995e33a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16bff2e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa9e2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8dc7c40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b85bdbe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79006157)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23b28419)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5abbf67f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70edda43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76a394d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c1c5b0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f8bcea4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f833ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c32dce8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8755312)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e5d2ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d655cd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63776fde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16e918cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe690c5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e469f1a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(357d37b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7089ee8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0e69d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3071c1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(128eb754)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a022c37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49322553)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59ab7528)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ddedf4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0a3e71f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(816d070)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fbf5250)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3545268b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42a75fa5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bf74c3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e46ab81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a324cab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(383e8c3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(920a12ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c850b028)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91fad6d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6720869)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51dafc58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92dc7fd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d2213a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59308c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bea80ca1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f97f2b2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61e3459)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b776e5ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc3c38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce733cec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55b53f2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(865cbda4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8205fd9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd5830fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9d22644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d42b41e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
