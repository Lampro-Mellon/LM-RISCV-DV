//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_86_assert(
  input         _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [1:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [1:0]  _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input  [2:0]  _EVAL_8,
  input         _EVAL_9,
  input  [1:0]  _EVAL_10,
  input  [3:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [2:0]  _EVAL_13,
  input  [29:0] _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18
);
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire [29:0] _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire [4:0] _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire [30:0] _EVAL_34;
  wire  _EVAL_35;
  wire [1:0] _EVAL_36;
  wire [1:0] _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire [29:0] _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  reg  _EVAL_47;
  reg [31:0] _RAND_0;
  wire  _EVAL_48;
  wire [3:0] _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire [7:0] _EVAL_53;
  wire  _EVAL_54;
  wire [1:0] _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire [4:0] _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  reg  _EVAL_62;
  reg [31:0] _RAND_1;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  reg [29:0] _EVAL_71;
  reg [31:0] _RAND_2;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  reg [2:0] _EVAL_75;
  reg [31:0] _RAND_3;
  reg [1:0] _EVAL_76;
  reg [31:0] _RAND_4;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire [4:0] _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire [31:0] _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_89;
  wire [30:0] _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  reg [2:0] _EVAL_98;
  reg [31:0] _RAND_5;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire [3:0] _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire [4:0] _EVAL_106;
  wire  _EVAL_107;
  wire [29:0] _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  reg [31:0] _EVAL_116;
  reg [31:0] _RAND_6;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire [1:0] _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire [7:0] _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  reg [1:0] _EVAL_138;
  reg [31:0] _RAND_7;
  wire [7:0] _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire [4:0] _EVAL_145;
  wire [3:0] _EVAL_146;
  reg [1:0] _EVAL_147;
  reg [31:0] _RAND_8;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire [4:0] _EVAL_150;
  reg  _EVAL_151;
  reg [31:0] _RAND_9;
  reg [4:0] _EVAL_152;
  reg [31:0] _RAND_10;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire [30:0] _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire [7:0] _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  reg  _EVAL_175;
  reg [31:0] _RAND_11;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire [1:0] _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  reg [2:0] _EVAL_211;
  reg [31:0] _RAND_12;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire [4:0] _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire [4:0] _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire [1:0] _EVAL_233;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  reg [2:0] _EVAL_241;
  reg [31:0] _RAND_13;
  wire  _EVAL_242;
  reg  _EVAL_243;
  reg [31:0] _RAND_14;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire [1:0] _EVAL_247;
  wire [32:0] _EVAL_248;
  wire  _EVAL_249;
  wire [3:0] _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire [4:0] _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire [1:0] _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  reg [2:0] _EVAL_268;
  reg [31:0] _RAND_15;
  wire  _EVAL_270;
  wire  _EVAL_271;
  reg  _EVAL_272;
  reg [31:0] _RAND_16;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_163 = ~_EVAL_6;
  assign _EVAL_40 = _EVAL_14 ^ 30'h20000000;
  assign _EVAL_162 = _EVAL_68 & _EVAL_230;
  assign _EVAL_215 = ~_EVAL_83;
  assign _EVAL_37 = _EVAL_175 - 1'h1;
  assign _EVAL_59 = ~_EVAL_106;
  assign _EVAL_251 = _EVAL_8 <= 3'h3;
  assign _EVAL_132 = 8'h1 << _EVAL_1;
  assign _EVAL_94 = ~_EVAL_104;
  assign _EVAL_213 = _EVAL_12 == 3'h4;
  assign _EVAL_134 = ~_EVAL_35;
  assign _EVAL_38 = _EVAL_250 == 4'h0;
  assign _EVAL_232 = _EVAL_93 | _EVAL_17;
  assign _EVAL_74 = _EVAL_200 | _EVAL_113;
  assign _EVAL_42 = _EVAL_67 | _EVAL_17;
  assign _EVAL_237 = _EVAL_15 == 3'h4;
  assign _EVAL_224 = _EVAL_21 | _EVAL_17;
  assign _EVAL_205 = ~_EVAL_201;
  assign _EVAL_253 = _EVAL_8 == _EVAL_241;
  assign _EVAL_91 = _EVAL_0 & _EVAL_263;
  assign _EVAL_227 = 5'h3 << _EVAL_10;
  assign _EVAL_72 = ~_EVAL_50;
  assign _EVAL_240 = _EVAL_4 & _EVAL;
  assign _EVAL_63 = ~_EVAL_232;
  assign _EVAL_129 = _EVAL & _EVAL_105;
  assign _EVAL_117 = _EVAL & _EVAL_137;
  assign _EVAL_84 = $signed(_EVAL_157) == 31'sh0;
  assign _EVAL_201 = _EVAL_20 | _EVAL_17;
  assign _EVAL_257 = _EVAL_153 & _EVAL_270;
  assign _EVAL_107 = _EVAL_130 | _EVAL_17;
  assign _EVAL_185 = ~_EVAL_36;
  assign _EVAL_124 = _EVAL_253 | _EVAL_17;
  assign _EVAL_85 = _EVAL_2 != 2'h2;
  assign _EVAL_226 = _EVAL_189 | _EVAL_17;
  assign _EVAL_208 = _EVAL_116 < plusarg_reader_out;
  assign _EVAL_122 = _EVAL_0 & _EVAL_236;
  assign _EVAL_118 = ~_EVAL_96;
  assign _EVAL_119 = ~_EVAL_17;
  assign _EVAL_190 = _EVAL_233[0];
  assign _EVAL_146 = _EVAL_11 & _EVAL_49;
  assign _EVAL_275 = _EVAL_77 | _EVAL_174;
  assign _EVAL_19 = _EVAL_14 == _EVAL_71;
  assign _EVAL_230 = ~_EVAL_260;
  assign _EVAL_102 = {_EVAL_275,_EVAL_159,_EVAL_74,_EVAL_186};
  assign _EVAL_206 = _EVAL_15 == 3'h1;
  assign _EVAL_267 = _EVAL_60 & _EVAL_142;
  assign _EVAL_133 = _EVAL_19 | _EVAL_17;
  assign _EVAL_194 = _EVAL_204 | _EVAL_17;
  assign _EVAL_34 = $signed(_EVAL_90) & -31'sh2000;
  assign _EVAL_168 = _EVAL_131 | _EVAL_17;
  assign _EVAL_171 = _EVAL_207 & _EVAL_199;
  assign _EVAL_172 = ~_EVAL_73;
  assign _EVAL_179 = _EVAL_38 | _EVAL_17;
  assign _EVAL_61 = _EVAL_39 | _EVAL_17;
  assign _EVAL_144 = _EVAL_0 & _EVAL_156;
  assign _EVAL_219 = ~_EVAL_168;
  assign _EVAL_31 = _EVAL_53[4:0];
  assign _EVAL_259 = _EVAL_150 & _EVAL_59;
  assign _EVAL_45 = _EVAL_68 & _EVAL_260;
  assign _EVAL_157 = _EVAL_34;
  assign _EVAL_89 = _EVAL_10 >= 2'h2;
  assign _EVAL_21 = _EVAL_12 == _EVAL_211;
  assign _EVAL_180 = _EVAL_8 <= 3'h2;
  assign _EVAL_109 = _EVAL & _EVAL_51;
  assign _EVAL_112 = ~_EVAL_178;
  assign _EVAL_78 = _EVAL_0 & _EVAL_57;
  assign _EVAL_93 = ~_EVAL_64;
  assign _EVAL_167 = _EVAL_240 & _EVAL_23;
  assign _EVAL_221 = _EVAL_196 | _EVAL_17;
  assign _EVAL_223 = ~_EVAL_160;
  assign _EVAL_49 = ~_EVAL_102;
  assign _EVAL_256 = ~_EVAL_225;
  assign _EVAL_181 = _EVAL_3 == _EVAL_272;
  assign _EVAL_27 = _EVAL_169 | _EVAL_208;
  assign _EVAL_145 = _EVAL_216 >> _EVAL_13;
  assign _EVAL_239 = _EVAL_153 & _EVAL_162;
  assign _EVAL_198 = _EVAL_222 | _EVAL_17;
  assign _EVAL_77 = _EVAL_89 | _EVAL_171;
  assign _EVAL_233 = _EVAL_47 - 1'h1;
  assign _EVAL_103 = ~_EVAL_133;
  assign _EVAL_46 = _EVAL_2 == _EVAL_147;
  assign _EVAL_218 = _EVAL_37[0];
  assign _EVAL_191 = _EVAL_15 == 3'h0;
  assign _EVAL_70 = ~_EVAL_69;
  assign _EVAL_41 = ~_EVAL_179;
  assign _EVAL_36 = _EVAL_227[1:0];
  assign _EVAL_123 = _EVAL_48 | _EVAL_17;
  assign _EVAL_255 = _EVAL_115 | _EVAL_17;
  assign _EVAL_197 = _EVAL & _EVAL_237;
  assign _EVAL_170 = _EVAL_148 | _EVAL_17;
  assign _EVAL_207 = _EVAL_55[1];
  assign _EVAL_225 = _EVAL_273 | _EVAL_17;
  assign _EVAL_100 = _EVAL_252 | _EVAL_17;
  assign _EVAL_158 = ~_EVAL_224;
  assign _EVAL_115 = _EVAL_8 <= 3'h4;
  assign _EVAL_80 = _EVAL_60 & _EVAL_149;
  assign _EVAL_33 = _EVAL_12 == 3'h2;
  assign _EVAL_81 = _EVAL_152 >> _EVAL_1;
  assign _EVAL_178 = _EVAL_181 | _EVAL_17;
  assign _EVAL_264 = _EVAL_29 | _EVAL_17;
  assign _EVAL_86 = _EVAL_248[31:0];
  assign _EVAL_128 = ~_EVAL_22;
  assign _EVAL_50 = _EVAL_180 | _EVAL_17;
  assign _EVAL_231 = ~_EVAL_264;
  assign _EVAL_187 = _EVAL_15 == 3'h7;
  assign _EVAL_99 = ~_EVAL_87;
  assign _EVAL_214 = ~_EVAL_54;
  assign _EVAL_30 = _EVAL_18 == _EVAL_151;
  assign _EVAL_54 = _EVAL_182 | _EVAL_17;
  assign _EVAL_209 = ~_EVAL_16;
  assign _EVAL_203 = _EVAL_0 & _EVAL_213;
  assign _EVAL_228 = _EVAL_207 & _EVAL_68;
  assign _EVAL_258 = ~_EVAL_198;
  assign _EVAL_48 = _EVAL_173 | _EVAL_261;
  assign _EVAL_184 = _EVAL_145[0];
  assign _EVAL_176 = ~_EVAL_65;
  assign _EVAL_101 = ~_EVAL_236;
  assign _EVAL_265 = 2'h1 << _EVAL_82;
  assign _EVAL_137 = _EVAL_15 == 3'h6;
  assign _EVAL_270 = _EVAL_199 & _EVAL_230;
  assign _EVAL_273 = _EVAL_10 == _EVAL_138;
  assign _EVAL_126 = ~_EVAL_243;
  assign _EVAL_236 = _EVAL_12 == 3'h6;
  assign _EVAL_79 = _EVAL & _EVAL_188;
  assign _EVAL_153 = _EVAL_55[0];
  assign _EVAL_90 = {1'b0,$signed(_EVAL_40)};
  assign _EVAL_58 = ~_EVAL_42;
  assign _EVAL_35 = _EVAL_85 | _EVAL_17;
  assign _EVAL_166 = ~_EVAL_123;
  assign _EVAL_177 = _EVAL_247[0];
  assign _EVAL_96 = _EVAL_32 | _EVAL_17;
  assign _EVAL_217 = _EVAL_13 <= 3'h4;
  assign _EVAL_200 = _EVAL_89 | _EVAL_228;
  assign _EVAL_113 = _EVAL_153 & _EVAL_45;
  assign _EVAL_55 = _EVAL_265 | 2'h1;
  assign _EVAL_92 = _EVAL_1 == _EVAL_75;
  assign _EVAL_183 = _EVAL_89 | _EVAL_17;
  assign _EVAL_229 = _EVAL_240 | _EVAL_60;
  assign _EVAL_182 = _EVAL_24 == 30'h0;
  assign _EVAL_66 = ~_EVAL_212;
  assign _EVAL_247 = _EVAL_243 - 1'h1;
  assign _EVAL_140 = ~_EVAL_44;
  assign _EVAL_136 = ~_EVAL_61;
  assign _EVAL_24 = _EVAL_14 & _EVAL_108;
  assign _EVAL_68 = ~_EVAL_199;
  assign _EVAL_216 = _EVAL_31 | _EVAL_152;
  assign _EVAL_261 = ~_EVAL_271;
  assign _EVAL_149 = ~_EVAL_175;
  assign _EVAL_114 = _EVAL_199 & _EVAL_260;
  assign _EVAL_212 = _EVAL_152 != 5'h0;
  assign _EVAL_22 = _EVAL_217 | _EVAL_17;
  assign _EVAL_202 = ~_EVAL_170;
  assign _EVAL_164 = _EVAL & _EVAL_187;
  assign _EVAL_87 = _EVAL_251 | _EVAL_17;
  assign _EVAL_195 = _EVAL_240 & _EVAL_126;
  assign _EVAL_53 = _EVAL_167 ? _EVAL_132 : 8'h0;
  assign _EVAL_169 = _EVAL_66 | _EVAL_266;
  assign _EVAL_156 = ~_EVAL_142;
  assign _EVAL_26 = _EVAL_13 == _EVAL_268;
  assign _EVAL_60 = _EVAL_9 & _EVAL_0;
  assign _EVAL_173 = _EVAL_31 != _EVAL_106;
  assign _EVAL_271 = _EVAL_31 != 5'h0;
  assign _EVAL_135 = _EVAL_0 & _EVAL_161;
  assign _EVAL_220 = _EVAL_154 & _EVAL_84;
  assign _EVAL_248 = _EVAL_116 + 32'h1;
  assign _EVAL_188 = _EVAL_15 == 3'h5;
  assign _EVAL_165 = 8'h1 << _EVAL_13;
  assign _EVAL_125 = _EVAL & _EVAL_191;
  assign _EVAL_244 = ~_EVAL_210;
  assign _EVAL_174 = _EVAL_153 & _EVAL_114;
  assign _EVAL_254 = ~_EVAL_194;
  assign _EVAL_196 = _EVAL_5 >= 2'h2;
  assign _EVAL_121 = _EVAL_127[0];
  assign _EVAL_23 = ~_EVAL_47;
  assign _EVAL_106 = _EVAL_139[4:0];
  assign _EVAL_238 = ~_EVAL_126;
  assign _EVAL_155 = ~_EVAL_107;
  assign _EVAL_143 = ~_EVAL_100;
  assign _EVAL_150 = _EVAL_152 | _EVAL_31;
  assign _EVAL_32 = _EVAL_11 == _EVAL_102;
  assign _EVAL_245 = ~_EVAL_226;
  assign _EVAL_250 = ~_EVAL_11;
  assign _EVAL_142 = ~_EVAL_62;
  assign _EVAL_39 = ~_EVAL_18;
  assign _EVAL_95 = ~_EVAL_124;
  assign _EVAL_44 = _EVAL_163 | _EVAL_17;
  assign _EVAL_82 = _EVAL_10[0];
  assign _EVAL_28 = ~_EVAL_221;
  assign _EVAL_64 = _EVAL_81[0];
  assign _EVAL_105 = _EVAL_15 == 3'h3;
  assign _EVAL_186 = _EVAL_200 | _EVAL_239;
  assign _EVAL_148 = _EVAL_8 != 3'h0;
  assign _EVAL_204 = _EVAL_8 <= 3'h1;
  assign _EVAL_25 = _EVAL_184 | _EVAL_17;
  assign _EVAL_127 = _EVAL_62 - 1'h1;
  assign _EVAL_274 = _EVAL_46 | _EVAL_17;
  assign _EVAL_161 = _EVAL_12 == 3'h1;
  assign _EVAL_235 = _EVAL_80 & _EVAL_101;
  assign _EVAL_260 = _EVAL_14[0];
  assign _EVAL_159 = _EVAL_77 | _EVAL_257;
  assign _EVAL_110 = ~_EVAL_255;
  assign _EVAL_67 = _EVAL_8 == 3'h0;
  assign _EVAL_56 = ~_EVAL_25;
  assign _EVAL_20 = _EVAL_15 == _EVAL_98;
  assign _EVAL_104 = _EVAL_27 | _EVAL_17;
  assign _EVAL_199 = _EVAL_14[1];
  assign _EVAL_210 = _EVAL_92 | _EVAL_17;
  assign _EVAL_249 = ~_EVAL_274;
  assign _EVAL_51 = _EVAL_15 == 3'h2;
  assign _EVAL_130 = _EVAL_5 == _EVAL_76;
  assign _EVAL_263 = _EVAL_12 == 3'h5;
  assign _EVAL_65 = _EVAL_220 | _EVAL_17;
  assign _EVAL_69 = _EVAL_262 | _EVAL_17;
  assign _EVAL_160 = _EVAL_209 | _EVAL_17;
  assign _EVAL_43 = _EVAL & _EVAL_238;
  assign _EVAL_141 = ~_EVAL_183;
  assign _EVAL_73 = _EVAL_30 | _EVAL_17;
  assign _EVAL_242 = _EVAL & _EVAL_206;
  assign _EVAL_189 = _EVAL_39 | _EVAL_6;
  assign _EVAL_252 = _EVAL_2 == 2'h0;
  assign _EVAL_262 = _EVAL_12 <= 3'h6;
  assign _EVAL_83 = _EVAL_26 | _EVAL_17;
  assign _EVAL_131 = _EVAL_2 <= 2'h2;
  assign _EVAL_222 = _EVAL_146 == 4'h0;
  assign _EVAL_266 = plusarg_reader_out == 32'h0;
  assign _EVAL_29 = _EVAL_1 <= 3'h4;
  assign _EVAL_139 = _EVAL_235 ? _EVAL_165 : 8'h0;
  assign _EVAL_52 = _EVAL_0 & _EVAL_33;
  assign _EVAL_108 = {{28'd0}, _EVAL_185};
  assign _EVAL_57 = _EVAL_12 == 3'h0;
  assign _EVAL_154 = _EVAL_10 <= 2'h2;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_47 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_62 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_71 = _RAND_2[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_75 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_76 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_98 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_116 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_138 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_147 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_151 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_152 = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_175 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_211 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_241 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_243 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_268 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_272 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_7) begin
    if (_EVAL_17) begin
      _EVAL_47 <= 1'h0;
    end else if (_EVAL_240) begin
      if (_EVAL_23) begin
        _EVAL_47 <= 1'h0;
      end else begin
        _EVAL_47 <= _EVAL_190;
      end
    end
    if (_EVAL_17) begin
      _EVAL_62 <= 1'h0;
    end else if (_EVAL_60) begin
      if (_EVAL_142) begin
        _EVAL_62 <= 1'h0;
      end else begin
        _EVAL_62 <= _EVAL_121;
      end
    end
    if (_EVAL_195) begin
      _EVAL_71 <= _EVAL_14;
    end
    if (_EVAL_195) begin
      _EVAL_75 <= _EVAL_1;
    end
    if (_EVAL_267) begin
      _EVAL_76 <= _EVAL_5;
    end
    if (_EVAL_195) begin
      _EVAL_98 <= _EVAL_15;
    end
    if (_EVAL_17) begin
      _EVAL_116 <= 32'h0;
    end else if (_EVAL_229) begin
      _EVAL_116 <= 32'h0;
    end else begin
      _EVAL_116 <= _EVAL_86;
    end
    if (_EVAL_195) begin
      _EVAL_138 <= _EVAL_10;
    end
    if (_EVAL_267) begin
      _EVAL_147 <= _EVAL_2;
    end
    if (_EVAL_267) begin
      _EVAL_151 <= _EVAL_18;
    end
    if (_EVAL_17) begin
      _EVAL_152 <= 5'h0;
    end else begin
      _EVAL_152 <= _EVAL_259;
    end
    if (_EVAL_17) begin
      _EVAL_175 <= 1'h0;
    end else if (_EVAL_60) begin
      if (_EVAL_149) begin
        _EVAL_175 <= 1'h0;
      end else begin
        _EVAL_175 <= _EVAL_218;
      end
    end
    if (_EVAL_267) begin
      _EVAL_211 <= _EVAL_12;
    end
    if (_EVAL_195) begin
      _EVAL_241 <= _EVAL_8;
    end
    if (_EVAL_17) begin
      _EVAL_243 <= 1'h0;
    end else if (_EVAL_240) begin
      if (_EVAL_126) begin
        _EVAL_243 <= 1'h0;
      end else begin
        _EVAL_243 <= _EVAL_177;
      end
    end
    if (_EVAL_267) begin
      _EVAL_268 <= _EVAL_13;
    end
    if (_EVAL_267) begin
      _EVAL_272 <= _EVAL_3;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8de6ccab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4baab8bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5260c9e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b49aef20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27ec16e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4128b46b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89b6e733)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bb966f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df7289e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc87850f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8697490)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d30fdbc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e355979)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(898026bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d3aaa50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d7b8b6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17066053)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55c64379)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e93557b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(392c1af7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b57e530c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27b0a6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f87b9ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48ae5507)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9db450eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33e580e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b76f52d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(348edefe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d6cd263)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb10b563)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf652462)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69292c9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72f091b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df3751d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8aaf0a84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19a37425)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8511dbfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e9aa495)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f43c5305)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(838b8227)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13061bc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db496915)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78a4af06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18d04357)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12a519c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f721f2da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ce68870)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea6a2753)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2cf342a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b52c267)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1341f9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6270016)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94a100ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2cdd3e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c2c28a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95abb7c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0569570)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab779d75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd081c58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6ae0142)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bab55e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7c3d417)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c453e93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cc790d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60d9a538)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46e987a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1292e2e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11e6a41c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce55d102)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de4f7044)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23f0d0eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d439edd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46855bab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b9b61bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16e39e0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(310af077)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31e8f82c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f352c46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6f1616e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87f6c1f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(132eb8c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d98f173f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cd4908a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb9f1138)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3db870d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35e993da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce421ddf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7949eb65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cb87bf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d79b5a8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10a1a41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aeea1a27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d18cc9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
