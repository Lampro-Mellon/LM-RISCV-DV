//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_78_assert(
  input         _EVAL_0,
  input         _EVAL_2,
  input  [1:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  input  [2:0]  _EVAL_9,
  input  [2:0]  _EVAL_15,
  input  [2:0]  _EVAL_16,
  input  [1:0]  _EVAL_17,
  input         _EVAL_19,
  input         _EVAL_22,
  input  [2:0]  _EVAL_25,
  input  [25:0] _EVAL_26,
  input  [3:0]  _EVAL_27,
  input         _EVAL_29,
  input         _EVAL_31,
  input         _EVAL_32
);
  wire [1:0] TLMonitor__EVAL;
  wire  TLMonitor__EVAL_0;
  wire [25:0] TLMonitor__EVAL_1;
  wire [2:0] TLMonitor__EVAL_2;
  wire [2:0] TLMonitor__EVAL_3;
  wire [1:0] TLMonitor__EVAL_4;
  wire  TLMonitor__EVAL_5;
  wire  TLMonitor__EVAL_6;
  wire [3:0] TLMonitor__EVAL_7;
  wire  TLMonitor__EVAL_8;
  wire  TLMonitor__EVAL_9;
  wire [2:0] TLMonitor__EVAL_10;
  wire  TLMonitor__EVAL_11;
  wire [2:0] TLMonitor__EVAL_12;
  wire [2:0] TLMonitor__EVAL_13;
  wire  TLMonitor__EVAL_14;
  _EVAL_77_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14)
  );
  assign TLMonitor__EVAL_4 = _EVAL_4;
  assign TLMonitor__EVAL_0 = _EVAL_32;
  assign TLMonitor__EVAL_5 = _EVAL_29;
  assign TLMonitor__EVAL = _EVAL_17;
  assign TLMonitor__EVAL_9 = _EVAL_19;
  assign TLMonitor__EVAL_12 = _EVAL_25;
  assign TLMonitor__EVAL_13 = _EVAL_5;
  assign TLMonitor__EVAL_11 = _EVAL_22;
  assign TLMonitor__EVAL_8 = _EVAL_31;
  assign TLMonitor__EVAL_3 = _EVAL_16;
  assign TLMonitor__EVAL_1 = _EVAL_26;
  assign TLMonitor__EVAL_10 = _EVAL_9;
  assign TLMonitor__EVAL_6 = _EVAL_0;
  assign TLMonitor__EVAL_2 = _EVAL_15;
  assign TLMonitor__EVAL_14 = _EVAL_2;
  assign TLMonitor__EVAL_7 = _EVAL_27;

endmodule
