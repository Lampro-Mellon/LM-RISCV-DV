//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_45(
  output        _EVAL,
  input         _EVAL_0,
  output [2:0]  _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  output        _EVAL_4,
  output        _EVAL_5,
  input         _EVAL_6,
  output [31:0] _EVAL_7,
  input         _EVAL_8,
  output        _EVAL_9,
  input  [3:0]  _EVAL_10,
  output        _EVAL_11,
  input  [31:0] _EVAL_12,
  output [31:0] _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input  [31:0] _EVAL_18,
  output        _EVAL_19,
  output [3:0]  _EVAL_20,
  output        _EVAL_21,
  output        _EVAL_22,
  input  [31:0] _EVAL_23,
  input         _EVAL_24,
  output [3:0]  _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  output        _EVAL_28,
  output        _EVAL_29,
  output [31:0] _EVAL_30,
  output [1:0]  _EVAL_31,
  input  [3:0]  _EVAL_32,
  output        _EVAL_33,
  input  [2:0]  _EVAL_34,
  output [3:0]  _EVAL_35,
  input  [3:0]  _EVAL_36,
  output        _EVAL_37,
  input  [2:0]  _EVAL_38,
  output [2:0]  _EVAL_39,
  output        _EVAL_40,
  output [2:0]  _EVAL_41,
  output        _EVAL_42,
  input         _EVAL_43,
  output        _EVAL_44,
  output        _EVAL_45,
  input  [1:0]  _EVAL_46,
  input         _EVAL_47,
  input         _EVAL_48,
  output        _EVAL_49
);
  wire  Queue__EVAL;
  wire  Queue__EVAL_0;
  wire  Queue__EVAL_1;
  wire  Queue__EVAL_2;
  wire [2:0] Queue__EVAL_3;
  wire  Queue__EVAL_4;
  wire  Queue__EVAL_5;
  wire  Queue__EVAL_6;
  wire  Queue__EVAL_7;
  wire  Queue__EVAL_8;
  wire [3:0] Queue__EVAL_9;
  wire [31:0] Queue__EVAL_10;
  wire [2:0] Queue__EVAL_11;
  wire [31:0] Queue__EVAL_12;
  wire  Queue__EVAL_13;
  wire  Queue__EVAL_14;
  wire [3:0] Queue__EVAL_15;
  wire  Queue__EVAL_16;
  wire [31:0] Queue__EVAL_17;
  wire  Queue__EVAL_18;
  wire  Queue__EVAL_19;
  wire  Queue__EVAL_20;
  wire  Queue__EVAL_21;
  wire  Queue__EVAL_22;
  wire  Queue__EVAL_23;
  wire [3:0] Queue__EVAL_24;
  wire  Queue__EVAL_25;
  wire [3:0] Queue__EVAL_26;
  wire  Queue__EVAL_27;
  wire [31:0] Queue__EVAL_28;
  wire  Queue__EVAL_29;
  wire  Queue__EVAL_30;
  wire  Queue__EVAL_31;
  wire [2:0] Queue__EVAL_32;
  wire [2:0] Queue__EVAL_33;
  wire  Queue__EVAL_34;
  wire [1:0] Queue_1__EVAL;
  wire  Queue_1__EVAL_0;
  wire [2:0] Queue_1__EVAL_1;
  wire  Queue_1__EVAL_2;
  wire  Queue_1__EVAL_3;
  wire  Queue_1__EVAL_4;
  wire [31:0] Queue_1__EVAL_5;
  wire  Queue_1__EVAL_6;
  wire [31:0] Queue_1__EVAL_7;
  wire [2:0] Queue_1__EVAL_8;
  wire  Queue_1__EVAL_9;
  wire  Queue_1__EVAL_10;
  wire  Queue_1__EVAL_11;
  wire [1:0] Queue_1__EVAL_12;
  wire  Queue_1__EVAL_13;
  wire  Queue_1__EVAL_14;
  wire  Queue_1__EVAL_15;
  wire  Queue_1__EVAL_16;
  wire  Queue_1__EVAL_17;
  wire [3:0] Queue_1__EVAL_18;
  wire [3:0] Queue_1__EVAL_19;
  _EVAL_43 Queue (
    ._EVAL(Queue__EVAL),
    ._EVAL_0(Queue__EVAL_0),
    ._EVAL_1(Queue__EVAL_1),
    ._EVAL_2(Queue__EVAL_2),
    ._EVAL_3(Queue__EVAL_3),
    ._EVAL_4(Queue__EVAL_4),
    ._EVAL_5(Queue__EVAL_5),
    ._EVAL_6(Queue__EVAL_6),
    ._EVAL_7(Queue__EVAL_7),
    ._EVAL_8(Queue__EVAL_8),
    ._EVAL_9(Queue__EVAL_9),
    ._EVAL_10(Queue__EVAL_10),
    ._EVAL_11(Queue__EVAL_11),
    ._EVAL_12(Queue__EVAL_12),
    ._EVAL_13(Queue__EVAL_13),
    ._EVAL_14(Queue__EVAL_14),
    ._EVAL_15(Queue__EVAL_15),
    ._EVAL_16(Queue__EVAL_16),
    ._EVAL_17(Queue__EVAL_17),
    ._EVAL_18(Queue__EVAL_18),
    ._EVAL_19(Queue__EVAL_19),
    ._EVAL_20(Queue__EVAL_20),
    ._EVAL_21(Queue__EVAL_21),
    ._EVAL_22(Queue__EVAL_22),
    ._EVAL_23(Queue__EVAL_23),
    ._EVAL_24(Queue__EVAL_24),
    ._EVAL_25(Queue__EVAL_25),
    ._EVAL_26(Queue__EVAL_26),
    ._EVAL_27(Queue__EVAL_27),
    ._EVAL_28(Queue__EVAL_28),
    ._EVAL_29(Queue__EVAL_29),
    ._EVAL_30(Queue__EVAL_30),
    ._EVAL_31(Queue__EVAL_31),
    ._EVAL_32(Queue__EVAL_32),
    ._EVAL_33(Queue__EVAL_33),
    ._EVAL_34(Queue__EVAL_34)
  );
  _EVAL_44 Queue_1 (
    ._EVAL(Queue_1__EVAL),
    ._EVAL_0(Queue_1__EVAL_0),
    ._EVAL_1(Queue_1__EVAL_1),
    ._EVAL_2(Queue_1__EVAL_2),
    ._EVAL_3(Queue_1__EVAL_3),
    ._EVAL_4(Queue_1__EVAL_4),
    ._EVAL_5(Queue_1__EVAL_5),
    ._EVAL_6(Queue_1__EVAL_6),
    ._EVAL_7(Queue_1__EVAL_7),
    ._EVAL_8(Queue_1__EVAL_8),
    ._EVAL_9(Queue_1__EVAL_9),
    ._EVAL_10(Queue_1__EVAL_10),
    ._EVAL_11(Queue_1__EVAL_11),
    ._EVAL_12(Queue_1__EVAL_12),
    ._EVAL_13(Queue_1__EVAL_13),
    ._EVAL_14(Queue_1__EVAL_14),
    ._EVAL_15(Queue_1__EVAL_15),
    ._EVAL_16(Queue_1__EVAL_16),
    ._EVAL_17(Queue_1__EVAL_17),
    ._EVAL_18(Queue_1__EVAL_18),
    ._EVAL_19(Queue_1__EVAL_19)
  );
  assign Queue_1__EVAL_15 = _EVAL_24;
  assign Queue__EVAL = 1'h0;
  assign Queue_1__EVAL_4 = _EVAL_16;
  assign Queue_1__EVAL_8 = _EVAL_34;
  assign _EVAL_39 = Queue__EVAL_11;
  assign Queue__EVAL_18 = _EVAL_0;
  assign _EVAL_7 = Queue_1__EVAL_7;
  assign _EVAL_49 = Queue__EVAL_19;
  assign Queue__EVAL_12 = _EVAL_12;
  assign _EVAL_41 = Queue_1__EVAL_1;
  assign _EVAL_40 = Queue__EVAL_20;
  assign _EVAL_21 = Queue_1__EVAL_17;
  assign _EVAL_28 = Queue_1__EVAL_16;
  assign Queue_1__EVAL_0 = _EVAL_3;
  assign Queue__EVAL_7 = _EVAL_27;
  assign Queue__EVAL_29 = _EVAL_8;
  assign Queue__EVAL_33 = _EVAL_38;
  assign Queue__EVAL_32 = 3'h0;
  assign _EVAL_30 = Queue__EVAL_28;
  assign Queue__EVAL_30 = _EVAL_48;
  assign _EVAL_5 = Queue_1__EVAL_9;
  assign Queue__EVAL_4 = _EVAL_43;
  assign Queue__EVAL_24 = _EVAL_32;
  assign _EVAL_37 = Queue__EVAL_23;
  assign _EVAL_19 = Queue_1__EVAL_3;
  assign _EVAL_11 = Queue__EVAL_31;
  assign _EVAL_33 = Queue_1__EVAL_2;
  assign Queue__EVAL_1 = 1'h0;
  assign Queue_1__EVAL_14 = _EVAL_6;
  assign _EVAL_29 = Queue__EVAL_14;
  assign _EVAL_45 = Queue_1__EVAL_13;
  assign _EVAL_35 = Queue_1__EVAL_19;
  assign Queue_1__EVAL_6 = _EVAL_14;
  assign Queue_1__EVAL_5 = _EVAL_23;
  assign _EVAL_9 = Queue__EVAL_13;
  assign Queue__EVAL_25 = _EVAL_16;
  assign Queue_1__EVAL_18 = _EVAL_36;
  assign _EVAL_22 = Queue__EVAL_8;
  assign _EVAL_44 = Queue__EVAL_5;
  assign _EVAL_4 = Queue__EVAL_21;
  assign Queue__EVAL_0 = _EVAL_47;
  assign Queue__EVAL_34 = _EVAL_2;
  assign _EVAL_42 = Queue__EVAL_27;
  assign _EVAL_25 = Queue__EVAL_9;
  assign Queue__EVAL_6 = _EVAL_26;
  assign _EVAL = Queue__EVAL_16;
  assign Queue_1__EVAL_10 = _EVAL_17;
  assign Queue__EVAL_22 = 1'h0;
  assign Queue_1__EVAL_11 = _EVAL_15;
  assign _EVAL_31 = Queue_1__EVAL_12;
  assign Queue__EVAL_26 = _EVAL_10;
  assign Queue_1__EVAL = _EVAL_46;
  assign _EVAL_1 = Queue__EVAL_3;
  assign _EVAL_20 = Queue__EVAL_15;
  assign Queue__EVAL_2 = _EVAL_15;
  assign _EVAL_13 = Queue__EVAL_17;
  assign Queue__EVAL_10 = _EVAL_18;
endmodule
