//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_117_assert(
  input  [1:0] _EVAL,
  input  [2:0] _EVAL_0,
  input  [1:0] _EVAL_1,
  input        _EVAL_2,
  input        _EVAL_3,
  input        _EVAL_4,
  input  [2:0] _EVAL_5,
  input        _EVAL_6,
  input        _EVAL_7,
  input        _EVAL_8,
  input        _EVAL_9,
  input        _EVAL_10,
  input        _EVAL_11,
  input  [8:0] _EVAL_12,
  input  [3:0] _EVAL_13
);
  wire  _EVAL_14;
  reg  _EVAL_15;
  reg [31:0] _RAND_0;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  reg  _EVAL_28;
  reg [31:0] _RAND_1;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire [1:0] _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  reg [2:0] _EVAL_37;
  reg [31:0] _RAND_2;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire [32:0] _EVAL_45;
  wire [1:0] _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  reg  _EVAL_50;
  reg [31:0] _RAND_3;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_55;
  wire [8:0] _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  reg [1:0] _EVAL_76;
  reg [31:0] _RAND_4;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  reg  _EVAL_80;
  reg [31:0] _RAND_5;
  reg  _EVAL_81;
  reg [31:0] _RAND_6;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  reg [31:0] _EVAL_85;
  reg [31:0] _RAND_7;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire [9:0] _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire [3:0] _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire [1:0] _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  reg  _EVAL_113;
  reg [31:0] _RAND_8;
  wire  _EVAL_114;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire [31:0] _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  reg [1:0] _EVAL_123;
  reg [31:0] _RAND_9;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire [1:0] _EVAL_128;
  wire [9:0] _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire [1:0] _EVAL_133;
  wire  _EVAL_134;
  reg [8:0] _EVAL_135;
  reg [31:0] _RAND_10;
  wire  _EVAL_136;
  wire [9:0] _EVAL_137;
  wire  _EVAL_138;
  reg [2:0] _EVAL_139;
  reg [31:0] _RAND_11;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire [1:0] _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  reg  _EVAL_163;
  reg [31:0] _RAND_12;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_93 = ~_EVAL_81;
  assign _EVAL_121 = _EVAL_0 == 3'h0;
  assign _EVAL_122 = ~_EVAL_48;
  assign _EVAL_41 = _EVAL_0 == 3'h4;
  assign _EVAL_74 = _EVAL_27 | _EVAL_16;
  assign _EVAL_101 = _EVAL_0 == 3'h7;
  assign _EVAL_73 = _EVAL_6 & _EVAL_31;
  assign _EVAL_154 = _EVAL_133[0];
  assign _EVAL_160 = _EVAL_6 & _EVAL_47;
  assign _EVAL_14 = _EVAL_4 & _EVAL_49;
  assign _EVAL_167 = ~_EVAL_91;
  assign _EVAL_134 = ~_EVAL_67;
  assign _EVAL_164 = _EVAL_70 | _EVAL_16;
  assign _EVAL_70 = _EVAL_11 == _EVAL_50;
  assign _EVAL_159 = _EVAL_6 & _EVAL_103;
  assign _EVAL_124 = ~_EVAL_80;
  assign _EVAL_24 = ~_EVAL_156;
  assign _EVAL_31 = _EVAL_5 == 3'h1;
  assign _EVAL_59 = _EVAL_46[0];
  assign _EVAL_89 = _EVAL_108[0];
  assign _EVAL_45 = _EVAL_85 + 32'h1;
  assign _EVAL_77 = _EVAL_107 & _EVAL_124;
  assign _EVAL_161 = _EVAL_25 | _EVAL_16;
  assign _EVAL_56 = _EVAL_12 & 9'h3;
  assign _EVAL_87 = _EVAL_33[0];
  assign _EVAL_114 = _EVAL_6 & _EVAL_65;
  assign _EVAL_27 = _EVAL_3 == _EVAL_163;
  assign _EVAL_49 = _EVAL_0 == 3'h5;
  assign _EVAL_26 = ~_EVAL_68;
  assign _EVAL_36 = _EVAL_13 == 4'hf;
  assign _EVAL_88 = ~_EVAL_69;
  assign _EVAL_19 = _EVAL_155 | _EVAL_16;
  assign _EVAL_30 = _EVAL_149 | _EVAL_16;
  assign _EVAL_102 = $signed(_EVAL_129) == 10'sh0;
  assign _EVAL_58 = _EVAL_0 == 3'h2;
  assign _EVAL_46 = _EVAL_15 - 1'h1;
  assign _EVAL_146 = _EVAL_5 == _EVAL_37;
  assign _EVAL_103 = _EVAL_5 == 3'h2;
  assign _EVAL_23 = ~_EVAL_18;
  assign _EVAL_111 = ~_EVAL_126;
  assign _EVAL_143 = _EVAL_128[0];
  assign _EVAL_78 = _EVAL_56 == 9'h0;
  assign _EVAL_71 = _EVAL_152 | _EVAL_20;
  assign _EVAL_44 = _EVAL_4 & _EVAL_117;
  assign _EVAL_162 = _EVAL_4 & _EVAL_121;
  assign _EVAL_133 = _EVAL_84 ? 2'h1 : 2'h0;
  assign _EVAL_99 = {1'b0,$signed(_EVAL_12)};
  assign _EVAL_42 = _EVAL_138 | _EVAL_7;
  assign _EVAL_138 = ~_EVAL_11;
  assign _EVAL_150 = _EVAL_28 - 1'h1;
  assign _EVAL_61 = _EVAL_138 | _EVAL_16;
  assign _EVAL_157 = _EVAL_22 | _EVAL_16;
  assign _EVAL_75 = _EVAL_93 | _EVAL_16;
  assign _EVAL_136 = _EVAL_6 & _EVAL_88;
  assign _EVAL_131 = ~_EVAL_7;
  assign _EVAL_94 = _EVAL_86 | _EVAL_16;
  assign _EVAL_18 = _EVAL_35 | _EVAL_16;
  assign _EVAL_40 = ~_EVAL_161;
  assign _EVAL_32 = ~_EVAL_157;
  assign _EVAL_128 = _EVAL_66 ? 2'h1 : 2'h0;
  assign _EVAL_98 = _EVAL_0 == 3'h1;
  assign _EVAL_145 = _EVAL_150[0];
  assign _EVAL_106 = ~_EVAL_74;
  assign _EVAL_104 = _EVAL_92 | _EVAL_16;
  assign _EVAL_38 = ~_EVAL_61;
  assign _EVAL_60 = ~_EVAL_19;
  assign _EVAL_57 = ~_EVAL_75;
  assign _EVAL_21 = _EVAL_4 & _EVAL_101;
  assign _EVAL_129 = _EVAL_137;
  assign _EVAL_84 = _EVAL_53 & _EVAL_158;
  assign _EVAL_108 = _EVAL_80 - 1'h1;
  assign _EVAL_72 = ~_EVAL_164;
  assign _EVAL_33 = _EVAL_113 - 1'h1;
  assign _EVAL_141 = _EVAL_36 | _EVAL_16;
  assign _EVAL_137 = $signed(_EVAL_99) & -10'sh200;
  assign _EVAL_35 = _EVAL_1 <= 2'h2;
  assign _EVAL_100 = ~_EVAL_147;
  assign _EVAL_151 = _EVAL_4 & _EVAL_58;
  assign _EVAL_166 = _EVAL_1 != 2'h2;
  assign _EVAL_53 = _EVAL_39 & _EVAL_83;
  assign _EVAL_67 = _EVAL_166 | _EVAL_16;
  assign _EVAL_48 = _EVAL_78 | _EVAL_16;
  assign _EVAL_97 = _EVAL_131 | _EVAL_16;
  assign _EVAL_54 = _EVAL >= 2'h2;
  assign _EVAL_65 = _EVAL_5 == 3'h5;
  assign _EVAL_82 = _EVAL_4 & _EVAL_118;
  assign _EVAL_112 = ~_EVAL_51;
  assign _EVAL_34 = ~_EVAL_104;
  assign _EVAL_22 = _EVAL_1 == 2'h0;
  assign _EVAL_17 = _EVAL_4 & _EVAL_41;
  assign _EVAL_51 = _EVAL_109 | _EVAL_16;
  assign _EVAL_110 = _EVAL_5 == 3'h6;
  assign _EVAL_152 = _EVAL_93 | _EVAL_132;
  assign _EVAL_127 = _EVAL_6 & _EVAL_110;
  assign _EVAL_153 = _EVAL_39 & _EVAL_69;
  assign _EVAL_90 = _EVAL_146 | _EVAL_16;
  assign _EVAL_16 = _EVAL_2;
  assign _EVAL_25 = _EVAL_143 | _EVAL_81;
  assign _EVAL_86 = _EVAL_1 == _EVAL_76;
  assign _EVAL_147 = _EVAL_42 | _EVAL_16;
  assign _EVAL_69 = ~_EVAL_28;
  assign _EVAL_118 = _EVAL_0 == 3'h6;
  assign _EVAL_63 = ~_EVAL_90;
  assign _EVAL_109 = _EVAL_5 <= 3'h6;
  assign _EVAL_117 = ~_EVAL_124;
  assign _EVAL_105 = ~_EVAL_13;
  assign _EVAL_91 = _EVAL_71 | _EVAL_16;
  assign _EVAL_155 = _EVAL_0 == _EVAL_139;
  assign _EVAL_158 = ~_EVAL_110;
  assign _EVAL_55 = ~_EVAL_141;
  assign _EVAL_62 = _EVAL_6 & _EVAL_52;
  assign _EVAL_20 = _EVAL_85 < plusarg_reader_out;
  assign _EVAL_83 = ~_EVAL_15;
  assign _EVAL_66 = _EVAL_107 & _EVAL_165;
  assign _EVAL_52 = _EVAL_5 == 3'h0;
  assign _EVAL_39 = _EVAL_8 & _EVAL_6;
  assign _EVAL_126 = _EVAL_95 | _EVAL_16;
  assign _EVAL_142 = _EVAL_81 | _EVAL_143;
  assign _EVAL_120 = _EVAL_45[31:0];
  assign _EVAL_148 = _EVAL_4 & _EVAL_79;
  assign _EVAL_149 = _EVAL_12 == _EVAL_135;
  assign _EVAL_130 = ~_EVAL_94;
  assign _EVAL_64 = ~_EVAL_30;
  assign _EVAL_119 = ~_EVAL_97;
  assign _EVAL_68 = _EVAL_102 | _EVAL_16;
  assign _EVAL_156 = _EVAL_54 | _EVAL_16;
  assign _EVAL_95 = _EVAL == _EVAL_123;
  assign _EVAL_92 = _EVAL_105 == 4'h0;
  assign _EVAL_79 = _EVAL_0 == 3'h3;
  assign _EVAL_47 = _EVAL_5 == 3'h4;
  assign _EVAL_29 = ~_EVAL_16;
  assign _EVAL_165 = ~_EVAL_113;
  assign _EVAL_125 = _EVAL_107 | _EVAL_39;
  assign _EVAL_116 = _EVAL_4 & _EVAL_98;
  assign _EVAL_132 = plusarg_reader_out == 32'h0;
  assign _EVAL_43 = ~_EVAL_154;
  assign _EVAL_107 = _EVAL_10 & _EVAL_4;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_28 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_37 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_50 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_76 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_80 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_81 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_85 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_113 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_123 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_135 = _RAND_10[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_139 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_163 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  if (_EVAL_2) begin
    _EVAL_15 = 1'h0;
  end
  if (_EVAL_2) begin
    _EVAL_28 = 1'h0;
  end
  if (_EVAL_2) begin
    _EVAL_80 = 1'h0;
  end
  if (_EVAL_2) begin
    _EVAL_81 = 1'h0;
  end
  if (_EVAL_2) begin
    _EVAL_85 = 32'h0;
  end
  if (_EVAL_2) begin
    _EVAL_113 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_9) begin
    if (_EVAL_153) begin
      _EVAL_37 <= _EVAL_5;
    end
    if (_EVAL_153) begin
      _EVAL_50 <= _EVAL_11;
    end
    if (_EVAL_153) begin
      _EVAL_76 <= _EVAL_1;
    end
    if (_EVAL_153) begin
      _EVAL_123 <= _EVAL;
    end
    if (_EVAL_77) begin
      _EVAL_135 <= _EVAL_12;
    end
    if (_EVAL_77) begin
      _EVAL_139 <= _EVAL_0;
    end
    if (_EVAL_153) begin
      _EVAL_163 <= _EVAL_3;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1ec2fa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47c0262e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad505ef0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19c3930a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f56d784e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(543d727b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4005fd0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1f36b7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(412a66d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb623721)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d0a88a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f415309c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(390f60fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a17cbab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(195d83e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da9f1d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd8449a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b65d73b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48d9b615)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f8582)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(caecec5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f79b7a8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcfe01e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8b6d7d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21a6a828)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef242ed5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3cd82ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7fe1346)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e90c14db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ebf9f81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd0d650e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11881bbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e40cb47e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(172674c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8205e43e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba86b81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20abaf66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6328756)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(902750c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1482ab4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e377f34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c72d938)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be6f55b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e584df8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fd23de3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a54ed39e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d76d673e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4a3038e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f040e8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37c4b639)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b8c4cef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f47ff4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47cb3f55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bc1cd2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f493ca8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(201fcf3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a4b008c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge _EVAL_9 or posedge _EVAL_2) begin
    if (_EVAL_2) begin
      _EVAL_15 <= 1'h0;
    end else if (_EVAL_39) begin
      if (_EVAL_83) begin
        _EVAL_15 <= 1'h0;
      end else begin
        _EVAL_15 <= _EVAL_59;
      end
    end
  end
  always @(posedge _EVAL_9 or posedge _EVAL_2) begin
    if (_EVAL_2) begin
      _EVAL_28 <= 1'h0;
    end else if (_EVAL_39) begin
      if (_EVAL_69) begin
        _EVAL_28 <= 1'h0;
      end else begin
        _EVAL_28 <= _EVAL_145;
      end
    end
  end
  always @(posedge _EVAL_9 or posedge _EVAL_2) begin
    if (_EVAL_2) begin
      _EVAL_80 <= 1'h0;
    end else if (_EVAL_107) begin
      if (_EVAL_124) begin
        _EVAL_80 <= 1'h0;
      end else begin
        _EVAL_80 <= _EVAL_89;
      end
    end
  end
  always @(posedge _EVAL_9 or posedge _EVAL_2) begin
    if (_EVAL_2) begin
      _EVAL_81 <= 1'h0;
    end else begin
      _EVAL_81 <= _EVAL_142 & _EVAL_43;
    end
  end
  always @(posedge _EVAL_9 or posedge _EVAL_2) begin
    if (_EVAL_2) begin
      _EVAL_85 <= 32'h0;
    end else if (_EVAL_125) begin
      _EVAL_85 <= 32'h0;
    end else begin
      _EVAL_85 <= _EVAL_120;
    end
  end
  always @(posedge _EVAL_9 or posedge _EVAL_2) begin
    if (_EVAL_2) begin
      _EVAL_113 <= 1'h0;
    end else if (_EVAL_107) begin
      if (_EVAL_165) begin
        _EVAL_113 <= 1'h0;
      end else begin
        _EVAL_113 <= _EVAL_87;
      end
    end
  end

endmodule
