//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_137_assert(
  input  [1:0] _EVAL,
  input        _EVAL_0,
  input        _EVAL_1,
  input        _EVAL_2,
  input        _EVAL_3,
  input        _EVAL_4,
  input  [1:0] _EVAL_5,
  input  [2:0] _EVAL_6,
  input  [3:0] _EVAL_7,
  input        _EVAL_8,
  input        _EVAL_9,
  input        _EVAL_10,
  input  [2:0] _EVAL_11,
  input  [2:0] _EVAL_12,
  input        _EVAL_13,
  input  [8:0] _EVAL_14
);
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire [9:0] _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire [3:0] _EVAL_21;
  wire [1:0] _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  reg [2:0] _EVAL_31;
  reg [31:0] _RAND_0;
  wire [1:0] _EVAL_32;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire [8:0] _EVAL_39;
  reg  _EVAL_40;
  reg [31:0] _RAND_1;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire [4:0] _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire [1:0] _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire [9:0] _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire [9:0] _EVAL_73;
  wire [1:0] _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire [9:0] _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire [8:0] _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  reg  _EVAL_97;
  reg [31:0] _RAND_2;
  wire [1:0] _EVAL_98;
  wire [31:0] _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire [3:0] _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire [3:0] _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire [9:0] _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire [9:0] _EVAL_134;
  reg [1:0] _EVAL_135;
  reg [31:0] _RAND_3;
  wire  _EVAL_136;
  wire [9:0] _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire [1:0] _EVAL_140;
  wire [1:0] _EVAL_141;
  wire  _EVAL_142;
  reg  _EVAL_143;
  reg [31:0] _RAND_4;
  wire  _EVAL_144;
  wire [9:0] _EVAL_145;
  wire [8:0] _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_149;
  wire [3:0] _EVAL_150;
  wire  _EVAL_151;
  wire [1:0] _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire [9:0] _EVAL_157;
  wire [9:0] _EVAL_158;
  wire  _EVAL_159;
  reg [31:0] _EVAL_161;
  reg [31:0] _RAND_5;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire [9:0] _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire [9:0] _EVAL_177;
  reg [2:0] _EVAL_178;
  reg [31:0] _RAND_6;
  wire  _EVAL_179;
  wire [9:0] _EVAL_180;
  wire  _EVAL_181;
  wire [32:0] _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_187;
  reg  _EVAL_188;
  reg [31:0] _RAND_7;
  wire  _EVAL_189;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  reg  _EVAL_196;
  reg [31:0] _RAND_8;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire [8:0] _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire [8:0] _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire [1:0] _EVAL_215;
  reg  _EVAL_216;
  reg [31:0] _RAND_9;
  wire [1:0] _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire [9:0] _EVAL_223;
  reg [1:0] _EVAL_224;
  reg [31:0] _RAND_10;
  wire [1:0] _EVAL_225;
  wire [9:0] _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  reg [8:0] _EVAL_236;
  reg [31:0] _RAND_11;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire [9:0] _EVAL_243;
  wire [9:0] _EVAL_244;
  wire  _EVAL_245;
  reg [2:0] _EVAL_246;
  reg [31:0] _RAND_12;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire [8:0] _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_252;
  wire [9:0] _EVAL_253;
  wire [8:0] _EVAL_254;
  wire  _EVAL_256;
  wire  _EVAL_257;
  reg  _EVAL_258;
  reg [31:0] _RAND_13;
  wire  _EVAL_259;
  wire [1:0] _EVAL_260;
  wire  _EVAL_261;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_197 = _EVAL_6 == 3'h6;
  assign _EVAL_58 = _EVAL_208 & _EVAL_212;
  assign _EVAL_165 = _EVAL_8 == _EVAL_97;
  assign _EVAL_95 = _EVAL_168 | _EVAL_2;
  assign _EVAL_114 = _EVAL_3 & _EVAL_238;
  assign _EVAL_209 = _EVAL_14 ^ 9'h100;
  assign _EVAL_123 = _EVAL_138 & _EVAL_239;
  assign _EVAL_261 = _EVAL_6 == 3'h3;
  assign _EVAL_118 = _EVAL_7 & _EVAL_21;
  assign _EVAL_223 = _EVAL_126;
  assign _EVAL_228 = _EVAL_43 | _EVAL_2;
  assign _EVAL_62 = _EVAL_213 | _EVAL_2;
  assign _EVAL_185 = _EVAL_75 | _EVAL_2;
  assign _EVAL_57 = _EVAL_4 & _EVAL_49;
  assign _EVAL_16 = ~_EVAL_237;
  assign _EVAL_215 = _EVAL_188 - 1'h1;
  assign _EVAL_17 = $signed(_EVAL_243) & -10'sh100;
  assign _EVAL_241 = _EVAL_4 & _EVAL_195;
  assign _EVAL_126 = $signed(_EVAL_226) & -10'sh40;
  assign _EVAL_189 = ~_EVAL_234;
  assign _EVAL_44 = ~_EVAL_40;
  assign _EVAL_206 = _EVAL_163 & _EVAL_153;
  assign _EVAL_39 = {{7'd0}, _EVAL_98};
  assign _EVAL_122 = _EVAL_6 == 3'h5;
  assign _EVAL_111 = _EVAL_162 | _EVAL_2;
  assign _EVAL_110 = _EVAL_11 != 3'h0;
  assign _EVAL_54 = ~_EVAL_147;
  assign _EVAL_71 = _EVAL_254 == 9'h0;
  assign _EVAL_82 = _EVAL_12 == 3'h0;
  assign _EVAL_49 = _EVAL_12 == 3'h1;
  assign _EVAL_51 = ~_EVAL_61;
  assign _EVAL_100 = ~_EVAL_94;
  assign _EVAL_98 = ~_EVAL_141;
  assign _EVAL_229 = _EVAL_6 == _EVAL_31;
  assign _EVAL_141 = _EVAL_45[1:0];
  assign _EVAL_234 = _EVAL_165 | _EVAL_2;
  assign _EVAL_85 = _EVAL_121 >> _EVAL_0;
  assign _EVAL_237 = _EVAL_92 | _EVAL_2;
  assign _EVAL_43 = ~_EVAL_8;
  assign _EVAL_90 = _EVAL_138 & _EVAL_170;
  assign _EVAL_175 = ~_EVAL_218;
  assign _EVAL_145 = $signed(_EVAL_68) & -10'sh4;
  assign _EVAL_164 = _EVAL_12 == _EVAL_246;
  assign _EVAL_180 = {1'b0,$signed(_EVAL_201)};
  assign _EVAL_200 = _EVAL_161 < plusarg_reader_out;
  assign _EVAL_194 = _EVAL_20 | _EVAL_124;
  assign _EVAL_173 = $signed(_EVAL_244) & -10'sh80;
  assign _EVAL_195 = _EVAL_12 == 3'h2;
  assign _EVAL_96 = plusarg_reader_out == 32'h0;
  assign _EVAL_238 = _EVAL_6 == 3'h0;
  assign _EVAL_177 = $signed(_EVAL_180) & -10'sh18;
  assign _EVAL_243 = {1'b0,$signed(_EVAL_209)};
  assign _EVAL_167 = ~_EVAL_107;
  assign _EVAL_193 = _EVAL_69 | _EVAL_123;
  assign _EVAL_30 = ~_EVAL_0;
  assign _EVAL_66 = _EVAL_13 & _EVAL_3;
  assign _EVAL_88 = _EVAL_14 == _EVAL_236;
  assign _EVAL_73 = _EVAL_173;
  assign _EVAL_198 = _EVAL_250 | _EVAL_136;
  assign _EVAL_69 = _EVAL_15 | _EVAL_64;
  assign _EVAL_138 = _EVAL_53[0];
  assign _EVAL_146 = _EVAL_14 ^ 9'h44;
  assign _EVAL_101 = _EVAL_3 & _EVAL_54;
  assign _EVAL_108 = _EVAL_74[0];
  assign _EVAL_251 = _EVAL_3 & _EVAL_154;
  assign _EVAL_252 = _EVAL_3 & _EVAL_23;
  assign _EVAL_214 = _EVAL_11 <= 3'h4;
  assign _EVAL_170 = _EVAL_245 & _EVAL_174;
  assign _EVAL_254 = _EVAL_14 & _EVAL_39;
  assign _EVAL_151 = _EVAL_198 | _EVAL_248;
  assign _EVAL_86 = _EVAL_14 ^ 9'h60;
  assign _EVAL_81 = _EVAL_4 & _EVAL_104;
  assign _EVAL_149 = _EVAL_66 & _EVAL_147;
  assign _EVAL_259 = ~_EVAL_139;
  assign _EVAL_157 = _EVAL_177;
  assign _EVAL_156 = _EVAL_143 | _EVAL_204;
  assign _EVAL_226 = {1'b0,$signed(_EVAL_14)};
  assign _EVAL_36 = _EVAL_199 & _EVAL_159;
  assign _EVAL_55 = ~_EVAL_63;
  assign _EVAL_248 = $signed(_EVAL_80) == 10'sh0;
  assign _EVAL_119 = $signed(_EVAL_137) == 10'sh0;
  assign _EVAL_201 = _EVAL_14 ^ 9'h48;
  assign _EVAL_67 = _EVAL_52 | _EVAL_200;
  assign _EVAL_84 = _EVAL_156 & _EVAL_169;
  assign _EVAL_99 = _EVAL_182[31:0];
  assign _EVAL_213 = _EVAL_166 & _EVAL_151;
  assign _EVAL_220 = _EVAL_91 | _EVAL_2;
  assign _EVAL_174 = ~_EVAL_212;
  assign _EVAL_247 = _EVAL_140[0];
  assign _EVAL_48 = _EVAL_131 & _EVAL_208;
  assign _EVAL_144 = _EVAL_66 | _EVAL_163;
  assign _EVAL_115 = _EVAL_225[0];
  assign _EVAL_79 = _EVAL_66 & _EVAL_83;
  assign _EVAL_222 = ~_EVAL_2;
  assign _EVAL_153 = ~_EVAL_216;
  assign _EVAL_26 = _EVAL_118 == 4'h0;
  assign _EVAL_23 = _EVAL_6 == 3'h1;
  assign _EVAL_78 = ~_EVAL_19;
  assign _EVAL_249 = _EVAL_14 ^ 9'h80;
  assign _EVAL_131 = _EVAL_53[1];
  assign _EVAL_217 = 2'h1 << _EVAL_8;
  assign _EVAL_199 = _EVAL_163 & _EVAL_44;
  assign _EVAL_83 = ~_EVAL_258;
  assign _EVAL_210 = _EVAL_4 & _EVAL_35;
  assign _EVAL_235 = _EVAL_187 | _EVAL_2;
  assign _EVAL_244 = {1'b0,$signed(_EVAL_249)};
  assign _EVAL_240 = _EVAL_6 == 3'h4;
  assign _EVAL_137 = _EVAL_134;
  assign _EVAL_202 = _EVAL_11 == _EVAL_178;
  assign _EVAL_187 = _EVAL_0 == _EVAL_196;
  assign _EVAL_134 = $signed(_EVAL_158) & -10'sh20;
  assign _EVAL_63 = _EVAL_202 | _EVAL_2;
  assign _EVAL_163 = _EVAL_9 & _EVAL_4;
  assign _EVAL_38 = _EVAL_138 & _EVAL_116;
  assign _EVAL_53 = _EVAL_22 | 2'h1;
  assign _EVAL_94 = _EVAL_41 | _EVAL_2;
  assign _EVAL_104 = _EVAL_12 == 3'h6;
  assign _EVAL_253 = _EVAL_145;
  assign _EVAL_102 = _EVAL_215[0];
  assign _EVAL_207 = ~_EVAL_181;
  assign _EVAL_52 = _EVAL_133 | _EVAL_96;
  assign _EVAL_42 = _EVAL_12 == 3'h4;
  assign _EVAL_45 = 5'h3 << _EVAL;
  assign _EVAL_68 = {1'b0,$signed(_EVAL_146)};
  assign _EVAL_120 = _EVAL_4 & _EVAL_132;
  assign _EVAL_80 = _EVAL_17;
  assign _EVAL_233 = ~_EVAL_257;
  assign _EVAL_179 = _EVAL_6 == 3'h2;
  assign _EVAL_158 = {1'b0,$signed(_EVAL_86)};
  assign _EVAL_35 = ~_EVAL_153;
  assign _EVAL_64 = _EVAL_131 & _EVAL_245;
  assign _EVAL_166 = _EVAL <= 2'h2;
  assign _EVAL_37 = _EVAL_242 | _EVAL_60;
  assign _EVAL_130 = ~_EVAL_235;
  assign _EVAL_257 = _EVAL_67 | _EVAL_2;
  assign _EVAL_116 = _EVAL_208 & _EVAL_174;
  assign _EVAL_133 = ~_EVAL_143;
  assign _EVAL_150 = ~_EVAL_7;
  assign _EVAL_77 = ~_EVAL_111;
  assign _EVAL_106 = $signed(_EVAL_253) == 10'sh0;
  assign _EVAL_121 = _EVAL_204 | _EVAL_143;
  assign _EVAL_204 = _EVAL_152[0];
  assign _EVAL_136 = $signed(_EVAL_73) == 10'sh0;
  assign _EVAL_260 = _EVAL_216 - 1'h1;
  assign _EVAL_47 = _EVAL_214 | _EVAL_2;
  assign _EVAL_176 = _EVAL_11 <= 3'h1;
  assign _EVAL_230 = _EVAL_26 | _EVAL_2;
  assign _EVAL_19 = _EVAL_205 | _EVAL_2;
  assign _EVAL_155 = _EVAL_3 & _EVAL_240;
  assign _EVAL_219 = ~_EVAL_70;
  assign _EVAL_72 = _EVAL_71 | _EVAL_2;
  assign _EVAL_227 = ~_EVAL_29;
  assign _EVAL_192 = _EVAL_150 == 4'h0;
  assign _EVAL_28 = _EVAL_5 >= 2'h2;
  assign _EVAL_41 = _EVAL_5 == _EVAL_135;
  assign _EVAL_105 = {_EVAL_193,_EVAL_65,_EVAL_37,_EVAL_93};
  assign _EVAL_171 = _EVAL_110 | _EVAL_2;
  assign _EVAL_124 = $signed(_EVAL_157) == 10'sh0;
  assign _EVAL_242 = _EVAL_15 | _EVAL_48;
  assign _EVAL_93 = _EVAL_242 | _EVAL_38;
  assign _EVAL_154 = _EVAL_6 == 3'h7;
  assign _EVAL_129 = ~_EVAL_228;
  assign _EVAL_70 = _EVAL_183 | _EVAL_2;
  assign _EVAL_125 = _EVAL_260[0];
  assign _EVAL_87 = _EVAL_143 >> _EVAL_8;
  assign _EVAL_218 = _EVAL_30 | _EVAL_2;
  assign _EVAL_27 = _EVAL_85 | _EVAL_2;
  assign _EVAL_76 = ~_EVAL_171;
  assign _EVAL_142 = _EVAL[0];
  assign _EVAL_208 = ~_EVAL_245;
  assign _EVAL_203 = ~_EVAL_230;
  assign _EVAL_211 = ~_EVAL_47;
  assign _EVAL_182 = _EVAL_161 + 32'h1;
  assign _EVAL_162 = _EVAL_12 <= 3'h6;
  assign _EVAL_169 = ~_EVAL_108;
  assign _EVAL_221 = _EVAL_3 & _EVAL_197;
  assign _EVAL_20 = _EVAL_113 | _EVAL_106;
  assign _EVAL_183 = _EVAL_11 <= 3'h3;
  assign _EVAL_245 = _EVAL_14[1];
  assign _EVAL_59 = ~_EVAL_87;
  assign _EVAL_139 = _EVAL_15 | _EVAL_2;
  assign _EVAL_91 = ~_EVAL_10;
  assign _EVAL_15 = _EVAL >= 2'h2;
  assign _EVAL_132 = _EVAL_12 == 3'h5;
  assign _EVAL_65 = _EVAL_69 | _EVAL_90;
  assign _EVAL_232 = _EVAL_4 & _EVAL_82;
  assign _EVAL_103 = ~_EVAL_95;
  assign _EVAL_147 = ~_EVAL_188;
  assign _EVAL_74 = _EVAL_36 ? _EVAL_32 : 2'h0;
  assign _EVAL_89 = ~_EVAL_220;
  assign _EVAL_61 = _EVAL_229 | _EVAL_2;
  assign _EVAL_205 = _EVAL_11 == 3'h0;
  assign _EVAL_29 = _EVAL_192 | _EVAL_2;
  assign _EVAL_22 = 2'h1 << _EVAL_142;
  assign _EVAL_212 = _EVAL_14[0];
  assign _EVAL_75 = _EVAL_7 == _EVAL_105;
  assign _EVAL_25 = ~_EVAL_62;
  assign _EVAL_21 = ~_EVAL_105;
  assign _EVAL_60 = _EVAL_138 & _EVAL_58;
  assign _EVAL_32 = 2'h1 << _EVAL_0;
  assign _EVAL_18 = ~_EVAL_72;
  assign _EVAL_113 = $signed(_EVAL_223) == 10'sh0;
  assign _EVAL_250 = _EVAL_194 | _EVAL_119;
  assign _EVAL_127 = ~_EVAL_24;
  assign _EVAL_231 = ~_EVAL_185;
  assign _EVAL_191 = ~_EVAL_27;
  assign _EVAL_168 = _EVAL == _EVAL_224;
  assign _EVAL_92 = _EVAL_11 <= 3'h2;
  assign _EVAL_184 = _EVAL_4 & _EVAL_42;
  assign _EVAL_46 = _EVAL_59 | _EVAL_2;
  assign _EVAL_239 = _EVAL_245 & _EVAL_212;
  assign _EVAL_34 = ~_EVAL_256;
  assign _EVAL_181 = _EVAL_164 | _EVAL_2;
  assign _EVAL_159 = ~_EVAL_104;
  assign _EVAL_172 = ~_EVAL_46;
  assign _EVAL_107 = _EVAL_28 | _EVAL_2;
  assign _EVAL_152 = _EVAL_79 ? _EVAL_217 : 2'h0;
  assign _EVAL_24 = _EVAL_88 | _EVAL_2;
  assign _EVAL_140 = _EVAL_258 - 1'h1;
  assign _EVAL_256 = _EVAL_176 | _EVAL_2;
  assign _EVAL_128 = _EVAL_3 & _EVAL_122;
  assign _EVAL_112 = _EVAL_3 & _EVAL_261;
  assign _EVAL_56 = _EVAL_3 & _EVAL_179;
  assign _EVAL_225 = _EVAL_40 - 1'h1;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_31 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_40 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_97 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_135 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_143 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_161 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_178 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_188 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_196 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_216 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_224 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_236 = _RAND_11[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_246 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_258 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_1) begin
    if (_EVAL_149) begin
      _EVAL_31 <= _EVAL_6;
    end
    if (_EVAL_2) begin
      _EVAL_40 <= 1'h0;
    end else if (_EVAL_163) begin
      if (_EVAL_44) begin
        _EVAL_40 <= 1'h0;
      end else begin
        _EVAL_40 <= _EVAL_115;
      end
    end
    if (_EVAL_149) begin
      _EVAL_97 <= _EVAL_8;
    end
    if (_EVAL_206) begin
      _EVAL_135 <= _EVAL_5;
    end
    if (_EVAL_2) begin
      _EVAL_143 <= 1'h0;
    end else begin
      _EVAL_143 <= _EVAL_84;
    end
    if (_EVAL_2) begin
      _EVAL_161 <= 32'h0;
    end else if (_EVAL_144) begin
      _EVAL_161 <= 32'h0;
    end else begin
      _EVAL_161 <= _EVAL_99;
    end
    if (_EVAL_149) begin
      _EVAL_178 <= _EVAL_11;
    end
    if (_EVAL_2) begin
      _EVAL_188 <= 1'h0;
    end else if (_EVAL_66) begin
      if (_EVAL_147) begin
        _EVAL_188 <= 1'h0;
      end else begin
        _EVAL_188 <= _EVAL_102;
      end
    end
    if (_EVAL_206) begin
      _EVAL_196 <= _EVAL_0;
    end
    if (_EVAL_2) begin
      _EVAL_216 <= 1'h0;
    end else if (_EVAL_163) begin
      if (_EVAL_153) begin
        _EVAL_216 <= 1'h0;
      end else begin
        _EVAL_216 <= _EVAL_125;
      end
    end
    if (_EVAL_149) begin
      _EVAL_224 <= _EVAL;
    end
    if (_EVAL_149) begin
      _EVAL_236 <= _EVAL_14;
    end
    if (_EVAL_206) begin
      _EVAL_246 <= _EVAL_12;
    end
    if (_EVAL_2) begin
      _EVAL_258 <= 1'h0;
    end else if (_EVAL_66) begin
      if (_EVAL_83) begin
        _EVAL_258 <= 1'h0;
      end else begin
        _EVAL_258 <= _EVAL_247;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96ad3069)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38f03c62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ae9dd8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d81bf4d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3dd3843f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42e0c193)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51ae211)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24bbc611)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(146642d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(778de31f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cb56083)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91cfcf48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a07ebe8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed69e68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72f15626)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca183a51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6ec8c4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5654c69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a96dbfd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f676ca3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(721da699)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_211) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0c3b97b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77c77d38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37690cd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f46e25e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_211) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1fd181d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa9d2834)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb49a010)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4038c66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73fe57e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7637236)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b71d61c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a864f9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f907601)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7199586)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bf5fca2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_16) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e96f39be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(283039c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_16) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f90c35a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2414cee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f219016)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28e99c18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c7639ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e4fc712)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_16) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe687202)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c342aaf8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0eff1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8513e2dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20b0d224)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86bb27eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0b4375a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd93daec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17acafd9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46be8d7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee7f68a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa451766)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c605e64a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3af4071f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb6da62b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(262ac9e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(929e11d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92f89521)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c0189f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_16) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(926bee20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca955536)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5346c246)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c6ed55b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a932772f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2db1630a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d0e6bd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f00354e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_251 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f517400)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
