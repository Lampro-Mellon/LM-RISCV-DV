//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_65(
  output        _EVAL,
  input         _EVAL_0,
  output        _EVAL_1,
  output [29:0] _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  output [3:0]  _EVAL_5,
  output [2:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  output        _EVAL_9,
  output        _EVAL_10,
  output        _EVAL_11,
  output        _EVAL_12,
  output [31:0] _EVAL_13,
  input         _EVAL_14,
  output        _EVAL_15,
  input  [3:0]  _EVAL_16,
  input  [31:0] _EVAL_17,
  output [3:0]  _EVAL_18,
  input  [2:0]  _EVAL_19,
  input         _EVAL_20,
  input  [29:0] _EVAL_21,
  output [2:0]  _EVAL_22,
  input  [3:0]  _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  output [2:0]  _EVAL_26,
  input  [2:0]  _EVAL_27,
  input         _EVAL_28
);
  reg [31:0] _EVAL_29 [0:1];
  reg [31:0] _RAND_0;
  wire [31:0] _EVAL_29__EVAL_30_data;
  wire  _EVAL_29__EVAL_30_addr;
  wire [31:0] _EVAL_29__EVAL_31_data;
  wire  _EVAL_29__EVAL_31_addr;
  wire  _EVAL_29__EVAL_31_mask;
  wire  _EVAL_29__EVAL_31_en;
  reg  _EVAL_32 [0:1];
  reg [31:0] _RAND_1;
  wire  _EVAL_32__EVAL_33_data;
  wire  _EVAL_32__EVAL_33_addr;
  wire  _EVAL_32__EVAL_34_data;
  wire  _EVAL_32__EVAL_34_addr;
  wire  _EVAL_32__EVAL_34_mask;
  wire  _EVAL_32__EVAL_34_en;
  reg [2:0] _EVAL_35 [0:1];
  reg [31:0] _RAND_2;
  wire [2:0] _EVAL_35__EVAL_36_data;
  wire  _EVAL_35__EVAL_36_addr;
  wire [2:0] _EVAL_35__EVAL_37_data;
  wire  _EVAL_35__EVAL_37_addr;
  wire  _EVAL_35__EVAL_37_mask;
  wire  _EVAL_35__EVAL_37_en;
  reg  _EVAL_38;
  reg [31:0] _RAND_3;
  wire [1:0] _EVAL_39;
  wire [1:0] _EVAL_40;
  wire  _EVAL_41;
  reg [2:0] _EVAL_42 [0:1];
  reg [31:0] _RAND_4;
  wire [2:0] _EVAL_42__EVAL_43_data;
  wire  _EVAL_42__EVAL_43_addr;
  wire [2:0] _EVAL_42__EVAL_44_data;
  wire  _EVAL_42__EVAL_44_addr;
  wire  _EVAL_42__EVAL_44_mask;
  wire  _EVAL_42__EVAL_44_en;
  wire  _EVAL_45;
  wire  _EVAL_46;
  reg  _EVAL_47;
  reg [31:0] _RAND_5;
  reg  _EVAL_49;
  reg [31:0] _RAND_6;
  wire  _EVAL_50;
  reg [2:0] _EVAL_51 [0:1];
  reg [31:0] _RAND_7;
  wire [2:0] _EVAL_51__EVAL_52_data;
  wire  _EVAL_51__EVAL_52_addr;
  wire [2:0] _EVAL_51__EVAL_53_data;
  wire  _EVAL_51__EVAL_53_addr;
  wire  _EVAL_51__EVAL_53_mask;
  wire  _EVAL_51__EVAL_53_en;
  reg  _EVAL_54 [0:1];
  reg [31:0] _RAND_8;
  wire  _EVAL_54__EVAL_55_data;
  wire  _EVAL_54__EVAL_55_addr;
  wire  _EVAL_54__EVAL_56_data;
  wire  _EVAL_54__EVAL_56_addr;
  wire  _EVAL_54__EVAL_56_mask;
  wire  _EVAL_54__EVAL_56_en;
  reg [3:0] _EVAL_57 [0:1];
  reg [31:0] _RAND_9;
  wire [3:0] _EVAL_57__EVAL_58_data;
  wire  _EVAL_57__EVAL_58_addr;
  wire [3:0] _EVAL_57__EVAL_59_data;
  wire  _EVAL_57__EVAL_59_addr;
  wire  _EVAL_57__EVAL_59_mask;
  wire  _EVAL_57__EVAL_59_en;
  reg [3:0] _EVAL_60 [0:1];
  reg [31:0] _RAND_10;
  wire [3:0] _EVAL_60__EVAL_61_data;
  wire  _EVAL_60__EVAL_61_addr;
  wire [3:0] _EVAL_60__EVAL_62_data;
  wire  _EVAL_60__EVAL_62_addr;
  wire  _EVAL_60__EVAL_62_mask;
  wire  _EVAL_60__EVAL_62_en;
  wire  _EVAL_63;
  reg  _EVAL_64 [0:1];
  reg [31:0] _RAND_11;
  wire  _EVAL_64__EVAL_65_data;
  wire  _EVAL_64__EVAL_65_addr;
  wire  _EVAL_64__EVAL_66_data;
  wire  _EVAL_64__EVAL_66_addr;
  wire  _EVAL_64__EVAL_66_mask;
  wire  _EVAL_64__EVAL_66_en;
  reg  _EVAL_68 [0:1];
  reg [31:0] _RAND_12;
  wire  _EVAL_68__EVAL_69_data;
  wire  _EVAL_68__EVAL_69_addr;
  wire  _EVAL_68__EVAL_70_data;
  wire  _EVAL_68__EVAL_70_addr;
  wire  _EVAL_68__EVAL_70_mask;
  wire  _EVAL_68__EVAL_70_en;
  reg [29:0] _EVAL_72 [0:1];
  reg [31:0] _RAND_13;
  wire [29:0] _EVAL_72__EVAL_73_data;
  wire  _EVAL_72__EVAL_73_addr;
  wire [29:0] _EVAL_72__EVAL_74_data;
  wire  _EVAL_72__EVAL_74_addr;
  wire  _EVAL_72__EVAL_74_mask;
  wire  _EVAL_72__EVAL_74_en;
  wire  _EVAL_75;
  wire  _EVAL_76;
  reg  _EVAL_77 [0:1];
  reg [31:0] _RAND_14;
  wire  _EVAL_77__EVAL_78_data;
  wire  _EVAL_77__EVAL_78_addr;
  wire  _EVAL_77__EVAL_79_data;
  wire  _EVAL_77__EVAL_79_addr;
  wire  _EVAL_77__EVAL_79_mask;
  wire  _EVAL_77__EVAL_79_en;
  wire  _EVAL_80;
  wire  _EVAL_81;
  assign _EVAL_29__EVAL_30_addr = _EVAL_49;
  assign _EVAL_29__EVAL_30_data = _EVAL_29[_EVAL_29__EVAL_30_addr];
  assign _EVAL_29__EVAL_31_data = _EVAL_17;
  assign _EVAL_29__EVAL_31_addr = _EVAL_47;
  assign _EVAL_29__EVAL_31_mask = 1'h1;
  assign _EVAL_29__EVAL_31_en = _EVAL_11 & _EVAL_8;
  assign _EVAL_32__EVAL_33_addr = _EVAL_49;
  assign _EVAL_32__EVAL_33_data = _EVAL_32[_EVAL_32__EVAL_33_addr];
  assign _EVAL_32__EVAL_34_data = _EVAL_24;
  assign _EVAL_32__EVAL_34_addr = _EVAL_47;
  assign _EVAL_32__EVAL_34_mask = 1'h1;
  assign _EVAL_32__EVAL_34_en = _EVAL_11 & _EVAL_8;
  assign _EVAL_35__EVAL_36_addr = _EVAL_49;
  assign _EVAL_35__EVAL_36_data = _EVAL_35[_EVAL_35__EVAL_36_addr];
  assign _EVAL_35__EVAL_37_data = _EVAL_3;
  assign _EVAL_35__EVAL_37_addr = _EVAL_47;
  assign _EVAL_35__EVAL_37_mask = 1'h1;
  assign _EVAL_35__EVAL_37_en = _EVAL_11 & _EVAL_8;
  assign _EVAL_42__EVAL_43_addr = _EVAL_49;
  assign _EVAL_42__EVAL_43_data = _EVAL_42[_EVAL_42__EVAL_43_addr];
  assign _EVAL_42__EVAL_44_data = _EVAL_27;
  assign _EVAL_42__EVAL_44_addr = _EVAL_47;
  assign _EVAL_42__EVAL_44_mask = 1'h1;
  assign _EVAL_42__EVAL_44_en = _EVAL_11 & _EVAL_8;
  assign _EVAL_51__EVAL_52_addr = _EVAL_49;
  assign _EVAL_51__EVAL_52_data = _EVAL_51[_EVAL_51__EVAL_52_addr];
  assign _EVAL_51__EVAL_53_data = _EVAL_19;
  assign _EVAL_51__EVAL_53_addr = _EVAL_47;
  assign _EVAL_51__EVAL_53_mask = 1'h1;
  assign _EVAL_51__EVAL_53_en = _EVAL_11 & _EVAL_8;
  assign _EVAL_54__EVAL_55_addr = _EVAL_49;
  assign _EVAL_54__EVAL_55_data = _EVAL_54[_EVAL_54__EVAL_55_addr];
  assign _EVAL_54__EVAL_56_data = _EVAL_20;
  assign _EVAL_54__EVAL_56_addr = _EVAL_47;
  assign _EVAL_54__EVAL_56_mask = 1'h1;
  assign _EVAL_54__EVAL_56_en = _EVAL_11 & _EVAL_8;
  assign _EVAL_57__EVAL_58_addr = _EVAL_49;
  assign _EVAL_57__EVAL_58_data = _EVAL_57[_EVAL_57__EVAL_58_addr];
  assign _EVAL_57__EVAL_59_data = _EVAL_16;
  assign _EVAL_57__EVAL_59_addr = _EVAL_47;
  assign _EVAL_57__EVAL_59_mask = 1'h1;
  assign _EVAL_57__EVAL_59_en = _EVAL_11 & _EVAL_8;
  assign _EVAL_60__EVAL_61_addr = _EVAL_49;
  assign _EVAL_60__EVAL_61_data = _EVAL_60[_EVAL_60__EVAL_61_addr];
  assign _EVAL_60__EVAL_62_data = _EVAL_23;
  assign _EVAL_60__EVAL_62_addr = _EVAL_47;
  assign _EVAL_60__EVAL_62_mask = 1'h1;
  assign _EVAL_60__EVAL_62_en = _EVAL_11 & _EVAL_8;
  assign _EVAL_64__EVAL_65_addr = _EVAL_49;
  assign _EVAL_64__EVAL_65_data = _EVAL_64[_EVAL_64__EVAL_65_addr];
  assign _EVAL_64__EVAL_66_data = _EVAL_4;
  assign _EVAL_64__EVAL_66_addr = _EVAL_47;
  assign _EVAL_64__EVAL_66_mask = 1'h1;
  assign _EVAL_64__EVAL_66_en = _EVAL_11 & _EVAL_8;
  assign _EVAL_68__EVAL_69_addr = _EVAL_49;
  assign _EVAL_68__EVAL_69_data = _EVAL_68[_EVAL_68__EVAL_69_addr];
  assign _EVAL_68__EVAL_70_data = _EVAL_0;
  assign _EVAL_68__EVAL_70_addr = _EVAL_47;
  assign _EVAL_68__EVAL_70_mask = 1'h1;
  assign _EVAL_68__EVAL_70_en = _EVAL_11 & _EVAL_8;
  assign _EVAL_72__EVAL_73_addr = _EVAL_49;
  assign _EVAL_72__EVAL_73_data = _EVAL_72[_EVAL_72__EVAL_73_addr];
  assign _EVAL_72__EVAL_74_data = _EVAL_21;
  assign _EVAL_72__EVAL_74_addr = _EVAL_47;
  assign _EVAL_72__EVAL_74_mask = 1'h1;
  assign _EVAL_72__EVAL_74_en = _EVAL_11 & _EVAL_8;
  assign _EVAL_77__EVAL_78_addr = _EVAL_49;
  assign _EVAL_77__EVAL_78_data = _EVAL_77[_EVAL_77__EVAL_78_addr];
  assign _EVAL_77__EVAL_79_data = _EVAL_28;
  assign _EVAL_77__EVAL_79_addr = _EVAL_47;
  assign _EVAL_77__EVAL_79_mask = 1'h1;
  assign _EVAL_77__EVAL_79_en = _EVAL_11 & _EVAL_8;
  assign _EVAL_9 = _EVAL_32__EVAL_33_data;
  assign _EVAL = _EVAL_77__EVAL_78_data;
  assign _EVAL_11 = ~_EVAL_63;
  assign _EVAL_63 = _EVAL_81 & _EVAL_38;
  assign _EVAL_12 = ~_EVAL_50;
  assign _EVAL_50 = _EVAL_81 & _EVAL_41;
  assign _EVAL_13 = _EVAL_29__EVAL_30_data;
  assign _EVAL_15 = _EVAL_64__EVAL_65_data;
  assign _EVAL_45 = _EVAL_25 & _EVAL_12;
  assign _EVAL_80 = _EVAL_40[0];
  assign _EVAL_46 = _EVAL_11 & _EVAL_8;
  assign _EVAL_10 = _EVAL_68__EVAL_69_data;
  assign _EVAL_76 = _EVAL_39[0];
  assign _EVAL_75 = _EVAL_46 != _EVAL_45;
  assign _EVAL_41 = ~_EVAL_38;
  assign _EVAL_6 = _EVAL_42__EVAL_43_data;
  assign _EVAL_18 = _EVAL_60__EVAL_61_data;
  assign _EVAL_26 = _EVAL_35__EVAL_36_data;
  assign _EVAL_1 = _EVAL_54__EVAL_55_data;
  assign _EVAL_40 = _EVAL_47 + 1'h1;
  assign _EVAL_5 = _EVAL_57__EVAL_58_data;
  assign _EVAL_81 = _EVAL_47 == _EVAL_49;
  assign _EVAL_22 = _EVAL_51__EVAL_52_data;
  assign _EVAL_2 = _EVAL_72__EVAL_73_data;
  assign _EVAL_39 = _EVAL_49 + 1'h1;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_29[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_32[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_35[initvar] = _RAND_2[2:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_38 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_42[initvar] = _RAND_4[2:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_47 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_49 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_51[initvar] = _RAND_7[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_54[initvar] = _RAND_8[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_57[initvar] = _RAND_9[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_60[initvar] = _RAND_10[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_11 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_64[initvar] = _RAND_11[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_68[initvar] = _RAND_12[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_13 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_72[initvar] = _RAND_13[29:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_14 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_77[initvar] = _RAND_14[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_14) begin
    if(_EVAL_29__EVAL_31_en & _EVAL_29__EVAL_31_mask) begin
      _EVAL_29[_EVAL_29__EVAL_31_addr] <= _EVAL_29__EVAL_31_data;
    end
    if(_EVAL_32__EVAL_34_en & _EVAL_32__EVAL_34_mask) begin
      _EVAL_32[_EVAL_32__EVAL_34_addr] <= _EVAL_32__EVAL_34_data;
    end
    if(_EVAL_35__EVAL_37_en & _EVAL_35__EVAL_37_mask) begin
      _EVAL_35[_EVAL_35__EVAL_37_addr] <= _EVAL_35__EVAL_37_data;
    end
    if (_EVAL_7) begin
      _EVAL_38 <= 1'h0;
    end else if (_EVAL_75) begin
      _EVAL_38 <= _EVAL_46;
    end
    if(_EVAL_42__EVAL_44_en & _EVAL_42__EVAL_44_mask) begin
      _EVAL_42[_EVAL_42__EVAL_44_addr] <= _EVAL_42__EVAL_44_data;
    end
    if (_EVAL_7) begin
      _EVAL_47 <= 1'h0;
    end else if (_EVAL_46) begin
      _EVAL_47 <= _EVAL_80;
    end
    if (_EVAL_7) begin
      _EVAL_49 <= 1'h0;
    end else if (_EVAL_45) begin
      _EVAL_49 <= _EVAL_76;
    end
    if(_EVAL_51__EVAL_53_en & _EVAL_51__EVAL_53_mask) begin
      _EVAL_51[_EVAL_51__EVAL_53_addr] <= _EVAL_51__EVAL_53_data;
    end
    if(_EVAL_54__EVAL_56_en & _EVAL_54__EVAL_56_mask) begin
      _EVAL_54[_EVAL_54__EVAL_56_addr] <= _EVAL_54__EVAL_56_data;
    end
    if(_EVAL_57__EVAL_59_en & _EVAL_57__EVAL_59_mask) begin
      _EVAL_57[_EVAL_57__EVAL_59_addr] <= _EVAL_57__EVAL_59_data;
    end
    if(_EVAL_60__EVAL_62_en & _EVAL_60__EVAL_62_mask) begin
      _EVAL_60[_EVAL_60__EVAL_62_addr] <= _EVAL_60__EVAL_62_data;
    end
    if(_EVAL_64__EVAL_66_en & _EVAL_64__EVAL_66_mask) begin
      _EVAL_64[_EVAL_64__EVAL_66_addr] <= _EVAL_64__EVAL_66_data;
    end
    if(_EVAL_68__EVAL_70_en & _EVAL_68__EVAL_70_mask) begin
      _EVAL_68[_EVAL_68__EVAL_70_addr] <= _EVAL_68__EVAL_70_data;
    end
    if(_EVAL_72__EVAL_74_en & _EVAL_72__EVAL_74_mask) begin
      _EVAL_72[_EVAL_72__EVAL_74_addr] <= _EVAL_72__EVAL_74_data;
    end
    if(_EVAL_77__EVAL_79_en & _EVAL_77__EVAL_79_mask) begin
      _EVAL_77[_EVAL_77__EVAL_79_addr] <= _EVAL_77__EVAL_79_data;
    end
  end
endmodule
