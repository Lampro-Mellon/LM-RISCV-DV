//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_32(
  output        _EVAL,
  input  [2:0]  _EVAL_0,
  output        _EVAL_1,
  input  [31:0] _EVAL_2,
  input  [2:0]  _EVAL_3,
  output        _EVAL_4,
  input  [3:0]  _EVAL_5,
  output        _EVAL_6,
  output [3:0]  _EVAL_7,
  input         _EVAL_8,
  output        _EVAL_9,
  input         _EVAL_10,
  output [2:0]  _EVAL_11,
  input  [3:0]  _EVAL_12,
  output        _EVAL_13,
  output [2:0]  _EVAL_14,
  input         _EVAL_15,
  output [1:0]  _EVAL_16,
  output        _EVAL_17,
  input  [2:0]  _EVAL_18,
  output [31:0] _EVAL_19,
  input         _EVAL_20,
  output        _EVAL_21,
  input         _EVAL_22,
  output        _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input  [3:0]  _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input  [2:0]  _EVAL_32,
  output        _EVAL_33,
  input  [29:0] _EVAL_34,
  input  [31:0] _EVAL_35,
  output [29:0] _EVAL_36,
  output        _EVAL_37,
  output        _EVAL_38,
  output [2:0]  _EVAL_39,
  input         _EVAL_40,
  input  [2:0]  _EVAL_41,
  input         _EVAL_42,
  input         _EVAL_43,
  output [3:0]  _EVAL_44,
  output        _EVAL_45,
  input         _EVAL_46,
  output        _EVAL_47,
  output [31:0] _EVAL_48,
  input  [1:0]  _EVAL_49,
  output [2:0]  _EVAL_50,
  output [3:0]  _EVAL_51,
  input         _EVAL_52,
  output [2:0]  _EVAL_53,
  output        _EVAL_54
);
  assign _EVAL_45 = _EVAL_15;
  assign _EVAL_7 = _EVAL_12;
  assign _EVAL_44 = _EVAL_5;
  assign _EVAL_13 = _EVAL_42;
  assign _EVAL_17 = _EVAL_26;
  assign _EVAL_50 = _EVAL_32;
  assign _EVAL_19 = _EVAL_2;
  assign _EVAL_47 = _EVAL_8;
  assign _EVAL = _EVAL_46;
  assign _EVAL_33 = _EVAL_22;
  assign _EVAL_21 = _EVAL_52;
  assign _EVAL_48 = _EVAL_35;
  assign _EVAL_4 = _EVAL_40;
  assign _EVAL_11 = _EVAL_41;
  assign _EVAL_16 = _EVAL_49;
  assign _EVAL_14 = _EVAL_3;
  assign _EVAL_39 = _EVAL_0;
  assign _EVAL_54 = _EVAL_24;
  assign _EVAL_1 = _EVAL_10;
  assign _EVAL_38 = _EVAL_27;
  assign _EVAL_36 = _EVAL_34;
  assign _EVAL_9 = _EVAL_29;
  assign _EVAL_53 = _EVAL_18;
  assign _EVAL_6 = _EVAL_43;
  assign _EVAL_51 = _EVAL_28;
  assign _EVAL_23 = _EVAL_31;
  assign _EVAL_37 = _EVAL_20;
endmodule
