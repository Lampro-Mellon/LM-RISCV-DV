//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_119(
  input         _EVAL,
  input  [6:0]  _EVAL_0,
  input         _EVAL_1,
  output        _EVAL_2,
  input  [31:0] _EVAL_3,
  input         _EVAL_4,
  output [1:0]  _EVAL_5,
  output [2:0]  _EVAL_6,
  output [31:0] _EVAL_7,
  output        _EVAL_8,
  input         _EVAL_9,
  input  [31:0] _EVAL_10,
  output        _EVAL_11,
  input         _EVAL_12,
  output [31:0] _EVAL_13,
  output [3:0]  _EVAL_14,
  input         _EVAL_15,
  output        _EVAL_16,
  output [8:0]  _EVAL_17,
  input  [1:0]  _EVAL_18
);
  wire  _EVAL_19;
  wire [3:0] _EVAL_20;
  wire [8:0] _EVAL_21;
  wire [8:0] _EVAL_22;
  wire [2:0] _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  assign _EVAL_5 = {{1'd0}, _EVAL_25};
  assign _EVAL_19 = _EVAL_18 == 2'h1;
  assign _EVAL_2 = _EVAL_15;
  assign _EVAL_13 = _EVAL_24 ? _EVAL_3 : 32'h0;
  assign _EVAL_25 = _EVAL | _EVAL_1;
  assign _EVAL_20 = _EVAL_19 ? 4'hf : 4'h0;
  assign _EVAL_16 = _EVAL_4;
  assign _EVAL_8 = _EVAL_12;
  assign _EVAL_7 = _EVAL_10;
  assign _EVAL_22 = {_EVAL_0, 2'h0};
  assign _EVAL_24 = _EVAL_18 == 2'h2;
  assign _EVAL_23 = _EVAL_19 ? 3'h4 : 3'h1;
  assign _EVAL_6 = _EVAL_24 ? 3'h0 : _EVAL_23;
  assign _EVAL_14 = _EVAL_24 ? 4'hf : _EVAL_20;
  assign _EVAL_11 = _EVAL_9;
  assign _EVAL_17 = _EVAL_24 ? _EVAL_22 : _EVAL_21;
  assign _EVAL_21 = _EVAL_19 ? _EVAL_22 : 9'h40;
endmodule
