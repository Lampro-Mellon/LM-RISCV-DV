//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_19(
  input  [3:0]  _EVAL,
  output [2:0]  _EVAL_0,
  output        _EVAL_1,
  output [31:0] _EVAL_2,
  input         _EVAL_3,
  output        _EVAL_4,
  input  [31:0] _EVAL_5,
  output [1:0]  _EVAL_6,
  output [31:0] _EVAL_7,
  input  [31:0] _EVAL_8,
  output [2:0]  _EVAL_9,
  output        _EVAL_10,
  output [2:0]  _EVAL_11,
  input         _EVAL_12,
  input  [2:0]  _EVAL_13,
  input  [2:0]  _EVAL_14,
  input  [1:0]  _EVAL_15,
  output [2:0]  _EVAL_16,
  output [3:0]  _EVAL_17,
  output [31:0] _EVAL_18,
  output [2:0]  _EVAL_19,
  input         _EVAL_20,
  input         _EVAL_21,
  output        _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  output [1:0]  _EVAL_25,
  output        _EVAL_26,
  input         _EVAL_27,
  input  [2:0]  _EVAL_28,
  input  [31:0] _EVAL_29,
  input  [2:0]  _EVAL_30,
  input  [1:0]  _EVAL_31,
  input  [2:0]  _EVAL_32
);
  wire [2:0] buffer__EVAL;
  wire [2:0] buffer__EVAL_0;
  wire [31:0] buffer__EVAL_1;
  wire  buffer__EVAL_2;
  wire  buffer__EVAL_3;
  wire  buffer__EVAL_4;
  wire [31:0] buffer__EVAL_5;
  wire [3:0] buffer__EVAL_6;
  wire  buffer__EVAL_7;
  wire [2:0] buffer__EVAL_8;
  wire [31:0] buffer__EVAL_9;
  wire  buffer__EVAL_10;
  wire [31:0] buffer__EVAL_11;
  wire [2:0] buffer__EVAL_12;
  wire [2:0] buffer__EVAL_13;
  wire [3:0] buffer__EVAL_14;
  wire [1:0] buffer__EVAL_15;
  wire  buffer__EVAL_16;
  wire [2:0] buffer__EVAL_17;
  wire [2:0] buffer__EVAL_18;
  wire [31:0] buffer__EVAL_19;
  wire [1:0] buffer__EVAL_20;
  wire [2:0] buffer__EVAL_21;
  wire  buffer__EVAL_22;
  wire [1:0] buffer__EVAL_23;
  wire [31:0] buffer__EVAL_24;
  wire [2:0] buffer__EVAL_25;
  wire  buffer__EVAL_26;
  wire  buffer__EVAL_27;
  wire [2:0] buffer__EVAL_28;
  wire  buffer__EVAL_29;
  wire [1:0] buffer__EVAL_30;
  wire  buffer__EVAL_31;
  wire  buffer__EVAL_32;
  wire [1:0] fragmenter__EVAL;
  wire [31:0] fragmenter__EVAL_0;
  wire [1:0] fragmenter__EVAL_1;
  wire  fragmenter__EVAL_2;
  wire [1:0] fragmenter__EVAL_3;
  wire  fragmenter__EVAL_4;
  wire [2:0] fragmenter__EVAL_5;
  wire [2:0] fragmenter__EVAL_6;
  wire [2:0] fragmenter__EVAL_7;
  wire  fragmenter__EVAL_8;
  wire [3:0] fragmenter__EVAL_9;
  wire [2:0] fragmenter__EVAL_10;
  wire  fragmenter__EVAL_11;
  wire [2:0] fragmenter__EVAL_12;
  wire [2:0] fragmenter__EVAL_13;
  wire [31:0] fragmenter__EVAL_14;
  wire  fragmenter__EVAL_15;
  wire  fragmenter__EVAL_16;
  wire [31:0] fragmenter__EVAL_17;
  wire  fragmenter__EVAL_18;
  wire  fragmenter__EVAL_19;
  wire  fragmenter__EVAL_20;
  wire [2:0] fragmenter__EVAL_21;
  wire  fragmenter__EVAL_22;
  wire [2:0] fragmenter__EVAL_23;
  wire [1:0] fragmenter__EVAL_24;
  wire [2:0] fragmenter__EVAL_25;
  wire [31:0] fragmenter__EVAL_26;
  wire [2:0] fragmenter__EVAL_27;
  wire [31:0] fragmenter__EVAL_28;
  wire  fragmenter__EVAL_29;
  wire  fragmenter__EVAL_30;
  wire [3:0] fragmenter__EVAL_31;
  wire [31:0] fragmenter__EVAL_32;
  _EVAL_18 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32)
  );
  _EVAL_16 fragmenter (
    ._EVAL(fragmenter__EVAL),
    ._EVAL_0(fragmenter__EVAL_0),
    ._EVAL_1(fragmenter__EVAL_1),
    ._EVAL_2(fragmenter__EVAL_2),
    ._EVAL_3(fragmenter__EVAL_3),
    ._EVAL_4(fragmenter__EVAL_4),
    ._EVAL_5(fragmenter__EVAL_5),
    ._EVAL_6(fragmenter__EVAL_6),
    ._EVAL_7(fragmenter__EVAL_7),
    ._EVAL_8(fragmenter__EVAL_8),
    ._EVAL_9(fragmenter__EVAL_9),
    ._EVAL_10(fragmenter__EVAL_10),
    ._EVAL_11(fragmenter__EVAL_11),
    ._EVAL_12(fragmenter__EVAL_12),
    ._EVAL_13(fragmenter__EVAL_13),
    ._EVAL_14(fragmenter__EVAL_14),
    ._EVAL_15(fragmenter__EVAL_15),
    ._EVAL_16(fragmenter__EVAL_16),
    ._EVAL_17(fragmenter__EVAL_17),
    ._EVAL_18(fragmenter__EVAL_18),
    ._EVAL_19(fragmenter__EVAL_19),
    ._EVAL_20(fragmenter__EVAL_20),
    ._EVAL_21(fragmenter__EVAL_21),
    ._EVAL_22(fragmenter__EVAL_22),
    ._EVAL_23(fragmenter__EVAL_23),
    ._EVAL_24(fragmenter__EVAL_24),
    ._EVAL_25(fragmenter__EVAL_25),
    ._EVAL_26(fragmenter__EVAL_26),
    ._EVAL_27(fragmenter__EVAL_27),
    ._EVAL_28(fragmenter__EVAL_28),
    ._EVAL_29(fragmenter__EVAL_29),
    ._EVAL_30(fragmenter__EVAL_30),
    ._EVAL_31(fragmenter__EVAL_31),
    ._EVAL_32(fragmenter__EVAL_32)
  );
  assign buffer__EVAL_4 = _EVAL_27;
  assign _EVAL_22 = fragmenter__EVAL_8;
  assign _EVAL_10 = fragmenter__EVAL_29;
  assign buffer__EVAL_6 = _EVAL;
  assign _EVAL_6 = fragmenter__EVAL_24;
  assign fragmenter__EVAL_28 = buffer__EVAL_5;
  assign fragmenter__EVAL_20 = _EVAL_20;
  assign fragmenter__EVAL_0 = _EVAL_29;
  assign _EVAL_11 = buffer__EVAL_12;
  assign fragmenter__EVAL = buffer__EVAL_23;
  assign _EVAL_1 = buffer__EVAL_3;
  assign buffer__EVAL_13 = _EVAL_30;
  assign _EVAL_0 = fragmenter__EVAL_23;
  assign buffer__EVAL_11 = fragmenter__EVAL_14;
  assign fragmenter__EVAL_2 = buffer__EVAL_7;
  assign fragmenter__EVAL_6 = buffer__EVAL_17;
  assign buffer__EVAL_27 = _EVAL_12;
  assign fragmenter__EVAL_11 = _EVAL_24;
  assign _EVAL_18 = fragmenter__EVAL_26;
  assign fragmenter__EVAL_18 = buffer__EVAL_22;
  assign _EVAL_9 = buffer__EVAL_21;
  assign buffer__EVAL_26 = fragmenter__EVAL_16;
  assign fragmenter__EVAL_15 = buffer__EVAL_2;
  assign buffer__EVAL_9 = _EVAL_5;
  assign fragmenter__EVAL_19 = _EVAL_12;
  assign _EVAL_16 = fragmenter__EVAL_5;
  assign buffer__EVAL_8 = _EVAL_14;
  assign fragmenter__EVAL_22 = _EVAL_21;
  assign _EVAL_4 = buffer__EVAL_32;
  assign buffer__EVAL_19 = _EVAL_8;
  assign fragmenter__EVAL_1 = _EVAL_31;
  assign fragmenter__EVAL_27 = buffer__EVAL_25;
  assign buffer__EVAL_10 = _EVAL_3;
  assign _EVAL_19 = fragmenter__EVAL_25;
  assign _EVAL_17 = fragmenter__EVAL_31;
  assign buffer__EVAL_30 = fragmenter__EVAL_3;
  assign _EVAL_25 = buffer__EVAL_15;
  assign buffer__EVAL_20 = _EVAL_15;
  assign fragmenter__EVAL_9 = buffer__EVAL_14;
  assign _EVAL_2 = fragmenter__EVAL_32;
  assign fragmenter__EVAL_21 = _EVAL_28;
  assign buffer__EVAL_29 = fragmenter__EVAL_30;
  assign _EVAL_7 = buffer__EVAL_1;
  assign buffer__EVAL_31 = _EVAL_23;
  assign buffer__EVAL_16 = _EVAL_24;
  assign buffer__EVAL_28 = fragmenter__EVAL_12;
  assign fragmenter__EVAL_7 = buffer__EVAL;
  assign fragmenter__EVAL_13 = _EVAL_13;
  assign buffer__EVAL_0 = fragmenter__EVAL_10;
  assign fragmenter__EVAL_17 = buffer__EVAL_24;
  assign _EVAL_26 = fragmenter__EVAL_4;
  assign buffer__EVAL_18 = _EVAL_32;
endmodule
