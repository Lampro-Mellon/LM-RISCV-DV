//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_62_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [3:0]  _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [3:0]  _EVAL_11,
  input  [3:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input  [1:0]  _EVAL_16,
  input         _EVAL_17,
  input  [29:0] _EVAL_18
);
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire [32:0] _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  reg [2:0] _EVAL_31;
  reg [31:0] _RAND_0;
  wire [4:0] _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire [7:0] _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire [3:0] _EVAL_49;
  wire  _EVAL_50;
  wire [31:0] _EVAL_51;
  wire [6:0] _EVAL_52;
  wire [7:0] _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire [30:0] _EVAL_61;
  wire  _EVAL_62;
  reg [3:0] _EVAL_63;
  reg [31:0] _RAND_1;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire [4:0] _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire [22:0] _EVAL_71;
  wire  _EVAL_72;
  wire [3:0] _EVAL_73;
  wire  _EVAL_75;
  wire  _EVAL_76;
  reg [2:0] _EVAL_77;
  reg [31:0] _RAND_2;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_80;
  wire [4:0] _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire [1:0] _EVAL_95;
  wire [1:0] _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire [30:0] _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire [5:0] _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire [30:0] _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire [4:0] _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire [30:0] _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire [7:0] _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire [5:0] _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  reg [1:0] _EVAL_142;
  reg [31:0] _RAND_3;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire [7:0] _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire [5:0] _EVAL_155;
  wire [30:0] _EVAL_156;
  wire  _EVAL_157;
  wire [30:0] _EVAL_158;
  wire [6:0] _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire [30:0] _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  reg [2:0] _EVAL_168;
  reg [31:0] _RAND_4;
  reg [3:0] _EVAL_169;
  reg [31:0] _RAND_5;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  reg  _EVAL_176;
  reg [31:0] _RAND_6;
  reg [31:0] _EVAL_177;
  reg [31:0] _RAND_7;
  wire  _EVAL_178;
  wire [4:0] _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire [6:0] _EVAL_187;
  wire  _EVAL_188;
  wire [30:0] _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire [7:0] _EVAL_196;
  wire  _EVAL_197;
  wire [3:0] _EVAL_198;
  wire  _EVAL_199;
  wire [7:0] _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire [29:0] _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire [7:0] _EVAL_216;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  reg [4:0] _EVAL_224;
  reg [31:0] _RAND_8;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire [29:0] _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire [6:0] _EVAL_235;
  wire [22:0] _EVAL_236;
  wire [7:0] _EVAL_237;
  wire  _EVAL_238;
  wire [4:0] _EVAL_239;
  wire  _EVAL_240;
  reg [2:0] _EVAL_241;
  reg [31:0] _RAND_9;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  reg [2:0] _EVAL_247;
  reg [31:0] _RAND_10;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire [4:0] _EVAL_253;
  wire [5:0] _EVAL_254;
  wire  _EVAL_255;
  wire [30:0] _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire [3:0] _EVAL_260;
  wire [29:0] _EVAL_261;
  wire  _EVAL_262;
  reg [5:0] _EVAL_263;
  reg [31:0] _RAND_11;
  reg [29:0] _EVAL_264;
  reg [31:0] _RAND_12;
  wire  _EVAL_265;
  reg [5:0] _EVAL_266;
  reg [31:0] _RAND_13;
  wire [30:0] _EVAL_267;
  wire [29:0] _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire [4:0] _EVAL_276;
  wire [5:0] _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  reg [5:0] _EVAL_283;
  reg [31:0] _RAND_14;
  wire  _EVAL_284;
  wire [30:0] _EVAL_285;
  wire  _EVAL_286;
  wire [5:0] _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire [1:0] _EVAL_293;
  wire  _EVAL_294;
  reg  _EVAL_295;
  reg [31:0] _RAND_15;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire [29:0] _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  reg [5:0] _EVAL_308;
  reg [31:0] _RAND_16;
  wire [1:0] _EVAL_310;
  wire  _EVAL_311;
  wire [30:0] _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_36 = _EVAL_87 | _EVAL_230;
  assign _EVAL_95 = 2'h1 << _EVAL_64;
  assign _EVAL_73 = ~_EVAL_12;
  assign _EVAL_27 = _EVAL_9 == 3'h2;
  assign _EVAL_109 = ~_EVAL_5;
  assign _EVAL_78 = ~_EVAL_116;
  assign _EVAL_84 = _EVAL_70 & _EVAL_292;
  assign _EVAL_136 = _EVAL_128[7:2];
  assign _EVAL_207 = _EVAL_302 | _EVAL_15;
  assign _EVAL_60 = _EVAL_313 & _EVAL_288;
  assign _EVAL_271 = _EVAL_10 <= 3'h2;
  assign _EVAL_205 = _EVAL_273 & _EVAL_41;
  assign _EVAL_313 = _EVAL_2 <= 4'h8;
  assign _EVAL_261 = _EVAL_18 ^ 30'h20000000;
  assign _EVAL_141 = plusarg_reader_out == 32'h0;
  assign _EVAL_249 = _EVAL_1 == _EVAL_247;
  assign _EVAL_251 = _EVAL_4 == 3'h6;
  assign _EVAL_310 = _EVAL_95 | 2'h1;
  assign _EVAL_191 = _EVAL_160 | _EVAL_15;
  assign _EVAL_33 = _EVAL_0 == _EVAL_241;
  assign _EVAL_234 = _EVAL_293 == 2'h1;
  assign _EVAL_282 = _EVAL_8 & _EVAL_57;
  assign _EVAL_143 = _EVAL_226 & _EVAL_79;
  assign _EVAL_119 = ~_EVAL_98;
  assign _EVAL_194 = _EVAL_9 == 3'h4;
  assign _EVAL_149 = _EVAL_199 & _EVAL_97;
  assign _EVAL_97 = _EVAL_273 & _EVAL_68;
  assign _EVAL_230 = _EVAL_115 & _EVAL_273;
  assign _EVAL_98 = _EVAL_146 | _EVAL_15;
  assign _EVAL_115 = _EVAL_310[1];
  assign _EVAL_268 = _EVAL_18 ^ 30'h2000000;
  assign _EVAL_162 = $signed(_EVAL_158) & -31'sh1000;
  assign _EVAL_32 = _EVAL_200[4:0];
  assign _EVAL_88 = _EVAL_91 | _EVAL_15;
  assign _EVAL_213 = _EVAL_9 == 3'h6;
  assign _EVAL_44 = 8'h1 << _EVAL_1;
  assign _EVAL_103 = _EVAL_292 | _EVAL_135;
  assign _EVAL_66 = ~_EVAL_102;
  assign _EVAL_300 = _EVAL_18 & _EVAL_204;
  assign _EVAL_211 = ~_EVAL_21;
  assign _EVAL_100 = _EVAL_61;
  assign _EVAL_212 = ~_EVAL_273;
  assign _EVAL_185 = _EVAL_87 | _EVAL_131;
  assign _EVAL_101 = _EVAL_234 | _EVAL_39;
  assign _EVAL_262 = _EVAL_9 == 3'h5;
  assign _EVAL_188 = _EVAL_18 == _EVAL_264;
  assign _EVAL_123 = _EVAL & _EVAL_167;
  assign _EVAL_134 = _EVAL_300 == 30'h0;
  assign _EVAL_186 = _EVAL_184 | _EVAL_15;
  assign _EVAL_157 = $signed(_EVAL_125) == 31'sh0;
  assign _EVAL_219 = _EVAL_96 == 2'h0;
  assign _EVAL_126 = $signed(_EVAL_113) == 31'sh0;
  assign _EVAL_294 = _EVAL_1 == 3'h4;
  assign _EVAL_293 = _EVAL_0[2:1];
  assign _EVAL_202 = ~_EVAL_22;
  assign _EVAL_50 = _EVAL_70 & _EVAL_288;
  assign _EVAL_317 = _EVAL_177 < plusarg_reader_out;
  assign _EVAL_62 = _EVAL_199 & _EVAL_205;
  assign _EVAL_298 = _EVAL_35 | _EVAL_15;
  assign _EVAL_22 = _EVAL_270 | _EVAL_15;
  assign _EVAL_43 = _EVAL_16 != 2'h2;
  assign _EVAL_248 = ~_EVAL_207;
  assign _EVAL_92 = ~_EVAL_191;
  assign _EVAL_291 = ~_EVAL_154;
  assign _EVAL_163 = ~_EVAL_299;
  assign _EVAL_304 = _EVAL_5 == _EVAL_295;
  assign _EVAL_70 = _EVAL_2 <= 4'h2;
  assign _EVAL_35 = _EVAL_10 <= 3'h1;
  assign _EVAL_302 = _EVAL_17 == _EVAL_176;
  assign _EVAL_166 = _EVAL_244 & _EVAL_40;
  assign _EVAL_240 = _EVAL_10 == _EVAL_168;
  assign _EVAL_129 = _EVAL_69 | _EVAL_15;
  assign _EVAL_278 = _EVAL_10 == 3'h0;
  assign _EVAL_116 = _EVAL_304 | _EVAL_15;
  assign _EVAL_37 = _EVAL & _EVAL_286;
  assign _EVAL_214 = ~_EVAL_206;
  assign _EVAL_274 = ~_EVAL_93;
  assign _EVAL_192 = _EVAL_249 | _EVAL_15;
  assign _EVAL_259 = _EVAL_185 | _EVAL_173;
  assign _EVAL_48 = _EVAL_29 | _EVAL_141;
  assign _EVAL_19 = _EVAL_212 & _EVAL_68;
  assign _EVAL_131 = _EVAL_115 & _EVAL_212;
  assign _EVAL_299 = _EVAL_80 | _EVAL_15;
  assign _EVAL_206 = _EVAL_164 | _EVAL_15;
  assign _EVAL_297 = ~_EVAL_290;
  assign _EVAL_303 = _EVAL_8 & _EVAL_27;
  assign _EVAL_155 = _EVAL_159[5:0];
  assign _EVAL_244 = _EVAL_13 & _EVAL;
  assign _EVAL_99 = _EVAL & _EVAL_170;
  assign _EVAL_225 = _EVAL_12 == _EVAL_198;
  assign _EVAL_67 = _EVAL_32 | _EVAL_224;
  assign _EVAL_164 = _EVAL_109 | _EVAL_7;
  assign _EVAL_145 = _EVAL_134 | _EVAL_15;
  assign _EVAL_215 = _EVAL_224 != 5'h0;
  assign _EVAL_72 = _EVAL_265 | _EVAL_15;
  assign _EVAL_167 = _EVAL_4 == 3'h0;
  assign _EVAL_139 = _EVAL_11 >= 4'h2;
  assign _EVAL_61 = $signed(_EVAL_156) & -31'sh2000;
  assign _EVAL_199 = _EVAL_310[0];
  assign _EVAL_201 = ~_EVAL_88;
  assign _EVAL_20 = ~_EVAL_315;
  assign _EVAL_46 = ~_EVAL_186;
  assign _EVAL_311 = _EVAL_246 | _EVAL_15;
  assign _EVAL_216 = _EVAL_71[7:0];
  assign _EVAL_87 = _EVAL_2 >= 4'h2;
  assign _EVAL_171 = ~_EVAL_75;
  assign _EVAL_80 = _EVAL_101 | _EVAL_114;
  assign _EVAL_190 = _EVAL_107 | _EVAL_219;
  assign _EVAL_227 = _EVAL_109 | _EVAL_15;
  assign _EVAL_75 = _EVAL_305 | _EVAL_15;
  assign _EVAL_133 = _EVAL_8 & _EVAL_262;
  assign _EVAL_260 = _EVAL_12 & _EVAL_49;
  assign _EVAL_146 = _EVAL_190 | _EVAL_294;
  assign _EVAL_279 = _EVAL_11 == _EVAL_169;
  assign _EVAL_223 = _EVAL_8 & _EVAL_213;
  assign _EVAL_127 = _EVAL_4[0];
  assign _EVAL_314 = ~_EVAL_172;
  assign _EVAL_135 = $signed(_EVAL_100) == 31'sh0;
  assign _EVAL_226 = _EVAL_6 & _EVAL_8;
  assign _EVAL_118 = _EVAL_66 | _EVAL_15;
  assign _EVAL_267 = $signed(_EVAL_285) & -31'sh1000000;
  assign _EVAL_106 = _EVAL_144 | _EVAL_15;
  assign _EVAL_239 = _EVAL_224 >> _EVAL_0;
  assign _EVAL_235 = _EVAL_283 - 6'h1;
  assign _EVAL_170 = _EVAL_4 == 3'h1;
  assign _EVAL_94 = _EVAL_139 | _EVAL_15;
  assign _EVAL_144 = _EVAL_2 == _EVAL_63;
  assign _EVAL_41 = ~_EVAL_68;
  assign _EVAL_57 = _EVAL_9 == 3'h3;
  assign _EVAL_173 = _EVAL_199 & _EVAL_82;
  assign _EVAL_112 = ~_EVAL_250;
  assign _EVAL_153 = _EVAL_9 == 3'h0;
  assign _EVAL_221 = _EVAL_36 | _EVAL_62;
  assign _EVAL_148 = _EVAL_236[7:0];
  assign _EVAL_154 = _EVAL_279 | _EVAL_15;
  assign _EVAL_58 = _EVAL_197 | _EVAL_15;
  assign _EVAL_124 = _EVAL_8 & _EVAL_307;
  assign _EVAL_237 = 8'h1 << _EVAL_0;
  assign _EVAL_183 = ~_EVAL_298;
  assign _EVAL_158 = {1'b0,$signed(_EVAL_232)};
  assign _EVAL_287 = _EVAL_235[5:0];
  assign _EVAL_65 = _EVAL_185 | _EVAL_54;
  assign _EVAL_265 = _EVAL_73 == 4'h0;
  assign _EVAL_42 = ~_EVAL_243;
  assign _EVAL_38 = ~_EVAL_26;
  assign _EVAL_253 = _EVAL_53[4:0];
  assign _EVAL_175 = ~_EVAL_251;
  assign _EVAL_102 = _EVAL_239[0];
  assign _EVAL_55 = _EVAL_70 & _EVAL_103;
  assign _EVAL_284 = _EVAL_10 != 3'h0;
  assign _EVAL_34 = _EVAL_260 == 4'h0;
  assign _EVAL_45 = ~_EVAL_152;
  assign _EVAL_232 = _EVAL_18 ^ 30'h3000;
  assign _EVAL_151 = ~_EVAL_28;
  assign _EVAL_281 = _EVAL_60 | _EVAL_55;
  assign _EVAL_210 = _EVAL_70 & _EVAL_135;
  assign _EVAL_24 = ~_EVAL_255;
  assign _EVAL_79 = _EVAL_266 == 6'h0;
  assign _EVAL_204 = {{22'd0}, _EVAL_196};
  assign _EVAL_40 = _EVAL_263 == 6'h0;
  assign _EVAL_28 = _EVAL_33 | _EVAL_15;
  assign _EVAL_51 = _EVAL_23[31:0];
  assign _EVAL_152 = _EVAL_225 | _EVAL_15;
  assign _EVAL_296 = _EVAL_8 & _EVAL_59;
  assign _EVAL_130 = _EVAL_8 & _EVAL_203;
  assign _EVAL_222 = ~_EVAL_272;
  assign _EVAL_269 = ~_EVAL_72;
  assign _EVAL_290 = _EVAL_50 | _EVAL_15;
  assign _EVAL_187 = _EVAL_266 - 6'h1;
  assign _EVAL_113 = _EVAL_267;
  assign _EVAL_137 = _EVAL_226 | _EVAL_244;
  assign _EVAL_233 = _EVAL & _EVAL_111;
  assign _EVAL_47 = _EVAL_283 == 6'h0;
  assign _EVAL_286 = _EVAL_4 == 3'h5;
  assign _EVAL_277 = _EVAL_187[5:0];
  assign _EVAL_305 = _EVAL_10 <= 3'h4;
  assign _EVAL_181 = _EVAL & _EVAL_251;
  assign _EVAL_236 = 23'hff << _EVAL_2;
  assign _EVAL_250 = _EVAL_34 | _EVAL_15;
  assign _EVAL_29 = ~_EVAL_215;
  assign _EVAL_105 = ~_EVAL_192;
  assign _EVAL_56 = ~_EVAL_58;
  assign _EVAL_81 = _EVAL_122 & _EVAL_179;
  assign _EVAL_242 = _EVAL_16 == 2'h0;
  assign _EVAL_246 = _EVAL_9 == _EVAL_31;
  assign _EVAL_255 = _EVAL_43 | _EVAL_15;
  assign _EVAL_53 = _EVAL_110 ? _EVAL_44 : 8'h0;
  assign _EVAL_121 = _EVAL & _EVAL_86;
  assign _EVAL_107 = _EVAL_96 == 2'h1;
  assign _EVAL_218 = _EVAL_8 & _EVAL_153;
  assign _EVAL_252 = ~_EVAL_15;
  assign _EVAL_306 = ~_EVAL_227;
  assign _EVAL_150 = _EVAL_36 | _EVAL_149;
  assign _EVAL_203 = ~_EVAL_79;
  assign _EVAL_125 = _EVAL_256;
  assign _EVAL_319 = ~_EVAL_104;
  assign _EVAL_189 = {1'b0,$signed(_EVAL_18)};
  assign _EVAL_301 = ~_EVAL_180;
  assign _EVAL_229 = ~_EVAL_145;
  assign _EVAL_172 = _EVAL_271 | _EVAL_15;
  assign _EVAL_312 = _EVAL_162;
  assign _EVAL_110 = _EVAL_120 & _EVAL_175;
  assign _EVAL_231 = ~_EVAL_40;
  assign _EVAL_26 = _EVAL_178 | _EVAL_15;
  assign _EVAL_161 = ~_EVAL_238;
  assign _EVAL_307 = _EVAL_9 == 3'h7;
  assign _EVAL_68 = _EVAL_18[0];
  assign _EVAL_59 = _EVAL_9 == 3'h1;
  assign _EVAL_104 = _EVAL_278 | _EVAL_15;
  assign _EVAL_165 = ~_EVAL_94;
  assign _EVAL_96 = _EVAL_1[2:1];
  assign _EVAL_197 = ~_EVAL_7;
  assign _EVAL_69 = _EVAL_4 == _EVAL_77;
  assign _EVAL_316 = _EVAL_60 | _EVAL_210;
  assign _EVAL_257 = _EVAL_87 | _EVAL_15;
  assign _EVAL_120 = _EVAL_244 & _EVAL_258;
  assign _EVAL_178 = _EVAL_48 | _EVAL_317;
  assign _EVAL_220 = ~_EVAL_311;
  assign _EVAL_238 = _EVAL_242 | _EVAL_15;
  assign _EVAL_254 = _EVAL_196[7:2];
  assign _EVAL_292 = _EVAL_126 | _EVAL_157;
  assign _EVAL_132 = _EVAL & _EVAL_231;
  assign _EVAL_273 = _EVAL_18[1];
  assign _EVAL_198 = {_EVAL_150,_EVAL_221,_EVAL_65,_EVAL_259};
  assign _EVAL_114 = _EVAL_0 == 3'h4;
  assign _EVAL_122 = _EVAL_224 | _EVAL_32;
  assign _EVAL_64 = _EVAL_2[0];
  assign _EVAL_180 = _EVAL_284 | _EVAL_15;
  assign _EVAL_49 = ~_EVAL_198;
  assign _EVAL_140 = ~_EVAL_14;
  assign _EVAL_289 = ~_EVAL_118;
  assign _EVAL_318 = ~_EVAL_129;
  assign _EVAL_52 = _EVAL_308 - 6'h1;
  assign _EVAL_184 = _EVAL_16 <= 2'h2;
  assign _EVAL_30 = ~_EVAL_90;
  assign _EVAL_159 = _EVAL_263 - 6'h1;
  assign _EVAL_193 = _EVAL_8 & _EVAL_194;
  assign _EVAL_90 = _EVAL_9[2];
  assign _EVAL_256 = $signed(_EVAL_189) & -31'sh5000;
  assign _EVAL_21 = _EVAL_188 | _EVAL_15;
  assign _EVAL_315 = _EVAL_316 | _EVAL_15;
  assign _EVAL_200 = _EVAL_138 ? _EVAL_237 : 8'h0;
  assign _EVAL_54 = _EVAL_199 & _EVAL_19;
  assign _EVAL_156 = {1'b0,$signed(_EVAL_261)};
  assign _EVAL_280 = _EVAL_4 <= 3'h6;
  assign _EVAL_196 = ~_EVAL_148;
  assign _EVAL_71 = 23'hff << _EVAL_11;
  assign _EVAL_270 = _EVAL_10 <= 3'h3;
  assign _EVAL_272 = _EVAL_140 | _EVAL_15;
  assign _EVAL_108 = _EVAL_52[5:0];
  assign _EVAL_128 = ~_EVAL_216;
  assign _EVAL_245 = _EVAL_228 | _EVAL_15;
  assign _EVAL_138 = _EVAL_226 & _EVAL_47;
  assign _EVAL_174 = ~_EVAL_106;
  assign _EVAL_276 = _EVAL_67 >> _EVAL_1;
  assign _EVAL_243 = _EVAL_240 | _EVAL_15;
  assign _EVAL_25 = _EVAL_280 | _EVAL_15;
  assign _EVAL_147 = ~_EVAL_245;
  assign _EVAL_258 = _EVAL_308 == 6'h0;
  assign _EVAL_179 = ~_EVAL_253;
  assign _EVAL_288 = $signed(_EVAL_312) == 31'sh0;
  assign _EVAL_160 = _EVAL_60 | _EVAL_84;
  assign _EVAL_111 = _EVAL_4 == 3'h4;
  assign _EVAL_39 = _EVAL_293 == 2'h0;
  assign _EVAL_93 = _EVAL_281 | _EVAL_15;
  assign _EVAL_86 = _EVAL_4 == 3'h2;
  assign _EVAL_23 = _EVAL_177 + 32'h1;
  assign _EVAL_76 = ~_EVAL_257;
  assign _EVAL_82 = _EVAL_212 & _EVAL_41;
  assign _EVAL_91 = _EVAL_276[0];
  assign _EVAL_85 = ~_EVAL_25;
  assign _EVAL_228 = _EVAL_16 == _EVAL_142;
  assign _EVAL_285 = {1'b0,$signed(_EVAL_268)};
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_31 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_63 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_77 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_142 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_168 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_169 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_176 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_177 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_224 = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_241 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_247 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_263 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_264 = _RAND_12[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_266 = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_283 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_295 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_308 = _RAND_16[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_3) begin
    if (_EVAL_143) begin
      _EVAL_31 <= _EVAL_9;
    end
    if (_EVAL_143) begin
      _EVAL_63 <= _EVAL_2;
    end
    if (_EVAL_166) begin
      _EVAL_77 <= _EVAL_4;
    end
    if (_EVAL_166) begin
      _EVAL_142 <= _EVAL_16;
    end
    if (_EVAL_143) begin
      _EVAL_168 <= _EVAL_10;
    end
    if (_EVAL_166) begin
      _EVAL_169 <= _EVAL_11;
    end
    if (_EVAL_166) begin
      _EVAL_176 <= _EVAL_17;
    end
    if (_EVAL_15) begin
      _EVAL_177 <= 32'h0;
    end else if (_EVAL_137) begin
      _EVAL_177 <= 32'h0;
    end else begin
      _EVAL_177 <= _EVAL_51;
    end
    if (_EVAL_15) begin
      _EVAL_224 <= 5'h0;
    end else begin
      _EVAL_224 <= _EVAL_81;
    end
    if (_EVAL_143) begin
      _EVAL_241 <= _EVAL_0;
    end
    if (_EVAL_166) begin
      _EVAL_247 <= _EVAL_1;
    end
    if (_EVAL_15) begin
      _EVAL_263 <= 6'h0;
    end else if (_EVAL_244) begin
      if (_EVAL_40) begin
        if (_EVAL_127) begin
          _EVAL_263 <= _EVAL_136;
        end else begin
          _EVAL_263 <= 6'h0;
        end
      end else begin
        _EVAL_263 <= _EVAL_155;
      end
    end
    if (_EVAL_143) begin
      _EVAL_264 <= _EVAL_18;
    end
    if (_EVAL_15) begin
      _EVAL_266 <= 6'h0;
    end else if (_EVAL_226) begin
      if (_EVAL_79) begin
        if (_EVAL_30) begin
          _EVAL_266 <= _EVAL_254;
        end else begin
          _EVAL_266 <= 6'h0;
        end
      end else begin
        _EVAL_266 <= _EVAL_277;
      end
    end
    if (_EVAL_15) begin
      _EVAL_283 <= 6'h0;
    end else if (_EVAL_226) begin
      if (_EVAL_47) begin
        if (_EVAL_30) begin
          _EVAL_283 <= _EVAL_254;
        end else begin
          _EVAL_283 <= 6'h0;
        end
      end else begin
        _EVAL_283 <= _EVAL_287;
      end
    end
    if (_EVAL_166) begin
      _EVAL_295 <= _EVAL_5;
    end
    if (_EVAL_15) begin
      _EVAL_308 <= 6'h0;
    end else if (_EVAL_244) begin
      if (_EVAL_258) begin
        if (_EVAL_127) begin
          _EVAL_308 <= _EVAL_136;
        end else begin
          _EVAL_308 <= 6'h0;
        end
      end else begin
        _EVAL_308 <= _EVAL_108;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99f1e056)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_274) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b56fcdf5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e496c92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19120be6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_211) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e74370f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(281a97de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b6e717a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cf34932)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_211) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5762fbd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b283c4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e7f3b35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_319) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5faba071)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7585d69e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_274) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e06f8636)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1db8a3fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd96ddda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74e81818)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bfebaea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_319) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40bb65ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac078de1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77bc95fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aaad166d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_314) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(516402ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc63331f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_319) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_314) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32fa1e8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_319) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad723498)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f293344)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2068b47f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9fa468d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_301) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbb80f4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf00df60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f47d7f41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29da8e43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b58a4938)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cf23c74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_319) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97d33184)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36d3153)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45abd8a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee1ca09f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5678390)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a738b9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdbadc3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ac5d37d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebafc39c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_319) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7ccacd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3bfb977)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(210821ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9de13132)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a237bee2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad0ed30a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69e06d2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6cc61c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(196fe8b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_301) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a04c720)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc86bcd8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38147e75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f7e27b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(472a2e1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aeed1061)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e000cea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf1331cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba5a5b45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5be52d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f1ce96d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ceb07bc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_314) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4683d1b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c55e36b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3dc6e7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(141cfd66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84d5392a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dccc683)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d540a86d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6de37857)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12c3ff82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d51fad5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77c988c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98e48f4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94a914c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6535e6f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c902fa47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25a4139c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11a861a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f86704c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2320d025)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f767602)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee6baa6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_314) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e305f30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(269e622a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4a51673)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(983ee83c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
