//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_154(
  input         _EVAL,
  input         _EVAL_0,
  output [1:0]  _EVAL_1,
  output        _EVAL_2,
  input  [1:0]  _EVAL_3,
  output [31:0] _EVAL_4,
  output [31:0] _EVAL_5,
  input  [31:0] _EVAL_6,
  output        _EVAL_7,
  output        _EVAL_8,
  output        _EVAL_9,
  output        _EVAL_10,
  output        _EVAL_11,
  output        _EVAL_12,
  output        _EVAL_13,
  output        _EVAL_14,
  output [7:0]  _EVAL_15,
  input         _EVAL_16,
  input  [31:0] _EVAL_17,
  input  [31:0] _EVAL_18,
  output [31:0] _EVAL_19,
  output        _EVAL_20,
  output        _EVAL_21,
  output        _EVAL_22,
  output        _EVAL_23,
  output        _EVAL_24,
  output [29:0] _EVAL_25,
  output [31:0] _EVAL_26,
  output        _EVAL_27,
  output        _EVAL_28,
  output [31:0] _EVAL_29,
  output [31:0] _EVAL_30,
  output        _EVAL_31,
  output        _EVAL_32,
  output        _EVAL_33,
  output [31:0] _EVAL_34,
  output        _EVAL_35,
  output [1:0]  _EVAL_36,
  output [31:0] _EVAL_37,
  output [1:0]  _EVAL_38,
  input         _EVAL_39,
  input         _EVAL_40,
  output [1:0]  _EVAL_41,
  input         _EVAL_42,
  input         _EVAL_43,
  output        _EVAL_44,
  output        _EVAL_45,
  output [29:0] _EVAL_46,
  output [31:0] _EVAL_47,
  output        _EVAL_48,
  output        _EVAL_49,
  output        _EVAL_50,
  input  [31:0] _EVAL_51,
  output        _EVAL_52,
  output        _EVAL_53,
  output        _EVAL_54,
  input  [7:0]  _EVAL_55,
  output [1:0]  _EVAL_56,
  output        _EVAL_57,
  output        _EVAL_58,
  input         _EVAL_59,
  output        _EVAL_60,
  input         _EVAL_61,
  output [1:0]  _EVAL_62,
  input         _EVAL_63,
  output [31:0] _EVAL_64,
  output [1:0]  _EVAL_65,
  output        _EVAL_66,
  output        _EVAL_67,
  output [29:0] _EVAL_68,
  output        _EVAL_69,
  output        _EVAL_70,
  output        _EVAL_71,
  output        _EVAL_72,
  output [31:0] _EVAL_73,
  output        _EVAL_74,
  output        _EVAL_75,
  input  [11:0] _EVAL_76,
  output        _EVAL_77,
  output        _EVAL_78,
  output [31:0] _EVAL_79,
  output        _EVAL_80,
  output [31:0] _EVAL_81,
  output        _EVAL_82,
  output [31:0] _EVAL_83,
  output        _EVAL_84,
  output [31:0] _EVAL_85,
  output [29:0] _EVAL_86,
  input         _EVAL_87,
  output        _EVAL_88,
  output [1:0]  _EVAL_89,
  output [31:0] _EVAL_90,
  output [31:0] _EVAL_91,
  output        _EVAL_92,
  input         _EVAL_93,
  output        _EVAL_94,
  output [2:0]  _EVAL_95,
  output        _EVAL_96,
  output        _EVAL_97,
  input  [2:0]  _EVAL_98,
  output        _EVAL_99,
  output        _EVAL_100,
  input  [11:0] _EVAL_101,
  output        _EVAL_102,
  output        _EVAL_103,
  output [1:0]  _EVAL_104,
  output        _EVAL_105,
  output        _EVAL_106,
  input  [31:0] _EVAL_107,
  input  [7:0]  _EVAL_108,
  input  [31:0] _EVAL_109,
  output        _EVAL_110,
  output        _EVAL_111,
  output        _EVAL_112,
  input         _EVAL_113,
  output        _EVAL_114,
  output        _EVAL_115,
  output [1:0]  _EVAL_116,
  output        _EVAL_117,
  output        _EVAL_118,
  output        _EVAL_119,
  output        _EVAL_120,
  input         _EVAL_121,
  output        _EVAL_122,
  output        _EVAL_123,
  output        _EVAL_124,
  output [26:0] _EVAL_125,
  output        _EVAL_126,
  output [1:0]  _EVAL_127,
  output [1:0]  _EVAL_128,
  output [1:0]  _EVAL_129,
  output [1:0]  _EVAL_130,
  output        _EVAL_131,
  output        _EVAL_132,
  output [31:0] _EVAL_133,
  output        _EVAL_134,
  output [1:0]  _EVAL_135,
  output        _EVAL_136,
  output [1:0]  _EVAL_137,
  output        _EVAL_138,
  output        _EVAL_139,
  output        _EVAL_140,
  output [1:0]  _EVAL_141
);
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire [1:0] _EVAL_151;
  wire [33:0] _EVAL_152;
  reg  _EVAL_153;
  reg [31:0] _RAND_0;
  wire [7:0] _EVAL_155;
  reg [31:0] _EVAL_156;
  reg [31:0] _RAND_1;
  wire  _EVAL_157;
  wire [7:0] _EVAL_158;
  wire  _EVAL_159;
  wire [30:0] _EVAL_160;
  wire  _EVAL_162;
  reg  _EVAL_163;
  reg [31:0] _RAND_2;
  wire  _EVAL_164;
  wire  _EVAL_167;
  wire [29:0] _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire [5:0] _EVAL_172;
  wire  _EVAL_173;
  wire [31:0] _EVAL_176;
  wire  _EVAL_177;
  reg [31:0] _EVAL_178;
  reg [31:0] _RAND_3;
  wire  _EVAL_179;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_187;
  wire  _EVAL_189;
  wire [1:0] _EVAL_190;
  reg  _EVAL_192;
  reg [31:0] _RAND_4;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire [7:0] _EVAL_198;
  wire [7:0] _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire [31:0] _EVAL_204;
  wire [142:0] _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire [3:0] _EVAL_214;
  wire [39:0] _EVAL_215;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire [142:0] _EVAL_223;
  wire [7:0] _EVAL_224;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_230;
  wire  _EVAL_232;
  wire  _EVAL_234;
  wire [142:0] _EVAL_235;
  wire  _EVAL_236;
  wire [5:0] _EVAL_237;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire [1:0] _EVAL_243;
  wire [7:0] _EVAL_244;
  wire [6:0] _EVAL_245;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire [6:0] _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_256;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  reg  _EVAL_261;
  reg [31:0] _RAND_5;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire [1:0] _EVAL_266;
  wire  _EVAL_267;
  reg  _EVAL_269;
  reg [31:0] _RAND_6;
  wire  _EVAL_270;
  reg  _EVAL_272;
  reg [31:0] _RAND_7;
  wire  _EVAL_273;
  wire [7:0] _EVAL_274;
  wire [31:0] _EVAL_275;
  wire  _EVAL_277;
  wire [7:0] _EVAL_278;
  reg [31:0] _EVAL_279;
  reg [31:0] _RAND_8;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire [57:0] _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire [31:0] _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire [1:0] _EVAL_296;
  wire  _EVAL_297;
  wire [5:0] _EVAL_298;
  wire [25:0] _EVAL_299;
  wire [7:0] _EVAL_301;
  wire  _EVAL_302;
  wire [30:0] _EVAL_303;
  wire [31:0] _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_308;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  reg  _EVAL_315;
  reg [31:0] _RAND_9;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire [7:0] _EVAL_319;
  wire  _EVAL_320;
  wire  _EVAL_322;
  wire [142:0] _EVAL_325;
  wire  _EVAL_326;
  wire  _EVAL_327;
  wire  _EVAL_328;
  wire  _EVAL_329;
  wire [7:0] _EVAL_330;
  reg  _EVAL_331;
  reg [31:0] _RAND_10;
  wire  _EVAL_332;
  reg [29:0] _EVAL_333;
  reg [31:0] _RAND_11;
  reg  _EVAL_334;
  reg [31:0] _RAND_12;
  wire  _EVAL_335;
  wire  _EVAL_336;
  wire  _EVAL_337;
  wire [7:0] _EVAL_339;
  wire  _EVAL_340;
  wire  _EVAL_341;
  wire  _EVAL_344;
  wire  _EVAL_345;
  wire  _EVAL_350;
  wire  _EVAL_351;
  wire  _EVAL_353;
  wire [142:0] _EVAL_354;
  wire [7:0] _EVAL_356;
  wire  _EVAL_357;
  wire  _EVAL_361;
  wire  _EVAL_362;
  wire  _EVAL_363;
  wire [5:0] _EVAL_364;
  wire  _EVAL_365;
  wire [39:0] _EVAL_366;
  wire  _EVAL_367;
  wire  _EVAL_368;
  wire [31:0] _EVAL_369;
  wire  _EVAL_370;
  wire  _EVAL_373;
  wire  _EVAL_374;
  wire  _EVAL_375;
  wire  _EVAL_379;
  wire  _EVAL_380;
  wire  _EVAL_381;
  wire [7:0] _EVAL_382;
  wire  _EVAL_385;
  wire  _EVAL_386;
  wire [31:0] _EVAL_387;
  wire [31:0] _EVAL_388;
  wire  _EVAL_390;
  wire  _EVAL_391;
  wire  _EVAL_394;
  wire [6:0] _EVAL_397;
  wire  _EVAL_399;
  wire  _EVAL_402;
  wire  _EVAL_404;
  wire  _EVAL_405;
  reg  _EVAL_406;
  reg [31:0] _RAND_13;
  wire  _EVAL_407;
  wire  _EVAL_408;
  wire [7:0] _EVAL_409;
  wire  _EVAL_411;
  wire [31:0] _EVAL_412;
  wire  _EVAL_413;
  wire  _EVAL_414;
  wire  _EVAL_415;
  wire [1:0] _EVAL_417;
  wire [7:0] _EVAL_419;
  wire [7:0] _EVAL_420;
  wire  _EVAL_421;
  wire  _EVAL_422;
  wire  _EVAL_423;
  wire [63:0] _EVAL_424;
  wire  _EVAL_425;
  wire  _EVAL_427;
  wire  _EVAL_428;
  reg [5:0] _EVAL_429;
  reg [31:0] _RAND_14;
  wire  _EVAL_430;
  wire  _EVAL_431;
  wire [31:0] _EVAL_432;
  wire  _EVAL_435;
  wire  _EVAL_436;
  wire  _EVAL_437;
  reg [1:0] _EVAL_438;
  reg [31:0] _RAND_15;
  wire  _EVAL_439;
  reg [1:0] _EVAL_440;
  reg [31:0] _RAND_16;
  wire  _EVAL_441;
  wire [31:0] _EVAL_442;
  wire [5:0] _EVAL_444;
  wire  _EVAL_445;
  wire  _EVAL_446;
  wire  _EVAL_447;
  wire [3:0] _EVAL_448;
  wire  _EVAL_449;
  wire  _EVAL_452;
  wire [5:0] _EVAL_453;
  wire [7:0] _EVAL_454;
  wire  _EVAL_456;
  wire  _EVAL_457;
  reg [31:0] _EVAL_459;
  reg [31:0] _RAND_17;
  wire  _EVAL_460;
  wire  _EVAL_461;
  wire  _EVAL_463;
  wire [7:0] _EVAL_466;
  wire  _EVAL_467;
  wire  _EVAL_468;
  wire  _EVAL_469;
  wire  _EVAL_470;
  wire  _EVAL_471;
  wire [7:0] _EVAL_472;
  wire  _EVAL_473;
  wire  _EVAL_474;
  wire  _EVAL_475;
  wire  _EVAL_477;
  wire [6:0] _EVAL_478;
  wire [30:0] _EVAL_480;
  wire  _EVAL_481;
  wire [7:0] _EVAL_482;
  wire  _EVAL_483;
  reg  _EVAL_484;
  reg [31:0] _RAND_18;
  wire  _EVAL_486;
  wire  _EVAL_487;
  wire  _EVAL_489;
  wire  _EVAL_490;
  wire [6:0] _EVAL_491;
  wire [6:0] _EVAL_492;
  wire  _EVAL_493;
  reg  _EVAL_494;
  reg [31:0] _RAND_19;
  reg  _EVAL_495;
  reg [31:0] _RAND_20;
  wire [31:0] _EVAL_497;
  wire [7:0] _EVAL_498;
  wire  _EVAL_499;
  wire  _EVAL_500;
  wire  _EVAL_501;
  wire  _EVAL_502;
  wire [29:0] _EVAL_504;
  wire  _EVAL_505;
  wire  _EVAL_506;
  reg  _EVAL_507;
  reg [31:0] _RAND_21;
  wire [142:0] _EVAL_508;
  wire  _EVAL_509;
  wire  _EVAL_512;
  wire  _EVAL_513;
  wire  _EVAL_514;
  wire  _EVAL_515;
  wire [31:0] _EVAL_519;
  wire  _EVAL_520;
  wire  _EVAL_521;
  wire [30:0] _EVAL_522;
  wire  _EVAL_523;
  wire  _EVAL_524;
  reg  _EVAL_525;
  reg [31:0] _RAND_22;
  wire  _EVAL_526;
  wire [30:0] _EVAL_531;
  wire  _EVAL_532;
  wire  _EVAL_534;
  wire  _EVAL_535;
  wire  _EVAL_537;
  wire  _EVAL_539;
  wire  _EVAL_540;
  wire [7:0] _EVAL_542;
  wire  _EVAL_543;
  wire  _EVAL_544;
  wire  _EVAL_546;
  wire  _EVAL_547;
  wire  _EVAL_550;
  wire  _EVAL_551;
  wire  _EVAL_552;
  wire [33:0] _EVAL_553;
  wire  _EVAL_554;
  wire  _EVAL_555;
  wire  _EVAL_556;
  wire  _EVAL_557;
  wire  _EVAL_558;
  wire  _EVAL_559;
  wire [31:0] _EVAL_560;
  wire  _EVAL_562;
  wire [7:0] _EVAL_563;
  wire [6:0] _EVAL_564;
  wire [7:0] _EVAL_565;
  wire [6:0] _EVAL_567;
  wire  _EVAL_568;
  wire [6:0] _EVAL_570;
  wire [32:0] _EVAL_571;
  wire [142:0] _EVAL_572;
  wire  _EVAL_573;
  wire [39:0] _EVAL_576;
  wire [31:0] _EVAL_578;
  wire [63:0] _EVAL_581;
  wire  _EVAL_582;
  wire  _EVAL_583;
  wire  _EVAL_584;
  wire [7:0] _EVAL_586;
  wire  _EVAL_588;
  wire [30:0] _EVAL_589;
  wire [7:0] _EVAL_590;
  wire  _EVAL_591;
  wire  _EVAL_594;
  wire  _EVAL_596;
  wire [7:0] _EVAL_597;
  wire  _EVAL_598;
  wire [142:0] _EVAL_599;
  wire  _EVAL_601;
  wire [7:0] _EVAL_605;
  wire  _EVAL_606;
  wire [7:0] _EVAL_607;
  reg  _EVAL_608;
  reg [31:0] _RAND_23;
  wire  _EVAL_609;
  wire  _EVAL_610;
  wire [31:0] _EVAL_611;
  reg  _EVAL_612;
  reg [31:0] _RAND_24;
  wire  _EVAL_613;
  wire [31:0] _EVAL_616;
  wire  _EVAL_617;
  wire  _EVAL_618;
  reg [11:0] _EVAL_619;
  reg [31:0] _RAND_25;
  wire [31:0] _EVAL_620;
  wire  _EVAL_621;
  wire [7:0] _EVAL_624;
  wire  _EVAL_625;
  wire  _EVAL_626;
  wire [31:0] _EVAL_627;
  wire [142:0] _EVAL_628;
  wire [6:0] _EVAL_629;
  wire  _EVAL_631;
  wire  _EVAL_632;
  wire [142:0] _EVAL_634;
  wire  _EVAL_639;
  wire  _EVAL_640;
  wire  _EVAL_641;
  wire  _EVAL_642;
  wire [30:0] _EVAL_644;
  wire [6:0] _EVAL_645;
  wire  _EVAL_646;
  wire  _EVAL_648;
  wire [7:0] _EVAL_649;
  wire  _EVAL_650;
  wire  _EVAL_653;
  wire  _EVAL_655;
  wire [7:0] _EVAL_657;
  wire  _EVAL_659;
  wire  _EVAL_660;
  wire  _EVAL_661;
  wire  _EVAL_662;
  wire [31:0] _EVAL_663;
  wire  _EVAL_666;
  wire [4:0] _EVAL_667;
  wire [142:0] _EVAL_668;
  wire  _EVAL_669;
  wire [7:0] _EVAL_670;
  wire  _EVAL_671;
  wire  _EVAL_672;
  reg  _EVAL_673;
  reg [31:0] _RAND_26;
  wire [7:0] _EVAL_674;
  wire  _EVAL_675;
  wire  _EVAL_677;
  wire  _EVAL_681;
  wire [7:0] _EVAL_683;
  wire [7:0] _EVAL_684;
  reg  _EVAL_685;
  reg [31:0] _RAND_27;
  wire  _EVAL_686;
  wire  _EVAL_688;
  wire  _EVAL_690;
  wire  _EVAL_691;
  wire  _EVAL_692;
  wire  _EVAL_693;
  wire [25:0] _EVAL_694;
  wire [31:0] _EVAL_698;
  reg  _EVAL_699;
  reg [31:0] _RAND_28;
  wire  _EVAL_700;
  wire  _EVAL_701;
  wire  _EVAL_702;
  wire [25:0] _EVAL_703;
  wire  _EVAL_704;
  wire  _EVAL_705;
  wire [7:0] _EVAL_706;
  wire  _EVAL_707;
  wire [30:0] _EVAL_708;
  wire  _EVAL_710;
  wire  _EVAL_711;
  wire [6:0] _EVAL_712;
  wire [7:0] _EVAL_713;
  wire  _EVAL_714;
  wire [31:0] _EVAL_715;
  wire  _EVAL_716;
  wire  _EVAL_717;
  wire  _EVAL_718;
  wire  _EVAL_719;
  wire  _EVAL_721;
  wire  _EVAL_722;
  wire  _EVAL_724;
  wire [31:0] _EVAL_726;
  wire  _EVAL_727;
  reg [2:0] _EVAL_728;
  reg [31:0] _RAND_29;
  reg  _EVAL_729;
  reg [31:0] _RAND_30;
  wire  _EVAL_730;
  wire [1:0] _EVAL_731;
  wire [7:0] _EVAL_732;
  wire  _EVAL_733;
  wire [31:0] _EVAL_734;
  wire  _EVAL_736;
  wire [7:0] _EVAL_737;
  wire [31:0] _EVAL_739;
  wire  _EVAL_740;
  wire [7:0] _EVAL_741;
  wire  _EVAL_742;
  wire  _EVAL_743;
  wire  _EVAL_745;
  reg [57:0] _EVAL_746;
  reg [63:0] _RAND_31;
  wire [7:0] _EVAL_748;
  wire  _EVAL_749;
  wire [142:0] _EVAL_751;
  reg  _EVAL_753;
  reg [31:0] _RAND_32;
  wire [4:0] _EVAL_754;
  wire  _EVAL_758;
  wire  _EVAL_759;
  wire [31:0] _EVAL_761;
  reg  _EVAL_762;
  reg [31:0] _RAND_33;
  wire  _EVAL_763;
  wire  _EVAL_765;
  reg [31:0] _EVAL_767;
  reg [31:0] _RAND_34;
  wire [4:0] _EVAL_768;
  wire  _EVAL_769;
  wire [31:0] _EVAL_770;
  wire  _EVAL_771;
  wire [102:0] _EVAL_772;
  wire [6:0] _EVAL_773;
  reg [1:0] _EVAL_774;
  reg [31:0] _RAND_35;
  wire [7:0] _EVAL_775;
  wire [142:0] _EVAL_776;
  wire  _EVAL_777;
  wire [6:0] _EVAL_778;
  wire  _EVAL_779;
  wire [31:0] _EVAL_780;
  wire  _EVAL_781;
  wire [5:0] _EVAL_782;
  wire  _EVAL_785;
  wire [4:0] _EVAL_786;
  wire  _EVAL_787;
  wire  _EVAL_788;
  wire  _EVAL_789;
  wire  _EVAL_790;
  wire  _EVAL_791;
  wire  _EVAL_795;
  wire  _EVAL_798;
  wire  _EVAL_799;
  wire  _EVAL_800;
  wire [6:0] _EVAL_801;
  wire  _EVAL_802;
  wire  _EVAL_804;
  wire  _EVAL_805;
  wire  _EVAL_806;
  wire  _EVAL_808;
  wire  _EVAL_809;
  wire  _EVAL_810;
  wire  _EVAL_811;
  wire  _EVAL_813;
  wire [4:0] _EVAL_814;
  wire  _EVAL_815;
  wire  _EVAL_817;
  wire  _EVAL_818;
  reg  _EVAL_819;
  reg [31:0] _RAND_36;
  reg [1:0] _EVAL_820;
  reg [31:0] _RAND_37;
  wire  _EVAL_821;
  wire  _EVAL_822;
  wire  _EVAL_824;
  wire  _EVAL_825;
  wire  _EVAL_826;
  wire  _EVAL_828;
  wire  _EVAL_829;
  wire  _EVAL_830;
  wire  _EVAL_832;
  wire [11:0] _EVAL_834;
  wire  _EVAL_835;
  wire  _EVAL_836;
  wire [7:0] _EVAL_840;
  wire  _EVAL_841;
  wire  _EVAL_843;
  reg  _EVAL_845;
  reg [31:0] _RAND_38;
  wire [6:0] _EVAL_849;
  reg [29:0] _EVAL_850;
  reg [31:0] _RAND_39;
  wire  _EVAL_851;
  wire [142:0] _EVAL_852;
  wire [7:0] _EVAL_853;
  wire [142:0] _EVAL_854;
  wire  _EVAL_855;
  wire  _EVAL_856;
  wire [7:0] _EVAL_857;
  wire [7:0] _EVAL_859;
  wire [4:0] _EVAL_860;
  wire  _EVAL_861;
  wire [1:0] _EVAL_862;
  reg [7:0] _EVAL_864;
  reg [31:0] _RAND_40;
  wire [24:0] _EVAL_865;
  wire  _EVAL_866;
  wire  _EVAL_870;
  wire  _EVAL_871;
  wire  _EVAL_872;
  wire  _EVAL_873;
  wire  _EVAL_874;
  wire [1:0] _EVAL_875;
  wire  _EVAL_876;
  wire  _EVAL_877;
  wire [1:0] _EVAL_879;
  reg [31:0] _EVAL_880;
  reg [31:0] _RAND_41;
  wire [31:0] _EVAL_882;
  wire  _EVAL_883;
  wire  _EVAL_884;
  wire  _EVAL_885;
  wire [31:0] _EVAL_886;
  wire [7:0] _EVAL_887;
  wire  _EVAL_889;
  wire  _EVAL_890;
  reg  _EVAL_891;
  reg [31:0] _RAND_42;
  wire  _EVAL_892;
  wire  _EVAL_895;
  wire [142:0] _EVAL_896;
  wire [7:0] _EVAL_897;
  wire [142:0] _EVAL_899;
  wire  _EVAL_901;
  wire  _EVAL_902;
  wire  _EVAL_903;
  wire [7:0] _EVAL_904;
  wire  _EVAL_905;
  wire  _EVAL_906;
  wire [7:0] _EVAL_907;
  reg [1:0] _EVAL_908;
  reg [31:0] _RAND_43;
  wire  _EVAL_909;
  wire  _EVAL_910;
  wire [7:0] _EVAL_911;
  wire [6:0] _EVAL_912;
  wire [5:0] _EVAL_913;
  wire [2:0] _EVAL_914;
  wire [33:0] _EVAL_916;
  wire  _EVAL_917;
  wire  _EVAL_918;
  wire [6:0] _EVAL_919;
  reg  _EVAL_920;
  reg [31:0] _RAND_44;
  wire [31:0] _EVAL_922;
  wire  _EVAL_923;
  reg [26:0] _EVAL_924;
  reg [31:0] _RAND_45;
  wire  _EVAL_925;
  wire  _EVAL_926;
  wire  _EVAL_927;
  wire  _EVAL_928;
  wire  _EVAL_932;
  wire  _EVAL_933;
  wire  _EVAL_934;
  reg  _EVAL_935;
  reg [31:0] _RAND_46;
  wire [31:0] _EVAL_936;
  wire  _EVAL_937;
  wire [6:0] _EVAL_938;
  wire [31:0] _EVAL_941;
  wire  _EVAL_943;
  wire [31:0] _EVAL_944;
  wire  _EVAL_946;
  wire  _EVAL_947;
  wire [142:0] _EVAL_948;
  wire [6:0] _EVAL_950;
  wire  _EVAL_952;
  wire  _EVAL_953;
  wire  _EVAL_954;
  wire [7:0] _EVAL_956;
  wire [3:0] _EVAL_957;
  wire  _EVAL_959;
  wire  _EVAL_960;
  wire [6:0] _EVAL_961;
  wire  _EVAL_962;
  wire  _EVAL_964;
  wire  _EVAL_966;
  wire  _EVAL_967;
  wire  _EVAL_968;
  wire [142:0] _EVAL_969;
  wire  _EVAL_970;
  wire  _EVAL_971;
  wire  _EVAL_972;
  wire  _EVAL_973;
  wire [3:0] _EVAL_974;
  reg  _EVAL_975;
  reg [31:0] _RAND_47;
  wire  _EVAL_976;
  wire  _EVAL_977;
  wire  _EVAL_978;
  wire [7:0] _EVAL_979;
  wire [31:0] _EVAL_980;
  wire [7:0] _EVAL_981;
  wire  _EVAL_982;
  wire  _EVAL_985;
  wire  _EVAL_986;
  wire  _EVAL_993;
  wire  _EVAL_995;
  wire  _EVAL_996;
  wire  _EVAL_1000;
  wire  _EVAL_1001;
  wire  _EVAL_1004;
  wire  _EVAL_1006;
  wire [6:0] _EVAL_1007;
  wire  _EVAL_1009;
  wire  _EVAL_1010;
  wire [142:0] _EVAL_1011;
  wire  _EVAL_1012;
  wire [7:0] _EVAL_1013;
  wire  _EVAL_1015;
  wire  _EVAL_1016;
  wire  _EVAL_1017;
  wire [6:0] _EVAL_1018;
  reg  _EVAL_1019;
  reg [31:0] _RAND_48;
  wire [5:0] _EVAL_1020;
  wire [6:0] _EVAL_1021;
  wire  _EVAL_1024;
  wire  _EVAL_1026;
  wire  _EVAL_1027;
  wire  _EVAL_1029;
  wire  _EVAL_1030;
  wire  _EVAL_1031;
  wire [31:0] _EVAL_1032;
  wire [7:0] _EVAL_1033;
  wire [7:0] _EVAL_1035;
  wire  _EVAL_1036;
  wire  _EVAL_1037;
  wire  _EVAL_1039;
  wire [3:0] _EVAL_1040;
  wire  _EVAL_1044;
  wire [31:0] _EVAL_1045;
  reg [31:0] _EVAL_1047;
  reg [31:0] _RAND_49;
  wire  _EVAL_1050;
  wire [1:0] _EVAL_1051;
  wire [1:0] _EVAL_1054;
  wire  _EVAL_1056;
  wire [7:0] _EVAL_1058;
  wire [142:0] _EVAL_1060;
  wire [7:0] _EVAL_1061;
  wire  _EVAL_1062;
  wire  _EVAL_1063;
  wire  _EVAL_1064;
  wire [6:0] _EVAL_1065;
  wire  _EVAL_1069;
  wire [142:0] _EVAL_1070;
  wire  _EVAL_1071;
  wire [142:0] _EVAL_1073;
  wire [6:0] _EVAL_1074;
  wire [142:0] _EVAL_1077;
  wire [142:0] _EVAL_1078;
  wire [30:0] _EVAL_1079;
  reg  _EVAL_1080;
  reg [31:0] _RAND_50;
  wire  _EVAL_1081;
  wire  _EVAL_1083;
  wire [7:0] _EVAL_1085;
  wire [7:0] _EVAL_1087;
  wire [7:0] _EVAL_1088;
  wire  _EVAL_1089;
  wire  _EVAL_1090;
  wire [7:0] _EVAL_1093;
  wire [4:0] _EVAL_1094;
  wire  _EVAL_1095;
  wire [63:0] _EVAL_1097;
  wire  _EVAL_1098;
  wire  _EVAL_1099;
  wire  _EVAL_1104;
  wire  _EVAL_1105;
  wire  _EVAL_1106;
  wire  _EVAL_1107;
  wire  _EVAL_1108;
  wire  _EVAL_1110;
  wire [7:0] _EVAL_1112;
  wire  _EVAL_1113;
  wire  _EVAL_1114;
  wire [7:0] _EVAL_1115;
  wire [142:0] _EVAL_1116;
  wire  _EVAL_1117;
  wire  _EVAL_1118;
  wire  _EVAL_1119;
  wire  _EVAL_1121;
  wire  _EVAL_1122;
  wire  _EVAL_1123;
  wire [31:0] _EVAL_1124;
  wire  _EVAL_1125;
  wire [7:0] _EVAL_1126;
  wire  _EVAL_1127;
  wire  _EVAL_1128;
  wire  _EVAL_1129;
  wire  _EVAL_1130;
  wire [31:0] _EVAL_1131;
  wire [7:0] _EVAL_1132;
  wire  _EVAL_1133;
  wire  _EVAL_1134;
  wire [31:0] _EVAL_1136;
  wire  _EVAL_1137;
  wire  _EVAL_1141;
  reg [1:0] _EVAL_1142;
  reg [31:0] _RAND_51;
  wire [15:0] _EVAL_1144;
  wire  _EVAL_1146;
  wire  _EVAL_1148;
  wire  _EVAL_1149;
  wire  _EVAL_1150;
  wire [7:0] _EVAL_1152;
  wire  _EVAL_1154;
  wire  _EVAL_1157;
  wire  _EVAL_1158;
  wire  _EVAL_1159;
  wire [7:0] _EVAL_1163;
  wire [7:0] _EVAL_1164;
  wire  _EVAL_1165;
  wire  _EVAL_1169;
  wire  _EVAL_1171;
  reg  _EVAL_1172;
  reg [31:0] _RAND_52;
  wire  _EVAL_1173;
  wire  _EVAL_1174;
  wire  _EVAL_1175;
  wire  _EVAL_1176;
  wire  _EVAL_1177;
  wire  _EVAL_1179;
  wire [6:0] _EVAL_1181;
  wire  _EVAL_1184;
  wire  _EVAL_1185;
  wire [63:0] _EVAL_1187;
  wire  _EVAL_1189;
  wire [5:0] _EVAL_1190;
  wire  _EVAL_1191;
  wire [142:0] _EVAL_1192;
  wire  _EVAL_1193;
  wire  _EVAL_1194;
  wire  _EVAL_1195;
  wire [4:0] _EVAL_1197;
  wire  _EVAL_1199;
  wire  _EVAL_1200;
  wire  _EVAL_1201;
  wire  _EVAL_1202;
  wire  _EVAL_1203;
  wire [7:0] _EVAL_1204;
  wire  _EVAL_1205;
  wire  _EVAL_1207;
  wire  _EVAL_1208;
  wire  _EVAL_1209;
  wire  _EVAL_1212;
  wire  _EVAL_1213;
  wire  _EVAL_1214;
  wire  _EVAL_1215;
  wire  _EVAL_1217;
  wire [5:0] _EVAL_1218;
  wire  _EVAL_1223;
  wire  _EVAL_1224;
  wire [7:0] _EVAL_1225;
  wire  _EVAL_1226;
  wire  _EVAL_1228;
  wire [32:0] _EVAL_1229;
  wire  _EVAL_1231;
  wire  _EVAL_1233;
  wire  _EVAL_1235;
  wire  _EVAL_1236;
  wire [31:0] _EVAL_1238;
  reg [31:0] _EVAL_1239;
  reg [31:0] _RAND_53;
  wire [7:0] _EVAL_1240;
  wire  _EVAL_1241;
  wire [9:0] _EVAL_1243;
  wire [63:0] _EVAL_1244;
  wire  _EVAL_1245;
  reg [1:0] _EVAL_1246;
  reg [31:0] _RAND_54;
  wire  _EVAL_1247;
  wire [1:0] _EVAL_1248;
  wire  _EVAL_1252;
  wire [63:0] _EVAL_1255;
  wire  _EVAL_1258;
  wire  _EVAL_1259;
  wire [4:0] _EVAL_1261;
  wire  _EVAL_1264;
  wire [30:0] _EVAL_1265;
  reg [7:0] _EVAL_1267;
  reg [31:0] _RAND_55;
  reg  _EVAL_1268;
  reg [31:0] _RAND_56;
  wire  _EVAL_1269;
  wire  _EVAL_1270;
  reg [31:0] _EVAL_1271;
  reg [31:0] _RAND_57;
  wire  _EVAL_1272;
  wire  _EVAL_1273;
  wire  _EVAL_1274;
  wire  _EVAL_1275;
  wire [7:0] _EVAL_1276;
  wire [31:0] _EVAL_1277;
  wire  _EVAL_1278;
  reg [29:0] _EVAL_1279;
  reg [31:0] _RAND_58;
  wire  _EVAL_1280;
  wire  _EVAL_1281;
  wire  _EVAL_1282;
  wire [7:0] _EVAL_1283;
  wire  _EVAL_1286;
  wire  _EVAL_1287;
  wire  _EVAL_1289;
  wire [142:0] _EVAL_1290;
  wire  _EVAL_1291;
  wire  _EVAL_1292;
  wire [7:0] _EVAL_1293;
  wire  _EVAL_1294;
  wire  _EVAL_1295;
  wire  _EVAL_1297;
  wire  _EVAL_1298;
  wire [6:0] _EVAL_1299;
  wire  _EVAL_1300;
  wire  _EVAL_1302;
  wire  _EVAL_1303;
  wire  _EVAL_1305;
  wire  _EVAL_1306;
  wire  _EVAL_1308;
  wire  _EVAL_1310;
  wire [7:0] _EVAL_1312;
  wire [7:0] _EVAL_1313;
  wire  _EVAL_1315;
  reg  _EVAL_1318;
  reg [31:0] _RAND_59;
  wire  _EVAL_1319;
  wire  _EVAL_1321;
  wire  _EVAL_1322;
  wire  _EVAL_1323;
  wire  _EVAL_1324;
  wire  _EVAL_1325;
  wire [142:0] _EVAL_1326;
  wire [7:0] _EVAL_1327;
  wire  _EVAL_1329;
  wire  _EVAL_1330;
  wire  _EVAL_1331;
  wire [32:0] _EVAL_1332;
  wire [6:0] _EVAL_1333;
  wire  _EVAL_1334;
  wire  _EVAL_1335;
  wire [7:0] _EVAL_1337;
  wire [6:0] _EVAL_1338;
  wire [7:0] _EVAL_1343;
  wire  _EVAL_1344;
  wire  _EVAL_1347;
  wire  _EVAL_1348;
  wire [31:0] _EVAL_1349;
  wire  _EVAL_1350;
  reg [31:0] _EVAL_1351;
  reg [31:0] _RAND_60;
  reg  _EVAL_1353;
  reg [31:0] _RAND_61;
  wire  _EVAL_1356;
  wire [7:0] _EVAL_1359;
  wire [7:0] _EVAL_1360;
  wire  _EVAL_1362;
  wire  _EVAL_1364;
  wire  _EVAL_1365;
  wire  _EVAL_1366;
  wire  _EVAL_1367;
  wire  _EVAL_1371;
  wire [30:0] _EVAL_1372;
  wire  _EVAL_1375;
  wire  _EVAL_1376;
  wire  _EVAL_1377;
  wire [7:0] _EVAL_1379;
  wire  _EVAL_1380;
  wire [6:0] _EVAL_1381;
  wire  _EVAL_1382;
  wire  _EVAL_1383;
  wire  _EVAL_1384;
  wire  _EVAL_1385;
  wire  _EVAL_1386;
  wire  _EVAL_1387;
  wire  _EVAL_1388;
  wire  _EVAL_1389;
  wire  _EVAL_1390;
  wire  _EVAL_1391;
  wire  _EVAL_1392;
  wire  _EVAL_1393;
  wire  _EVAL_1394;
  wire [31:0] _EVAL_1395;
  wire  _EVAL_1396;
  wire  _EVAL_1397;
  wire  _EVAL_1398;
  wire [15:0] _EVAL_1399;
  wire  _EVAL_1400;
  wire [7:0] _EVAL_1401;
  wire [5:0] _EVAL_1403;
  wire  _EVAL_1404;
  wire [6:0] _EVAL_1405;
  wire  _EVAL_1407;
  wire  _EVAL_1408;
  wire  _EVAL_1410;
  wire  _EVAL_1411;
  wire  _EVAL_1412;
  wire [7:0] _EVAL_1413;
  wire  _EVAL_1414;
  wire  _EVAL_1415;
  wire  _EVAL_1416;
  wire  _EVAL_1418;
  wire  _EVAL_1419;
  wire [142:0] _EVAL_1420;
  wire [31:0] _EVAL_1421;
  wire [31:0] _EVAL_1422;
  wire  _EVAL_1423;
  wire  _EVAL_1424;
  wire  _EVAL_1427;
  wire [6:0] _EVAL_1428;
  wire  _EVAL_1429;
  wire [5:0] _EVAL_1433;
  wire [31:0] _EVAL_1435;
  wire [31:0] _EVAL_1436;
  wire  _EVAL_1439;
  wire  _EVAL_1440;
  wire  _EVAL_1446;
  reg [31:0] _EVAL_1447;
  reg [31:0] _RAND_62;
  wire  _EVAL_1448;
  reg  _EVAL_1450;
  reg [31:0] _RAND_63;
  reg [1:0] _EVAL_1451;
  reg [31:0] _RAND_64;
  wire  _EVAL_1452;
  wire  _EVAL_1453;
  wire [31:0] _EVAL_1454;
  wire  _EVAL_1455;
  wire  _EVAL_1457;
  wire  _EVAL_1458;
  wire  _EVAL_1459;
  wire [3:0] _EVAL_1460;
  wire  _EVAL_1462;
  wire  _EVAL_1463;
  wire  _EVAL_1464;
  wire [23:0] _EVAL_1465;
  reg  _EVAL_1466;
  reg [31:0] _RAND_65;
  reg  _EVAL_1467;
  reg [31:0] _RAND_66;
  wire  _EVAL_1469;
  wire [63:0] _EVAL_1472;
  wire [7:0] _EVAL_1473;
  wire  _EVAL_1474;
  wire  _EVAL_1475;
  wire  _EVAL_1476;
  wire  _EVAL_1478;
  wire  _EVAL_1479;
  wire [6:0] _EVAL_1480;
  wire [4:0] _EVAL_1482;
  wire [6:0] _EVAL_1484;
  wire [6:0] _EVAL_1485;
  wire [4:0] _EVAL_1486;
  wire [3:0] _EVAL_1487;
  wire  _EVAL_1488;
  wire  _EVAL_1489;
  reg  _EVAL_1491;
  reg [31:0] _RAND_67;
  wire  _EVAL_1492;
  reg  _EVAL_1493;
  reg [31:0] _RAND_68;
  wire [31:0] _EVAL_1494;
  wire [31:0] _EVAL_1495;
  wire  _EVAL_1499;
  wire [142:0] _EVAL_1500;
  wire [7:0] _EVAL_1501;
  wire  _EVAL_1502;
  wire  _EVAL_1505;
  wire [29:0] _EVAL_1506;
  reg  _EVAL_1507;
  reg [31:0] _RAND_69;
  wire  _EVAL_1508;
  wire [7:0] _EVAL_1510;
  reg [1:0] _EVAL_1512;
  reg [31:0] _RAND_70;
  wire  _EVAL_1513;
  wire  _EVAL_1514;
  wire [63:0] _EVAL_1515;
  wire  _EVAL_1517;
  wire  _EVAL_1518;
  wire  _EVAL_1519;
  wire [142:0] _EVAL_1520;
  wire  _EVAL_1523;
  wire [14:0] _EVAL_1525;
  wire  _EVAL_1526;
  wire  _EVAL_1528;
  wire  _EVAL_1529;
  wire [31:0] _EVAL_1530;
  wire [11:0] _EVAL_1532;
  wire [1:0] _EVAL_1533;
  wire  _EVAL_1534;
  wire  _EVAL_1537;
  wire  _EVAL_1539;
  wire  _EVAL_1541;
  wire  _EVAL_1543;
  wire [7:0] _EVAL_1544;
  wire  _EVAL_1545;
  wire  _EVAL_1546;
  wire [7:0] _EVAL_1548;
  wire  _EVAL_1549;
  wire [4:0] _EVAL_1550;
  wire [142:0] _EVAL_1551;
  wire  _EVAL_1553;
  wire  _EVAL_1554;
  wire  _EVAL_1557;
  wire [31:0] _EVAL_1558;
  wire  _EVAL_1559;
  wire  _EVAL_1560;
  wire  _EVAL_1562;
  wire [142:0] _EVAL_1563;
  wire  _EVAL_1564;
  wire  _EVAL_1566;
  wire  _EVAL_1568;
  wire  _EVAL_1569;
  wire [7:0] _EVAL_1571;
  wire  _EVAL_1573;
  wire  _EVAL_1577;
  wire  _EVAL_1578;
  wire  _EVAL_1579;
  wire [142:0] _EVAL_1580;
  wire  _EVAL_1581;
  wire [6:0] _EVAL_1584;
  wire  _EVAL_1585;
  wire  _EVAL_1586;
  wire [32:0] _EVAL_1587;
  wire  _EVAL_1588;
  wire  _EVAL_1589;
  wire [142:0] _EVAL_1591;
  wire  _EVAL_1592;
  wire [31:0] _EVAL_1593;
  wire  _EVAL_1594;
  reg  _EVAL_1595;
  reg [31:0] _RAND_71;
  wire  _EVAL_1596;
  wire  _EVAL_1599;
  wire [31:0] _EVAL_1600;
  wire  _EVAL_1601;
  wire [31:0] _EVAL_1603;
  wire  _EVAL_1604;
  reg  _EVAL_1608;
  reg [31:0] _RAND_72;
  wire  _EVAL_1609;
  wire  _EVAL_1610;
  wire  _EVAL_1611;
  wire  _EVAL_1614;
  wire  _EVAL_1616;
  wire  _EVAL_1617;
  wire  _EVAL_1618;
  wire  _EVAL_1619;
  wire [1:0] _EVAL_1620;
  wire  _EVAL_1621;
  wire  _EVAL_1626;
  wire [7:0] _EVAL_1627;
  wire  _EVAL_1628;
  wire  _EVAL_1630;
  wire [7:0] _EVAL_1631;
  wire  _EVAL_1634;
  wire  _EVAL_1635;
  wire  _EVAL_1636;
  wire  _EVAL_1637;
  wire  _EVAL_1642;
  wire  _EVAL_1643;
  wire  _EVAL_1644;
  wire  _EVAL_1646;
  wire  _EVAL_1651;
  wire [7:0] _EVAL_1656;
  wire  _EVAL_1658;
  wire  _EVAL_1659;
  wire  _EVAL_1660;
  wire  _EVAL_1665;
  wire  _EVAL_1666;
  wire [32:0] _EVAL_1671;
  wire  _EVAL_1672;
  wire  _EVAL_1673;
  wire  _EVAL_1675;
  wire [1:0] _EVAL_1676;
  wire [3:0] _EVAL_1677;
  wire  _EVAL_1678;
  wire  _EVAL_1679;
  wire  _EVAL_1680;
  wire  _EVAL_1681;
  wire  _EVAL_1682;
  wire [9:0] _EVAL_1683;
  wire  _EVAL_1684;
  wire  _EVAL_1685;
  wire [16:0] _EVAL_1686;
  wire [7:0] _EVAL_1688;
  wire [142:0] _EVAL_1689;
  wire [1:0] _EVAL_1692;
  wire  _EVAL_1693;
  wire [3:0] _EVAL_1694;
  wire  _EVAL_1695;
  wire  _EVAL_1697;
  wire [5:0] _EVAL_1698;
  wire [142:0] _EVAL_1699;
  wire  _EVAL_1700;
  wire  _EVAL_1704;
  wire [7:0] _EVAL_1705;
  wire  _EVAL_1706;
  wire  _EVAL_1707;
  wire [7:0] _EVAL_1710;
  wire  _EVAL_1714;
  wire [6:0] _EVAL_1715;
  wire  _EVAL_1716;
  wire  _EVAL_1717;
  wire [7:0] _EVAL_1719;
  wire  _EVAL_1720;
  wire [39:0] _EVAL_1721;
  reg  _EVAL_1722;
  reg [31:0] _RAND_73;
  wire  _EVAL_1723;
  wire [7:0] _EVAL_1724;
  wire  _EVAL_1725;
  wire  _EVAL_1727;
  wire  _EVAL_1729;
  wire  _EVAL_1730;
  wire [4:0] _EVAL_1731;
  wire  _EVAL_1734;
  wire  _EVAL_1735;
  wire  _EVAL_1736;
  wire [63:0] _EVAL_1737;
  wire  _EVAL_1738;
  wire [31:0] _EVAL_1739;
  wire  _EVAL_1740;
  wire  _EVAL_1742;
  wire [6:0] _EVAL_1743;
  wire [4:0] _EVAL_1744;
  wire [5:0] _EVAL_1746;
  wire  _EVAL_1749;
  wire  _EVAL_1750;
  wire [31:0] _EVAL_1751;
  wire  _EVAL_1752;
  wire [142:0] _EVAL_1753;
  reg  _EVAL_1755;
  reg [31:0] _RAND_74;
  wire [7:0] _EVAL_1756;
  wire  _EVAL_1757;
  wire  _EVAL_1758;
  wire [6:0] _EVAL_1759;
  wire [7:0] _EVAL_1760;
  wire  _EVAL_1761;
  wire  _EVAL_1762;
  wire  _EVAL_1763;
  wire  _EVAL_1764;
  wire  _EVAL_1766;
  wire  _EVAL_1767;
  wire  _EVAL_1770;
  wire  _EVAL_1771;
  wire  _EVAL_1772;
  wire  _EVAL_1773;
  wire  _EVAL_1774;
  wire  _EVAL_1777;
  wire  _EVAL_1778;
  wire [142:0] _EVAL_1781;
  wire  _EVAL_1782;
  wire  _EVAL_1783;
  wire  _EVAL_1788;
  wire  _EVAL_1790;
  wire  _EVAL_1792;
  wire [31:0] _EVAL_1793;
  wire  _EVAL_1794;
  wire  _EVAL_1795;
  wire  _EVAL_1796;
  wire  _EVAL_1799;
  wire [3:0] _EVAL_1800;
  wire [31:0] _EVAL_1802;
  wire [31:0] _EVAL_1803;
  wire  _EVAL_1805;
  wire  _EVAL_1807;
  wire [10:0] _EVAL_1808;
  wire  _EVAL_1811;
  wire  _EVAL_1812;
  wire  _EVAL_1813;
  wire [102:0] _EVAL_1814;
  wire  _EVAL_1815;
  wire [31:0] _EVAL_1816;
  wire  _EVAL_1817;
  wire  _EVAL_1818;
  wire  _EVAL_1819;
  wire [31:0] _EVAL_1821;
  wire  _EVAL_1823;
  wire  _EVAL_1825;
  wire  _EVAL_1829;
  wire  _EVAL_1830;
  wire  _EVAL_1831;
  wire [4:0] _EVAL_1832;
  wire  _EVAL_1835;
  wire  _EVAL_1837;
  wire [7:0] _EVAL_1838;
  wire  _EVAL_1839;
  wire  _EVAL_1841;
  wire  _EVAL_1842;
  wire  _EVAL_1843;
  wire  _EVAL_1844;
  wire  _EVAL_1846;
  wire  _EVAL_1847;
  wire [7:0] _EVAL_1848;
  wire  _EVAL_1849;
  reg  _EVAL_1850;
  reg [31:0] _RAND_75;
  wire  _EVAL_1851;
  wire  _EVAL_1852;
  wire [7:0] _EVAL_1853;
  wire  _EVAL_1856;
  wire  _EVAL_1857;
  wire  _EVAL_1858;
  wire [31:0] _EVAL_1859;
  wire [1:0] _EVAL_1860;
  wire  _EVAL_1862;
  wire [30:0] _EVAL_1863;
  wire  _EVAL_1864;
  wire [6:0] _EVAL_1866;
  wire [3:0] _EVAL_1868;
  wire  _EVAL_1869;
  wire  _EVAL_1871;
  wire  _EVAL_1873;
  wire  _EVAL_1877;
  wire  _EVAL_1878;
  wire [31:0] _EVAL_1881;
  wire [63:0] _EVAL_1882;
  wire  _EVAL_1884;
  wire  _EVAL_1885;
  wire  _EVAL_1886;
  wire [1:0] _EVAL_1887;
  reg [2:0] _EVAL_1888;
  reg [31:0] _RAND_76;
  wire  _EVAL_1890;
  wire  _EVAL_1892;
  wire  _EVAL_1893;
  wire [31:0] _EVAL_1894;
  wire  _EVAL_1895;
  wire [1:0] _EVAL_1896;
  wire  _EVAL_1898;
  wire  _EVAL_1899;
  wire  _EVAL_1900;
  wire [63:0] _EVAL_1901;
  wire [31:0] _EVAL_1905;
  wire [7:0] _EVAL_1906;
  wire [1:0] _EVAL_1907;
  wire [31:0] _EVAL_1908;
  wire  _EVAL_1909;
  wire  _EVAL_1910;
  wire  _EVAL_1911;
  wire [31:0] _EVAL_1913;
  wire  _EVAL_1914;
  wire  _EVAL_1915;
  wire [31:0] _EVAL_1916;
  wire  _EVAL_1917;
  wire  _EVAL_1918;
  wire  _EVAL_1919;
  wire  _EVAL_1920;
  wire [142:0] _EVAL_1924;
  wire  _EVAL_1925;
  wire  _EVAL_1927;
  wire  _EVAL_1928;
  wire  _EVAL_1929;
  wire  _EVAL_1930;
  wire  _EVAL_1931;
  wire  _EVAL_1933;
  wire  _EVAL_1934;
  wire [63:0] _EVAL_1935;
  wire [1:0] _EVAL_1936;
  wire [7:0] _EVAL_1937;
  wire  _EVAL_1939;
  wire [31:0] _EVAL_1940;
  wire [58:0] _EVAL_1941;
  wire  _EVAL_1942;
  wire  _EVAL_1944;
  wire  _EVAL_1945;
  wire  _EVAL_1947;
  reg  _EVAL_1948;
  reg [31:0] _RAND_77;
  wire  _EVAL_1949;
  wire  _EVAL_1951;
  wire  _EVAL_1952;
  wire [29:0] _EVAL_1953;
  wire [7:0] _EVAL_1955;
  wire  _EVAL_1956;
  wire [31:0] _EVAL_1957;
  wire [142:0] _EVAL_1958;
  wire [1:0] _EVAL_1960;
  wire  _EVAL_1961;
  wire  _EVAL_1963;
  wire [6:0] _EVAL_1964;
  wire [6:0] _EVAL_1965;
  wire  _EVAL_1966;
  wire [142:0] _EVAL_1967;
  reg [33:0] _EVAL_1969;
  reg [63:0] _RAND_78;
  wire [5:0] _EVAL_1970;
  wire [30:0] _EVAL_1971;
  wire [31:0] _EVAL_1972;
  wire  _EVAL_1974;
  wire [6:0] _EVAL_1975;
  wire  _EVAL_1976;
  wire  _EVAL_1978;
  wire  _EVAL_1979;
  wire [5:0] _EVAL_1980;
  wire  _EVAL_1982;
  wire  _EVAL_1983;
  wire [6:0] _EVAL_1984;
  wire [142:0] _EVAL_1985;
  wire  _EVAL_1986;
  wire  _EVAL_1987;
  wire [31:0] _EVAL_1988;
  wire  _EVAL_1989;
  wire  _EVAL_1992;
  wire [142:0] _EVAL_1993;
  wire  _EVAL_1995;
  wire  _EVAL_1996;
  wire [31:0] _EVAL_1998;
  wire [31:0] _EVAL_1999;
  wire  _EVAL_2000;
  wire  _EVAL_2001;
  wire  _EVAL_2002;
  wire  _EVAL_2003;
  wire  _EVAL_2005;
  wire  _EVAL_2008;
  wire  _EVAL_2009;
  wire [7:0] _EVAL_2011;
  wire [142:0] _EVAL_2013;
  wire  _EVAL_2014;
  wire  _EVAL_2016;
  wire  _EVAL_2019;
  wire  _EVAL_2020;
  wire [7:0] _EVAL_2023;
  wire [5:0] _EVAL_2026;
  wire  _EVAL_2029;
  wire  _EVAL_2030;
  wire [1:0] _EVAL_2031;
  wire  _EVAL_2034;
  wire [39:0] _EVAL_2037;
  wire  _EVAL_2039;
  wire  _EVAL_2041;
  wire  _EVAL_2042;
  wire [7:0] _EVAL_2046;
  wire  _EVAL_2047;
  wire [7:0] _EVAL_2048;
  wire  _EVAL_2049;
  wire [31:0] _EVAL_2050;
  wire [31:0] _EVAL_2053;
  wire  _EVAL_2054;
  wire [7:0] _EVAL_2056;
  wire [7:0] _EVAL_2057;
  wire  _EVAL_2058;
  wire [7:0] _EVAL_2059;
  wire  _EVAL_2060;
  wire  _EVAL_2061;
  wire  _EVAL_2062;
  wire  _EVAL_2063;
  wire  _EVAL_2064;
  wire  _EVAL_2065;
  wire [7:0] _EVAL_2067;
  wire [6:0] _EVAL_2069;
  wire  _EVAL_2070;
  wire  _EVAL_2072;
  wire  _EVAL_2073;
  wire  _EVAL_2075;
  wire  _EVAL_2076;
  wire [31:0] _EVAL_2077;
  wire  _EVAL_2081;
  reg  _EVAL_2083;
  reg [31:0] _RAND_79;
  wire  _EVAL_2085;
  wire  _EVAL_2086;
  wire  _EVAL_2087;
  wire  _EVAL_2088;
  wire  _EVAL_2089;
  wire [7:0] _EVAL_2090;
  wire [7:0] _EVAL_2092;
  wire  _EVAL_2093;
  wire [142:0] _EVAL_2094;
  wire  _EVAL_2095;
  wire  _EVAL_2096;
  wire  _EVAL_2097;
  wire  _EVAL_2098;
  wire  _EVAL_2100;
  wire [31:0] _EVAL_2101;
  wire [31:0] _EVAL_2102;
  wire  _EVAL_2105;
  wire  _EVAL_2106;
  wire  _EVAL_2107;
  wire [31:0] _EVAL_2108;
  wire  _EVAL_2111;
  wire  _EVAL_2113;
  wire [6:0] _EVAL_2114;
  wire [142:0] _EVAL_2115;
  wire  _EVAL_2117;
  wire  _EVAL_2118;
  wire [31:0] _EVAL_2119;
  wire  _EVAL_2121;
  wire [5:0] _EVAL_2122;
  wire  _EVAL_2123;
  wire  _EVAL_2124;
  wire [142:0] _EVAL_2125;
  wire  _EVAL_2127;
  wire [7:0] _EVAL_2128;
  reg  _EVAL_2129;
  reg [31:0] _RAND_80;
  wire  _EVAL_2130;
  wire  _EVAL_2133;
  wire  _EVAL_2134;
  wire  _EVAL_2135;
  wire  _EVAL_2138;
  wire  _EVAL_2139;
  wire  _EVAL_2141;
  wire  _EVAL_2142;
  wire  _EVAL_2145;
  wire  _EVAL_2146;
  reg [1:0] _EVAL_2147;
  reg [31:0] _RAND_81;
  reg  _EVAL_2148;
  reg [31:0] _RAND_82;
  wire  _EVAL_2149;
  wire [31:0] _EVAL_2150;
  wire  _EVAL_2151;
  wire [142:0] _EVAL_2152;
  wire [6:0] _EVAL_2155;
  wire [7:0] _EVAL_2156;
  wire  _EVAL_2157;
  reg  _EVAL_2158;
  reg [31:0] _RAND_83;
  wire [31:0] _EVAL_2159;
  wire [7:0] _EVAL_2160;
  wire  _EVAL_2161;
  wire [6:0] _EVAL_2162;
  wire  _EVAL_2163;
  wire  _EVAL_2164;
  wire  _EVAL_2165;
  wire  _EVAL_2166;
  wire [31:0] _EVAL_2168;
  wire [7:0] _EVAL_2169;
  wire  _EVAL_2170;
  wire [6:0] _EVAL_2171;
  wire  _EVAL_2172;
  wire [5:0] _EVAL_2173;
  wire  _EVAL_2175;
  wire [6:0] _EVAL_2178;
  wire  _EVAL_2179;
  wire  _EVAL_2182;
  wire  _EVAL_2184;
  wire [30:0] _EVAL_2185;
  wire  _EVAL_2186;
  wire [5:0] _EVAL_2188;
  wire  _EVAL_2189;
  wire [31:0] _EVAL_2190;
  wire [31:0] _EVAL_2191;
  wire  _EVAL_2192;
  wire  _EVAL_2193;
  wire [31:0] _EVAL_2195;
  wire  _EVAL_2196;
  wire  _EVAL_2199;
  wire [7:0] _EVAL_2201;
  wire [142:0] _EVAL_2202;
  wire  _EVAL_2203;
  wire [31:0] _EVAL_2204;
  wire  _EVAL_2205;
  wire  _EVAL_2206;
  wire  _EVAL_2208;
  wire  _EVAL_2209;
  wire  _EVAL_2210;
  wire [16:0] _EVAL_2211;
  wire [142:0] _EVAL_2213;
  wire [4:0] _EVAL_2215;
  wire  _EVAL_2216;
  wire  _EVAL_2217;
  wire  _EVAL_2218;
  wire  _EVAL_2219;
  wire  _EVAL_2221;
  wire [4:0] _EVAL_2222;
  wire  _EVAL_2223;
  wire [7:0] _EVAL_2224;
  wire  _EVAL_2225;
  wire  _EVAL_2227;
  wire  _EVAL_2228;
  wire  _EVAL_2229;
  wire  _EVAL_2231;
  wire  _EVAL_2233;
  wire  _EVAL_2234;
  wire  _EVAL_2235;
  wire  _EVAL_2236;
  wire [6:0] _EVAL_2239;
  wire [32:0] _EVAL_2241;
  wire  _EVAL_2247;
  wire  _EVAL_2248;
  wire  _EVAL_2250;
  reg [7:0] _EVAL_2251;
  reg [31:0] _RAND_84;
  wire  _EVAL_2252;
  wire  _EVAL_2255;
  wire  _EVAL_2256;
  wire  _EVAL_2257;
  wire [31:0] _EVAL_2258;
  wire [31:0] _EVAL_2260;
  wire  _EVAL_2261;
  wire  _EVAL_2262;
  wire  _EVAL_2263;
  wire  _EVAL_2264;
  wire  _EVAL_2265;
  wire [31:0] _EVAL_2267;
  reg  _EVAL_2268;
  reg [31:0] _RAND_85;
  wire [7:0] _EVAL_2269;
  wire  _EVAL_2271;
  wire  _EVAL_2274;
  wire  _EVAL_2276;
  wire  _EVAL_2277;
  wire  _EVAL_2278;
  wire [7:0] _EVAL_2279;
  wire [10:0] _EVAL_2280;
  wire [31:0] _EVAL_2281;
  wire [7:0] _EVAL_2284;
  wire  _EVAL_2285;
  wire [7:0] _EVAL_2286;
  wire  _EVAL_2287;
  wire  _EVAL_2289;
  wire  _EVAL_2290;
  wire  _EVAL_2293;
  wire  _EVAL_2294;
  wire  _EVAL_2295;
  wire [7:0] _EVAL_2296;
  wire [142:0] _EVAL_2297;
  wire  _EVAL_2298;
  wire  _EVAL_2299;
  wire [7:0] _EVAL_2300;
  wire  _EVAL_2302;
  wire [57:0] _EVAL_2304;
  wire  _EVAL_2305;
  reg [31:0] _EVAL_2306;
  reg [31:0] _RAND_86;
  wire  _EVAL_2308;
  wire [142:0] _EVAL_2309;
  wire  _EVAL_2310;
  wire [7:0] _EVAL_2311;
  wire  _EVAL_2314;
  wire [57:0] _EVAL_2315;
  wire [39:0] _EVAL_2317;
  wire  _EVAL_2318;
  wire  _EVAL_2319;
  wire  _EVAL_2320;
  wire  _EVAL_2321;
  wire [7:0] _EVAL_2322;
  wire  _EVAL_2323;
  wire  _EVAL_2324;
  wire [6:0] _EVAL_2325;
  wire  _EVAL_2326;
  wire  _EVAL_2327;
  wire  _EVAL_2330;
  wire  _EVAL_2333;
  wire  _EVAL_2335;
  wire [6:0] _EVAL_2338;
  wire [6:0] _EVAL_2340;
  wire [29:0] _EVAL_2342;
  wire  _EVAL_2343;
  wire [6:0] _EVAL_2344;
  wire  _EVAL_2345;
  wire  _EVAL_2346;
  wire  _EVAL_2347;
  wire  _EVAL_2348;
  reg  _EVAL_2349;
  reg [31:0] _RAND_87;
  wire  _EVAL_2350;
  wire  _EVAL_2351;
  wire [31:0] _EVAL_2352;
  wire  _EVAL_2354;
  reg [2:0] _EVAL_2355;
  reg [31:0] _RAND_88;
  reg  _EVAL_2356;
  reg [31:0] _RAND_89;
  wire [142:0] _EVAL_2358;
  wire  _EVAL_2359;
  wire  _EVAL_2360;
  wire  _EVAL_2362;
  wire [7:0] _EVAL_2363;
  wire  _EVAL_2364;
  wire  _EVAL_2366;
  wire  _EVAL_2367;
  wire [31:0] _EVAL_2369;
  wire  _EVAL_2372;
  wire [31:0] _EVAL_2374;
  reg  _EVAL_2375;
  reg [31:0] _RAND_90;
  wire  _EVAL_2376;
  wire  _EVAL_2378;
  wire [6:0] _EVAL_2379;
  reg  _EVAL_2380;
  reg [31:0] _RAND_91;
  wire  _EVAL_2381;
  wire  _EVAL_2382;
  wire [7:0] _EVAL_2384;
  wire  _EVAL_2385;
  wire  _EVAL_2386;
  reg  _EVAL_2387;
  reg [31:0] _RAND_92;
  wire [142:0] _EVAL_2388;
  wire  _EVAL_2389;
  wire  _EVAL_2391;
  reg [1:0] _EVAL_2392;
  reg [31:0] _RAND_93;
  wire  _EVAL_2394;
  wire  _EVAL_2395;
  wire  _EVAL_2396;
  wire  _EVAL_2397;
  wire  _EVAL_2400;
  wire  _EVAL_2404;
  wire [31:0] _EVAL_2405;
  reg  _EVAL_2406;
  reg [31:0] _RAND_94;
  wire  _EVAL_2407;
  wire [142:0] _EVAL_2408;
  wire  _EVAL_2409;
  wire  _EVAL_2410;
  wire  _EVAL_2411;
  wire [31:0] _EVAL_2413;
  wire  _EVAL_2414;
  wire  _EVAL_2416;
  wire  _EVAL_2418;
  wire [7:0] _EVAL_2419;
  wire  _EVAL_2420;
  wire  _EVAL_2421;
  wire  _EVAL_2422;
  wire  _EVAL_2423;
  wire  _EVAL_2425;
  wire  _EVAL_2427;
  wire  _EVAL_2428;
  wire  _EVAL_2429;
  wire  _EVAL_2430;
  wire  _EVAL_2431;
  wire  _EVAL_2433;
  wire  _EVAL_2434;
  wire [1:0] _EVAL_2435;
  wire [5:0] _EVAL_2440;
  wire [7:0] _EVAL_2441;
  wire  _EVAL_2442;
  wire  _EVAL_2443;
  wire [7:0] _EVAL_2444;
  reg [1:0] _EVAL_2445;
  reg [31:0] _RAND_95;
  wire [7:0] _EVAL_2446;
  wire [7:0] _EVAL_2447;
  wire [7:0] _EVAL_2448;
  wire  _EVAL_2449;
  wire [6:0] _EVAL_2451;
  wire  _EVAL_2452;
  wire  _EVAL_2453;
  wire  _EVAL_2454;
  wire [31:0] _EVAL_2455;
  wire  _EVAL_2457;
  wire  _EVAL_2458;
  wire  _EVAL_2460;
  wire  _EVAL_2461;
  wire  _EVAL_2462;
  wire  _EVAL_2463;
  wire [18:0] _EVAL_2464;
  wire  _EVAL_2466;
  wire  _EVAL_2467;
  wire  _EVAL_2468;
  wire  _EVAL_2469;
  wire  _EVAL_2470;
  reg [1:0] _EVAL_2471;
  reg [31:0] _RAND_96;
  wire  _EVAL_2472;
  wire  _EVAL_2474;
  wire  _EVAL_2477;
  reg [9:0] _EVAL_2479;
  reg [31:0] _RAND_97;
  wire [3:0] _EVAL_2480;
  wire  _EVAL_2481;
  wire  _EVAL_2482;
  wire  _EVAL_2484;
  wire  _EVAL_2485;
  reg  _EVAL_2486;
  reg [31:0] _RAND_98;
  wire  _EVAL_2487;
  wire [7:0] _EVAL_2488;
  wire [31:0] _EVAL_2489;
  wire  _EVAL_2490;
  wire  _EVAL_2492;
  wire  _EVAL_2493;
  wire [6:0] _EVAL_2494;
  wire  _EVAL_2495;
  wire  _EVAL_2496;
  wire [11:0] _EVAL_2498;
  wire  _EVAL_2500;
  wire  _EVAL_2501;
  wire  _EVAL_2502;
  wire  _EVAL_2504;
  wire  _EVAL_2505;
  wire  _EVAL_2506;
  wire [31:0] _EVAL_2507;
  wire [7:0] _EVAL_2508;
  wire  _EVAL_2509;
  wire [142:0] _EVAL_2510;
  wire  _EVAL_2511;
  wire  _EVAL_2513;
  wire [63:0] _EVAL_2516;
  wire [31:0] _EVAL_2517;
  wire  _EVAL_2519;
  wire  _EVAL_2521;
  wire  _EVAL_2524;
  wire [7:0] _EVAL_2525;
  wire [1:0] _EVAL_2527;
  wire [142:0] _EVAL_2528;
  wire [7:0] _EVAL_2529;
  wire  _EVAL_2533;
  wire  _EVAL_2534;
  wire  _EVAL_2535;
  wire  _EVAL_2536;
  wire  _EVAL_2537;
  wire  _EVAL_2538;
  wire  _EVAL_2539;
  wire  _EVAL_2540;
  wire  _EVAL_2541;
  reg  _EVAL_2542;
  reg [31:0] _RAND_99;
  wire  _EVAL_2543;
  wire  _EVAL_2544;
  wire [31:0] _EVAL_2545;
  wire [142:0] _EVAL_2546;
  wire  _EVAL_2548;
  wire [142:0] _EVAL_2549;
  wire [31:0] _EVAL_2550;
  wire [142:0] _EVAL_2551;
  wire  _EVAL_2557;
  wire  _EVAL_2558;
  wire  _EVAL_2561;
  wire [1:0] _EVAL_2562;
  wire [25:0] _EVAL_2563;
  wire [6:0] _EVAL_2564;
  wire  _EVAL_2567;
  wire  _EVAL_2568;
  wire  _EVAL_2569;
  wire  _EVAL_2571;
  wire [31:0] _EVAL_2573;
  wire  _EVAL_2574;
  reg  _EVAL_2579;
  reg [31:0] _RAND_100;
  wire  _EVAL_2580;
  wire  _EVAL_2581;
  wire  _EVAL_2582;
  wire [7:0] _EVAL_2583;
  wire  _EVAL_2584;
  wire [7:0] _EVAL_2586;
  wire  _EVAL_2587;
  wire  _EVAL_2588;
  wire  _EVAL_2589;
  wire [7:0] _EVAL_2590;
  wire  _EVAL_2591;
  wire  _EVAL_2592;
  reg  _EVAL_2593;
  reg [31:0] _RAND_101;
  wire  _EVAL_2594;
  wire [6:0] _EVAL_2595;
  wire [5:0] _EVAL_2597;
  wire  _EVAL_2599;
  wire  _EVAL_2602;
  wire  _EVAL_2604;
  wire [31:0] _EVAL_2605;
  wire  _EVAL_2606;
  wire  _EVAL_2607;
  wire [5:0] _EVAL_2608;
  reg [1:0] _EVAL_2609;
  reg [31:0] _RAND_102;
  wire [11:0] _EVAL_2611;
  wire [142:0] _EVAL_2613;
  wire [31:0] _EVAL_2614;
  wire  _EVAL_2615;
  wire [31:0] _EVAL_2616;
  wire [5:0] _EVAL_2617;
  wire  _EVAL_2620;
  wire  _EVAL_2621;
  wire [7:0] _EVAL_2622;
  wire [7:0] _EVAL_2624;
  wire [7:0] _EVAL_2627;
  wire  _EVAL_2628;
  wire  _EVAL_2629;
  wire [4:0] _EVAL_2631;
  wire  _EVAL_2632;
  wire  _EVAL_2636;
  wire  _EVAL_2637;
  wire [142:0] _EVAL_2638;
  wire [31:0] _EVAL_2640;
  reg [5:0] _EVAL_2644;
  reg [31:0] _RAND_103;
  wire [6:0] _EVAL_2645;
  reg  _EVAL_2647;
  reg [31:0] _RAND_104;
  wire [6:0] _EVAL_2648;
  wire [5:0] _EVAL_2649;
  wire  _EVAL_2650;
  wire [31:0] _EVAL_2651;
  wire [7:0] _EVAL_2652;
  wire  _EVAL_2653;
  reg  _EVAL_2654;
  reg [31:0] _RAND_105;
  wire  _EVAL_2655;
  wire [5:0] _EVAL_2656;
  wire  _EVAL_2657;
  wire  _EVAL_2658;
  wire  _EVAL_2659;
  wire  _EVAL_2660;
  wire [142:0] _EVAL_2661;
  wire [6:0] _EVAL_2662;
  wire  _EVAL_2663;
  reg [23:0] _EVAL_2665;
  reg [31:0] _RAND_106;
  wire  _EVAL_2666;
  wire [31:0] _EVAL_2667;
  wire  _EVAL_2668;
  wire  _EVAL_2669;
  wire  _EVAL_2670;
  wire [7:0] _EVAL_2671;
  reg  _EVAL_2673;
  reg [31:0] _RAND_107;
  reg  _EVAL_2674;
  reg [31:0] _RAND_108;
  reg  _EVAL_2676;
  reg [31:0] _RAND_109;
  wire [34:0] _EVAL_2677;
  wire  _EVAL_2678;
  wire  _EVAL_2680;
  wire  _EVAL_2681;
  wire  _EVAL_2685;
  wire  _EVAL_2688;
  reg [31:0] _EVAL_2689;
  reg [31:0] _RAND_110;
  wire [7:0] _EVAL_2690;
  wire [7:0] _EVAL_2691;
  wire [5:0] _EVAL_2692;
  wire  _EVAL_2694;
  wire  _EVAL_2695;
  wire  _EVAL_2696;
  wire  _EVAL_2697;
  wire  _EVAL_2698;
  wire [1:0] _EVAL_2699;
  wire  _EVAL_2701;
  wire [30:0] _EVAL_2702;
  wire [142:0] _EVAL_2703;
  wire  _EVAL_2704;
  wire [57:0] _EVAL_2705;
  wire  _EVAL_2707;
  reg [1:0] _EVAL_2708;
  reg [31:0] _RAND_111;
  wire  _EVAL_2709;
  wire  _EVAL_2711;
  wire  _EVAL_2712;
  wire [31:0] _EVAL_2713;
  wire [4:0] _EVAL_2715;
  wire  _EVAL_2716;
  wire  _EVAL_2717;
  wire [31:0] _EVAL_2719;
  wire  _EVAL_2720;
  wire [3:0] _EVAL_2722;
  wire  _EVAL_2725;
  wire [31:0] _EVAL_2727;
  wire  _EVAL_2728;
  wire  _EVAL_2729;
  wire [142:0] _EVAL_2730;
  wire  _EVAL_2731;
  reg [1:0] _EVAL_2732;
  reg [31:0] _RAND_112;
  wire  _EVAL_2733;
  wire [7:0] _EVAL_2735;
  wire  _EVAL_2736;
  wire  _EVAL_2737;
  wire [7:0] _EVAL_2738;
  wire [31:0] _EVAL_2740;
  wire  _EVAL_2741;
  wire  _EVAL_2743;
  wire  _EVAL_2744;
  wire  _EVAL_2746;
  wire  _EVAL_2747;
  wire  _EVAL_2748;
  wire  _EVAL_2750;
  wire [6:0] _EVAL_2752;
  wire [6:0] _EVAL_2753;
  wire  _EVAL_2754;
  wire [7:0] _EVAL_2755;
  wire  _EVAL_2757;
  wire  _EVAL_2760;
  wire  _EVAL_2761;
  reg  _EVAL_2764;
  reg [31:0] _RAND_113;
  wire [15:0] _EVAL_2766;
  wire  _EVAL_2767;
  wire [31:0] _EVAL_2769;
  wire [3:0] _EVAL_2770;
  wire  _EVAL_2771;
  wire  _EVAL_2772;
  wire  _EVAL_2774;
  wire [4:0] _EVAL_2775;
  wire  _EVAL_2778;
  wire  _EVAL_2779;
  reg  _EVAL_2784;
  reg [31:0] _RAND_114;
  wire  _EVAL_2786;
  wire [7:0] _EVAL_2787;
  wire  _EVAL_2788;
  wire  _EVAL_2789;
  wire [7:0] _EVAL_2790;
  reg [1:0] _EVAL_2791;
  reg [31:0] _RAND_115;
  wire  _EVAL_2792;
  wire  _EVAL_2793;
  wire  _EVAL_2794;
  wire  _EVAL_2796;
  reg [29:0] _EVAL_2799;
  reg [31:0] _RAND_116;
  wire  _EVAL_2802;
  wire [5:0] _EVAL_2803;
  wire  _EVAL_2804;
  wire  _EVAL_2805;
  wire  _EVAL_2806;
  wire  _EVAL_2808;
  wire  _EVAL_2809;
  wire  _EVAL_2810;
  wire  _EVAL_2813;
  wire [1:0] _EVAL_2814;
  wire  _EVAL_2815;
  wire  _EVAL_2817;
  wire  _EVAL_2818;
  wire  _EVAL_2819;
  wire [7:0] _EVAL_2821;
  wire [142:0] _EVAL_2822;
  wire  _EVAL_2823;
  wire  _EVAL_2824;
  wire  _EVAL_2827;
  reg [15:0] _EVAL_2828;
  reg [31:0] _RAND_117;
  wire  _EVAL_2830;
  wire  _EVAL_2831;
  wire [6:0] _EVAL_2833;
  wire [7:0] _EVAL_2834;
  wire [142:0] _EVAL_2836;
  wire  _EVAL_2837;
  wire  _EVAL_2838;
  wire [57:0] _EVAL_2841;
  reg  _EVAL_2842;
  reg [31:0] _RAND_118;
  wire [1:0] _EVAL_2843;
  reg  _EVAL_2844;
  reg [31:0] _RAND_119;
  wire  _EVAL_2845;
  wire  _EVAL_2846;
  wire  _EVAL_2848;
  wire  _EVAL_2849;
  wire  _EVAL_2850;
  wire  _EVAL_2851;
  wire  _EVAL_2853;
  wire [7:0] _EVAL_2856;
  wire  _EVAL_2857;
  wire [7:0] _EVAL_2858;
  wire [5:0] _EVAL_2859;
  wire [142:0] _EVAL_2861;
  wire [31:0] _EVAL_2862;
  wire  _EVAL_2863;
  wire  _EVAL_2865;
  wire  _EVAL_2866;
  wire [30:0] _EVAL_2867;
  wire  _EVAL_2868;
  wire  _EVAL_2869;
  reg [31:0] _EVAL_2870;
  reg [31:0] _RAND_120;
  wire [31:0] _EVAL_2872;
  wire [31:0] _EVAL_2873;
  wire [6:0] _EVAL_2875;
  wire  _EVAL_2876;
  wire  _EVAL_2877;
  wire  _EVAL_2878;
  wire [31:0] _EVAL_2880;
  wire  _EVAL_2881;
  wire  _EVAL_2884;
  wire  _EVAL_2887;
  wire [31:0] _EVAL_2888;
  wire  _EVAL_2889;
  wire  _EVAL_2890;
  wire [7:0] _EVAL_2893;
  wire [7:0] _EVAL_2895;
  wire [31:0] _EVAL_2896;
  wire  _EVAL_2898;
  wire  _EVAL_2899;
  wire  _EVAL_2900;
  wire [142:0] _EVAL_2901;
  wire [7:0] _EVAL_2902;
  wire  _EVAL_2903;
  wire  _EVAL_2904;
  wire [142:0] _EVAL_2906;
  reg  _EVAL_2907;
  reg [31:0] _RAND_121;
  wire [31:0] _EVAL_2908;
  wire  _EVAL_2909;
  wire [31:0] _EVAL_2913;
  reg [1:0] _EVAL_2914;
  reg [31:0] _RAND_122;
  wire  _EVAL_2915;
  wire  _EVAL_2917;
  wire [57:0] _EVAL_2918;
  wire  _EVAL_2920;
  reg  _EVAL_2927;
  reg [31:0] _RAND_123;
  wire  _EVAL_2928;
  wire  _EVAL_2929;
  reg [31:0] _EVAL_2931;
  reg [31:0] _RAND_124;
  wire  _EVAL_2933;
  wire  _EVAL_2934;
  wire [39:0] _EVAL_2937;
  wire  _EVAL_2939;
  wire [142:0] _EVAL_2940;
  wire  _EVAL_2941;
  wire [142:0] _EVAL_2942;
  wire  _EVAL_2944;
  wire  _EVAL_2945;
  wire [7:0] _EVAL_2946;
  wire  _EVAL_2949;
  wire  _EVAL_2950;
  wire [31:0] _EVAL_2951;
  wire  _EVAL_2953;
  wire  _EVAL_2954;
  wire  _EVAL_2955;
  wire [63:0] _EVAL_2956;
  wire  _EVAL_2958;
  wire  _EVAL_2960;
  wire [142:0] _EVAL_2962;
  wire  _EVAL_2964;
  wire  _EVAL_2965;
  wire [31:0] _EVAL_2966;
  wire  _EVAL_2968;
  wire [7:0] _EVAL_2970;
  wire [142:0] _EVAL_2971;
  wire  _EVAL_2972;
  wire  _EVAL_2974;
  wire  _EVAL_2975;
  wire [7:0] _EVAL_2976;
  wire  _EVAL_2977;
  wire  _EVAL_2978;
  wire [7:0] _EVAL_2981;
  wire  _EVAL_2983;
  wire  _EVAL_2985;
  wire  _EVAL_2986;
  reg [1:0] _EVAL_2987;
  reg [31:0] _RAND_125;
  wire  _EVAL_2988;
  wire [7:0] _EVAL_2989;
  wire [142:0] _EVAL_2990;
  wire  _EVAL_2991;
  wire [63:0] _EVAL_2993;
  wire [7:0] _EVAL_2994;
  wire [7:0] _EVAL_2996;
  wire  _EVAL_2998;
  wire [31:0] _EVAL_2999;
  wire  _EVAL_3000;
  wire  _EVAL_3002;
  wire  _EVAL_3005;
  wire [31:0] _EVAL_3006;
  wire  _EVAL_3007;
  wire  _EVAL_3008;
  wire [2:0] _EVAL_3011;
  wire [31:0] _EVAL_3012;
  wire  _EVAL_3013;
  wire  _EVAL_3014;
  wire [7:0] _EVAL_3015;
  wire  _EVAL_3016;
  wire  _EVAL_3018;
  wire [63:0] _EVAL_3020;
  wire [7:0] _EVAL_3021;
  wire  _EVAL_3022;
  wire  _EVAL_3025;
  wire [142:0] _EVAL_3026;
  wire  _EVAL_3027;
  wire [3:0] _EVAL_3029;
  wire  _EVAL_3031;
  wire  _EVAL_3033;
  wire  _EVAL_3034;
  wire [6:0] _EVAL_3035;
  wire  _EVAL_3036;
  wire  _EVAL_3037;
  wire [31:0] _EVAL_3040;
  wire [31:0] _EVAL_3042;
  wire [39:0] _EVAL_3043;
  wire [58:0] _EVAL_3044;
  wire  _EVAL_3046;
  wire  _EVAL_3048;
  wire [31:0] _EVAL_3049;
  wire [7:0] _EVAL_3051;
  reg  _EVAL_3052;
  reg [31:0] _RAND_126;
  wire [31:0] _EVAL_3053;
  wire [5:0] _EVAL_3055;
  wire  _EVAL_3057;
  reg  _EVAL_3058;
  reg [31:0] _RAND_127;
  wire  _EVAL_3059;
  wire  _EVAL_3060;
  wire [142:0] _EVAL_3062;
  wire  _EVAL_3063;
  wire [6:0] _EVAL_3064;
  wire  _EVAL_3065;
  wire [5:0] _EVAL_3066;
  wire [7:0] _EVAL_3067;
  reg [1:0] _EVAL_3068;
  reg [31:0] _RAND_128;
  wire  _EVAL_3069;
  reg [5:0] _EVAL_3070;
  reg [31:0] _RAND_129;
  wire  _EVAL_3074;
  wire  _EVAL_3075;
  wire [31:0] _EVAL_3076;
  wire [30:0] _EVAL_3078;
  wire [1:0] _EVAL_3079;
  wire [31:0] _EVAL_3080;
  wire  _EVAL_3081;
  wire [6:0] _EVAL_3082;
  wire [1:0] _EVAL_3084;
  wire [6:0] _EVAL_3086;
  wire [4:0] _EVAL_3087;
  wire  _EVAL_3088;
  wire [31:0] _EVAL_3089;
  wire  _EVAL_3090;
  wire  _EVAL_3091;
  wire [5:0] _EVAL_3095;
  wire [7:0] _EVAL_3096;
  wire  _EVAL_3097;
  wire  _EVAL_3099;
  wire [30:0] _EVAL_3100;
  wire [5:0] _EVAL_3101;
  wire  _EVAL_3102;
  wire  _EVAL_3105;
  wire  _EVAL_3106;
  wire  _EVAL_3109;
  wire [31:0] _EVAL_3110;
  wire [32:0] _EVAL_3112;
  wire [31:0] _EVAL_3113;
  wire  _EVAL_3114;
  reg  _EVAL_3115;
  reg [31:0] _RAND_130;
  wire [1:0] _EVAL_3116;
  wire  _EVAL_3117;
  wire [142:0] _EVAL_3119;
  wire [6:0] _EVAL_3120;
  wire  _EVAL_3121;
  wire [7:0] _EVAL_3122;
  wire  _EVAL_3123;
  wire  _EVAL_3125;
  wire  _EVAL_3127;
  wire  _EVAL_3128;
  wire [31:0] _EVAL_3129;
  wire [7:0] _EVAL_3131;
  wire  _EVAL_3133;
  wire  _EVAL_3134;
  wire  _EVAL_3136;
  wire  _EVAL_3139;
  wire  _EVAL_3140;
  reg  _EVAL_3143;
  reg [31:0] _RAND_131;
  wire [31:0] _EVAL_3144;
  wire  _EVAL_3147;
  wire  _EVAL_3148;
  wire  _EVAL_3149;
  wire  _EVAL_3150;
  reg [30:0] _EVAL_3152;
  reg [31:0] _RAND_132;
  wire  _EVAL_3153;
  wire  _EVAL_3156;
  wire  _EVAL_3157;
  wire  _EVAL_3158;
  wire [31:0] _EVAL_3160;
  wire [5:0] _EVAL_3162;
  wire  _EVAL_3163;
  wire  _EVAL_3164;
  wire  _EVAL_3165;
  wire  _EVAL_3166;
  wire  _EVAL_3167;
  wire [6:0] _EVAL_3168;
  wire  _EVAL_3169;
  reg [1:0] _EVAL_3170;
  reg [31:0] _RAND_133;
  wire [7:0] _EVAL_3171;
  wire  _EVAL_3172;
  wire  _EVAL_3173;
  wire [142:0] _EVAL_3175;
  wire  _EVAL_3179;
  wire  _EVAL_3180;
  wire [10:0] _EVAL_3181;
  wire  _EVAL_3182;
  reg  _EVAL_3183;
  reg [31:0] _RAND_134;
  reg [31:0] _EVAL_3184;
  reg [31:0] _RAND_135;
  wire  _EVAL_3186;
  wire  _EVAL_3187;
  wire  _EVAL_3189;
  wire  _EVAL_3193;
  wire  _EVAL_3194;
  reg [1:0] _EVAL_3195;
  reg [31:0] _RAND_136;
  wire  _EVAL_3196;
  wire [7:0] _EVAL_3197;
  wire  _EVAL_3198;
  wire  _EVAL_3199;
  wire [5:0] _EVAL_3201;
  wire  _EVAL_3202;
  wire  _EVAL_3203;
  wire  _EVAL_3206;
  wire  _EVAL_3207;
  wire  _EVAL_3208;
  wire  _EVAL_3209;
  wire  _EVAL_3210;
  reg  _EVAL_3213;
  reg [31:0] _RAND_137;
  wire  _EVAL_3214;
  wire  _EVAL_3215;
  wire [7:0] _EVAL_3216;
  reg  _EVAL_3217;
  reg [31:0] _RAND_138;
  wire  _EVAL_3218;
  wire  _EVAL_3219;
  wire  _EVAL_3224;
  wire [142:0] _EVAL_3225;
  wire  _EVAL_3228;
  wire  _EVAL_3229;
  reg [1:0] _EVAL_3231;
  reg [31:0] _RAND_139;
  wire [31:0] _EVAL_3233;
  wire  _EVAL_3235;
  wire  _EVAL_3236;
  wire  _EVAL_3237;
  reg [57:0] _EVAL_3239;
  reg [63:0] _RAND_140;
  reg  _EVAL_3242;
  reg [31:0] _RAND_141;
  wire  _EVAL_3243;
  wire  _EVAL_3245;
  wire  _EVAL_3246;
  wire  _EVAL_3248;
  wire  _EVAL_3249;
  wire  _EVAL_3250;
  wire [6:0] _EVAL_3251;
  wire [31:0] _EVAL_3254;
  reg [5:0] _EVAL_3256;
  reg [31:0] _RAND_142;
  assign _EVAL_2856 = _EVAL_1106 ? 8'h8 : _EVAL_1152;
  assign _EVAL_1113 = _EVAL_1611 | _EVAL_613;
  assign _EVAL_2 = _EVAL_2927;
  assign _EVAL_3162 = _EVAL_2319 ? 6'h37 : _EVAL_298;
  assign _EVAL_1835 = _EVAL_76 == 12'h3bb;
  assign _EVAL_151 = _EVAL_76[11:10];
  assign _EVAL_1630 = _EVAL_2659 & _EVAL_1790;
  assign _EVAL_3043 = {_EVAL_1906,_EVAL_2258};
  assign _EVAL_1282 = _EVAL_2298 | _EVAL_2175;
  assign _EVAL_2089 = _EVAL_76 == 12'h300;
  assign _EVAL_2118 = _EVAL_3090 | _EVAL_937;
  assign _EVAL_432 = _EVAL_176 | _EVAL_882;
  assign _EVAL_500 = _EVAL_640 | _EVAL_1707;
  assign _EVAL_2290 = _EVAL_76 == 12'hc92;
  assign _EVAL_282 = _EVAL_1187[63:6];
  assign _EVAL_572 = {{142'd0}, _EVAL_1134};
  assign _EVAL_772 = {{71'd0}, _EVAL_2258};
  assign _EVAL_736 = _EVAL_76 == 12'h325;
  assign _EVAL_430 = _EVAL_923 | _EVAL_327;
  assign _EVAL_67 = _EVAL_1450;
  assign _EVAL_1814 = {_EVAL_123,_EVAL_103,_EVAL_131,_EVAL_47,_EVAL_129,_EVAL_116,_EVAL_31,_EVAL_125,_EVAL_2211,_EVAL_2464};
  assign _EVAL_2039 = _EVAL_3189 & _EVAL_526;
  assign _EVAL_74 = _EVAL_2129;
  assign _EVAL_1706 = _EVAL_1095 & _EVAL_2524;
  assign _EVAL_2850 = _EVAL_1231 | _EVAL_769;
  assign _EVAL_1286 = _EVAL_1992 | _EVAL_1036;
  assign _EVAL_115 = _EVAL_891;
  assign _EVAL_2474 = _EVAL_76 == 12'hc80;
  assign _EVAL_168 = _EVAL_2605[31:2];
  assign _EVAL_123 = _EVAL_2647;
  assign _EVAL_1852 = _EVAL_2850 | _EVAL_1106;
  assign _EVAL_660 = _EVAL_2673 | _EVAL_1685;
  assign _EVAL_810 = _EVAL_776[56];
  assign _EVAL_2945 = _EVAL_1259 | _EVAL_2513;
  assign _EVAL_1890 = _EVAL_2013[93];
  assign _EVAL_1236 = _EVAL_1846 & _EVAL_473;
  assign _EVAL_90 = _EVAL_1239;
  assign _EVAL_1526 = _EVAL_975 | _EVAL_1396;
  assign _EVAL_742 = _EVAL_1774 | _EVAL_540;
  assign _EVAL_1058 = _EVAL_1171 ? 8'h57 : _EVAL_2444;
  assign _EVAL_328 = _EVAL_76 == 12'h7a1;
  assign _EVAL_1026 = _EVAL_2697 & _EVAL_1050;
  assign _EVAL_927 = _EVAL_526 | _EVAL_2647;
  assign _EVAL_3219 = _EVAL_1717 & _EVAL_452;
  assign _EVAL_2790 = _EVAL_1090 ? 8'h3e : _EVAL_981;
  assign _EVAL_471 = _EVAL_1001 | _EVAL_367;
  assign _EVAL_1544 = _EVAL_1362 ? 8'h4a : _EVAL_1359;
  assign _EVAL_1771 = _EVAL_108 > _EVAL_1267;
  assign _EVAL_686 = _EVAL_2636 | _EVAL_2416;
  assign _EVAL_140 = _EVAL_2268;
  assign _EVAL_2629 = _EVAL_2147 < _EVAL_2435;
  assign _EVAL_413 = _EVAL_2789 & _EVAL_1371;
  assign _EVAL_2490 = _EVAL_76 == 12'hb80;
  assign _EVAL_1853 = _EVAL_2258[31:24];
  assign _EVAL_3187 = _EVAL_211 | _EVAL_1734;
  assign _EVAL_128 = _EVAL_2392;
  assign _EVAL_2114 = _EVAL_2771 ? 7'h57 : _EVAL_2162;
  assign _EVAL_2248 = _EVAL_681 | _EVAL_1104;
  assign _EVAL_258 = _EVAL_425 | _EVAL_3235;
  assign _EVAL_1448 = _EVAL_2013[22];
  assign _EVAL_1164 = _EVAL_2505 ? 8'hb : _EVAL_1955;
  assign _EVAL_1118 = _EVAL_2013[70];
  assign _EVAL_3189 = _EVAL_2397 & _EVAL_1790;
  assign _EVAL_3123 = _EVAL_1725 & _EVAL_2443;
  assign _EVAL_3163 = _EVAL_2013[82];
  assign _EVAL_1980 = _EVAL_613 ? 6'h2c : _EVAL_3101;
  assign _EVAL_116 = _EVAL_2147;
  assign _EVAL_2893 = _EVAL_959 ? 8'h4 : _EVAL_1548;
  assign _EVAL_281 = _EVAL_776[43];
  assign _EVAL_634 = {{111'd0}, _EVAL_2896};
  assign _EVAL_969 = _EVAL_2309 | _EVAL_1689;
  assign _EVAL_2655 = _EVAL_76 == 12'h340;
  assign _EVAL_1324 = _EVAL_1839 | _EVAL_1900;
  assign _EVAL_565 = _EVAL_2900 ? 8'h85 : _EVAL_2384;
  assign _EVAL_2549 = _EVAL_2920 ? _EVAL_223 : {{127'd0}, _EVAL_2828};
  assign _EVAL_2534 = _EVAL_3013 | _EVAL_2793;
  assign _EVAL_1858 = _EVAL_1272 | _EVAL_197;
  assign _EVAL_1550 = _EVAL_2258[5:1];
  assign _EVAL_1942 = _EVAL_2210 | _EVAL_421;
  assign _EVAL_884 = _EVAL_2877 | _EVAL_1553;
  assign _EVAL_171 = _EVAL_1630 | _EVAL_2148;
  assign _EVAL_415 = _EVAL_776[50];
  assign _EVAL_478 = _EVAL_895 ? 7'h7a : _EVAL_2494;
  assign _EVAL_1699 = {{111'd0}, _EVAL_2951};
  assign _EVAL_2223 = _EVAL_2161 | _EVAL_2474;
  assign _EVAL_2929 = _EVAL_889 | _EVAL_373;
  assign _EVAL_2564 = _EVAL_390 ? 7'h65 : _EVAL_1428;
  assign _EVAL_2670 = _EVAL_101 == 12'h305;
  assign _EVAL_2544 = _EVAL_3031 | _EVAL_3117;
  assign _EVAL_1137 = _EVAL_776[70];
  assign _EVAL_2707 = _EVAL_2013[117];
  assign _EVAL_3087 = _EVAL_2411 ? 5'h1c : _EVAL_860;
  assign _EVAL_456 = _EVAL_1525[0];
  assign _EVAL_120 = _EVAL_2676;
  assign _EVAL_1723 = _EVAL_1927 | _EVAL_365;
  assign _EVAL_2011 = _EVAL_2317[39:32];
  assign _EVAL_2656 = _EVAL_2233 ? 6'h2d : _EVAL_1980;
  assign _EVAL_540 = _EVAL_776[109];
  assign _EVAL_1294 = _EVAL_101 == 12'hb03;
  assign _EVAL_832 = _EVAL_776[138];
  assign _EVAL_1134 = _EVAL_2680 & _EVAL_121;
  assign _EVAL_2121 = _EVAL_1569 | _EVAL_2771;
  assign _EVAL_1756 = _EVAL_2838 ? 8'h9 : _EVAL_1937;
  assign _EVAL_2418 = _EVAL_776[125];
  assign _EVAL_885 = _EVAL_461 | _EVAL_1415;
  assign _EVAL_1088 = _EVAL_2258[23:16];
  assign _EVAL_3202 = _EVAL_76 == 12'h7c1;
  assign _EVAL_1148 = _EVAL_251[6];
  assign _EVAL_447 = _EVAL_1635 | _EVAL_2813;
  assign _EVAL_874 = _EVAL_558 | _EVAL_1208;
  assign _EVAL_1313 = _EVAL_489 ? 8'h2b : _EVAL_2160;
  assign _EVAL_2587 = _EVAL_431 | _EVAL_1616;
  assign _EVAL_2824 = _EVAL_1907 == 2'h3;
  assign _EVAL_2363 = _EVAL_3163 ? 8'h52 : _EVAL_3171;
  assign _EVAL_1004 = _EVAL_776[137];
  assign _EVAL_1191 = _EVAL_2477 | _EVAL_810;
  assign _EVAL_2720 = _EVAL_785 | _EVAL_2728;
  assign _EVAL_2981 = _EVAL_582 ? 8'h78 : _EVAL_3067;
  assign _EVAL_2125 = _EVAL_1520 | _EVAL_2546;
  assign _EVAL_1163 = _EVAL_1782 ? 8'h7a : _EVAL_2976;
  assign _EVAL_337 = _EVAL_101 == 12'hc80;
  assign _EVAL_1684 = _EVAL_76 == 12'hc93;
  assign _EVAL_58 = _EVAL_334;
  assign _EVAL_2149 = _EVAL_76 == 12'h343;
  assign _EVAL_287 = _EVAL_1459 | _EVAL_829;
  assign _EVAL_2449 = _EVAL_1009 & _EVAL_526;
  assign _EVAL_2976 = _EVAL_3149 ? 8'h79 : _EVAL_2981;
  assign _EVAL_158 = _EVAL_1429 ? 8'h14 : _EVAL_2590;
  assign _EVAL_2680 = _EVAL_101 == 12'hf14;
  assign _EVAL_1831 = _EVAL_3075 | _EVAL_2647;
  assign _EVAL_44 = _EVAL_507;
  assign _EVAL_91 = _EVAL_17;
  assign _EVAL_1460 = {{2'd0}, _EVAL_2147};
  assign _EVAL_552 = _EVAL_776[116];
  assign _EVAL_463 = _EVAL_2842 | _EVAL_514;
  assign _EVAL_170 = _EVAL_776[58];
  assign _EVAL_2278 = _EVAL_446 | _EVAL_1659;
  assign _EVAL_813 = _EVAL_776[63];
  assign _EVAL_830 = _EVAL_1792 | _EVAL_954;
  assign _EVAL_2093 = _EVAL_2849 | _EVAL_1714;
  assign _EVAL_1149 = _EVAL_1245 | _EVAL_871;
  assign _EVAL_3067 = _EVAL_986 ? 8'h77 : _EVAL_1838;
  assign _EVAL_2550 = _EVAL_3049 | 32'h1;
  assign _EVAL_146 = _EVAL_2865 | _EVAL_2323;
  assign _EVAL_2151 = 2'h2 == _EVAL_1512 ? _EVAL_612 : _EVAL_2335;
  assign _EVAL_46 = _EVAL_850;
  assign _EVAL_3215 = 2'h3 == _EVAL_1512 ? _EVAL_1450 : _EVAL_2964;
  assign _EVAL_1495 = {{16'd0}, _EVAL_1144};
  assign _EVAL_374 = 2'h3 == _EVAL_1512 ? _EVAL_315 : _EVAL_3008;
  assign _EVAL_544 = _EVAL_1554 | _EVAL_2274;
  assign _EVAL_2041 = _EVAL_1610 ? 1'h0 : _EVAL_1722;
  assign _EVAL_677 = _EVAL_556 & _EVAL_1310;
  assign _EVAL_724 = _EVAL_2457 | _EVAL_170;
  assign _EVAL_769 = _EVAL_1525[5];
  assign _EVAL_2005 = _EVAL_3097 & _EVAL_1659;
  assign _EVAL_1478 = _EVAL_777 | _EVAL_2386;
  assign _EVAL_1656 = _EVAL_1289 ? 8'h74 : _EVAL_1360;
  assign _EVAL_2996 = _EVAL_1448 ? 8'h16 : _EVAL_1760;
  assign _EVAL_1599 = _EVAL_3097 & _EVAL_2227;
  assign _EVAL_1857 = _EVAL_76 == 12'h304;
  assign _EVAL_761 = _EVAL_700 ? _EVAL_1881 : 32'h0;
  assign _EVAL_512 = _EVAL_1777 | _EVAL_336;
  assign _EVAL_2917 = _EVAL_776[83];
  assign _EVAL_2621 = _EVAL_2787[2];
  assign _EVAL_1695 = _EVAL_76 == 12'hc06;
  assign _EVAL_2225 = _EVAL_776[89];
  assign _EVAL_22 = _EVAL_1507;
  assign _EVAL_1050 = _EVAL_1853[0];
  assign _EVAL_2190 = _EVAL_767 & 32'hf;
  assign _EVAL_509 = _EVAL_1157 ? 1'h0 : _EVAL_1324;
  assign _EVAL_1729 = _EVAL_525 & _EVAL_59;
  assign _EVAL_1731 = _EVAL_1592 ? 5'h18 : _EVAL_1744;
  assign _EVAL_758 = _EVAL_49 & _EVAL_39;
  assign _EVAL_1917 = _EVAL_1525[7];
  assign _EVAL_2901 = _EVAL_1060 | _EVAL_2661;
  assign _EVAL_1131 = {_EVAL_299, 6'h0};
  assign _EVAL_513 = _EVAL_76 == 12'h3b8;
  assign _EVAL_834 = {_EVAL_3143,_EVAL_2844,_EVAL_2593,_EVAL_2355,_EVAL_1888,_EVAL_1172,_EVAL_2609};
  assign _EVAL_3048 = _EVAL_1300 | _EVAL_499;
  assign _EVAL_407 = _EVAL_76 == 12'h33f;
  assign _EVAL_872 = _EVAL_2385 | _EVAL_2741;
  assign _EVAL_564 = _EVAL_3016 ? 7'h6e : _EVAL_3064;
  assign _EVAL_938 = _EVAL_2289 ? 7'h4b : _EVAL_1299;
  assign _EVAL_2009 = _EVAL_2013[54];
  assign _EVAL_2541 = ~_EVAL_3224;
  assign _EVAL_1933 = _EVAL_2013[19];
  assign _EVAL_1036 = _EVAL_76 == 12'hb83;
  assign _EVAL_556 = ~_EVAL_2299;
  assign _EVAL_1976 = _EVAL_2013[47];
  assign _EVAL_1244 = _EVAL_1878 ? _EVAL_1097 : _EVAL_424;
  assign _EVAL_1386 = _EVAL_3076 == 32'h20000000;
  assign _EVAL_1774 = _EVAL_1390 | _EVAL_3016;
  assign _EVAL_626 = _EVAL_76 == 12'hb8a;
  assign _EVAL_118 = _EVAL_269;
  assign _EVAL_3120 = _EVAL_1618 ? 7'h48 : _EVAL_2069;
  assign _EVAL_523 = _EVAL_76 == 12'hc91;
  assign _EVAL_773 = _EVAL_2075 ? 7'h5d : _EVAL_849;
  assign _EVAL_3127 = _EVAL_76 == 12'hc82;
  assign _EVAL_1093 = _EVAL_2853 ? 8'h72 : _EVAL_956;
  assign _EVAL_1528 = _EVAL_1578 & _EVAL_2227;
  assign _EVAL_718 = _EVAL_573 | _EVAL_2900;
  assign _EVAL_41 = _EVAL_3170;
  assign _EVAL_3186 = _EVAL_1545 | _EVAL_813;
  assign _EVAL_3248 = ~_EVAL_2904;
  assign _EVAL_2863 = _EVAL_76 == 12'h32c;
  assign _EVAL_303 = {_EVAL_333,_EVAL_2003};
  assign _EVAL_2502 = _EVAL_2139 | _EVAL_3193;
  assign _EVAL_2404 = _EVAL | _EVAL_2567;
  assign _EVAL_182 = _EVAL_2013[45];
  assign _EVAL_1752 = _EVAL_76 == 12'hb87;
  assign _EVAL_1302 = _EVAL_1202 & _EVAL_3036;
  assign _EVAL_594 = _EVAL_76 == 12'hc1b;
  assign _EVAL_362 = _EVAL_2350 | _EVAL_1599;
  assign _EVAL_712 = {_EVAL_926,1'h0,1'h0,_EVAL_3215,_EVAL_1122,_EVAL_2743,_EVAL_374};
  assign _EVAL_1044 = _EVAL_1594 | _EVAL_1560;
  assign _EVAL_1133 = _EVAL_76 == 12'h338;
  assign _EVAL_1489 = _EVAL_311 | _EVAL_1462;
  assign _EVAL_1558 = _EVAL_2991 ? _EVAL_2258 : {{2'd0}, _EVAL_333};
  assign _EVAL_3125 = _EVAL_76 == 12'hc05;
  assign _EVAL_2203 = _EVAL_776[67];
  assign _EVAL_353 = _EVAL_1585 | _EVAL_552;
  assign _EVAL_3100 = _EVAL_2862[30:0];
  assign _EVAL_2779 = _EVAL_2788 | _EVAL_1537;
  assign _EVAL_293 = _EVAL_2147 > 2'h1;
  assign _EVAL_177 = _EVAL_1628 | _EVAL_1365;
  assign _EVAL_419 = _EVAL_1004 ? 8'h89 : _EVAL_607;
  assign _EVAL_1915 = _EVAL_1829 | _EVAL_159;
  assign _EVAL_1698 = _EVAL_1637 ? 6'h33 : _EVAL_2026;
  assign _EVAL_204 = 2'h2 == _EVAL_1512 ? _EVAL_2306 : _EVAL_2352;
  assign _EVAL_505 = _EVAL_2453 | _EVAL_1448;
  assign _EVAL_1626 = _EVAL_705 | _EVAL_2164;
  assign _EVAL_3025 = _EVAL_2954 & _EVAL_526;
  assign _EVAL_1060 = _EVAL_508 | _EVAL_1699;
  assign _EVAL_1289 = _EVAL_2013[116];
  assign _EVAL_2794 = ~_EVAL_1329;
  assign _EVAL_2321 = _EVAL_2704 | _EVAL_2729;
  assign _EVAL_2261 = _EVAL_776[11];
  assign _EVAL_345 = _EVAL_2673 & _EVAL_2965;
  assign _EVAL_2314 = _EVAL_1795 | _EVAL_781;
  assign _EVAL_1918 = _EVAL_2013[129];
  assign _EVAL_1616 = _EVAL_2013[142];
  assign _EVAL_1914 = _EVAL_2000 | _EVAL_1693;
  assign _EVAL_1420 = _EVAL_2125 | _EVAL_634;
  assign _EVAL_663 = {_EVAL_2251,_EVAL_2665};
  assign _EVAL_1385 = _EVAL_76 == 12'h7b2;
  assign _EVAL_2300 = _EVAL_2848 ? _EVAL_1267 : 8'h0;
  assign _EVAL_3053 = {4'h2,_EVAL_2434,14'h400,_EVAL_821,_EVAL_2231,2'h0,_EVAL_2562,_EVAL_712};
  assign _EVAL_584 = _EVAL_2013[107];
  assign _EVAL_265 = _EVAL_76 == 12'h344;
  assign _EVAL_3237 = _EVAL_1016 | _EVAL_2029;
  assign _EVAL_1436 = _EVAL_1739 & 32'h20400000;
  assign _EVAL_2521 = _EVAL_2504 | _EVAL_2135;
  assign _EVAL_80 = _EVAL_2674;
  assign _EVAL_214 = _EVAL_226 ? 4'h5 : _EVAL_1040;
  assign _EVAL_2691 = _EVAL_2410 ? 8'h81 : _EVAL_1126;
  assign _EVAL_1844 = _EVAL_76 == 12'hb10;
  assign _EVAL_2205 = _EVAL_2848 & _EVAL_1722;
  assign _EVAL_3122 = _EVAL_336 ? 8'hd : _EVAL_498;
  assign _EVAL_1452 = _EVAL_261 & _EVAL_526;
  assign _EVAL_2138 = _EVAL_76 == 12'hc94;
  assign _EVAL_1817 = _EVAL_1914 | _EVAL_626;
  assign _EVAL_2632 = _EVAL_76 == 12'hb13;
  assign _EVAL_1264 = _EVAL_1986 | _EVAL_2009;
  assign _EVAL_270 = _EVAL_2013[55];
  assign _EVAL_625 = _EVAL_2013[125];
  assign _EVAL_655 = _EVAL_2013[68];
  assign _EVAL_2862 = _EVAL_589 + 31'h1;
  assign _EVAL_283 = _EVAL_2189 | _EVAL_164;
  assign _EVAL_1012 = _EVAL_776[113];
  assign _EVAL_618 = _EVAL_1411 | _EVAL_2761;
  assign _EVAL_947 = _EVAL_76 == 12'hc83;
  assign _EVAL_2956 = _EVAL_1681 ? _EVAL_1472 : {{57'd0}, _EVAL_397};
  assign _EVAL_1930 = _EVAL_1080 | _EVAL_2845;
  assign _EVAL_805 = _EVAL_76 == 12'h3bf;
  assign _EVAL_369 = _EVAL_2489 | _EVAL_2053;
  assign _EVAL_628 = {{111'd0}, _EVAL_3160};
  assign _EVAL_1760 = _EVAL_2939 ? 8'h15 : _EVAL_158;
  assign _EVAL_3081 = _EVAL_76 == 12'hc8d;
  assign _EVAL_2802 = _EVAL_1154 | _EVAL_1919;
  assign _EVAL_1334 = _EVAL_1228 | _EVAL_2568;
  assign _EVAL_2616 = {{30'd0}, _EVAL_1692};
  assign _EVAL_1821 = ~_EVAL_1999;
  assign _EVAL_1680 = _EVAL_734 == 32'h10000000;
  assign _EVAL_1083 = _EVAL_101[10];
  assign _EVAL_2650 = _EVAL_76 == 12'hc00;
  assign _EVAL_607 = _EVAL_1818 ? 8'h88 : _EVAL_605;
  assign _EVAL_674 = _EVAL_2567 ? _EVAL_319 : _EVAL_2251;
  assign _EVAL_779 = _EVAL_76 == 12'h334;
  assign _EVAL_980 = _EVAL_2119 | _EVAL_18;
  assign _EVAL_12 = _EVAL_272;
  assign _EVAL_662 = _EVAL_1291 | _EVAL_1118;
  assign _EVAL_2157 = _EVAL_776[29];
  assign _EVAL_2775 = _EVAL_2944 ? 5'h1f : _EVAL_768;
  assign _EVAL_1398 = _EVAL_2750 | _EVAL_1549;
  assign _EVAL_1554 = _EVAL_1757 | _EVAL_2228;
  assign _EVAL_1839 = _EVAL_427 | _EVAL_2107;
  assign _EVAL_3131 = _EVAL_539 ? 8'h63 : _EVAL_2690;
  assign _EVAL_1077 = {{111'd0}, _EVAL_1495};
  assign _EVAL_367 = _EVAL_76 == 12'h3a0;
  assign _EVAL_1207 = _EVAL_776[25];
  assign _EVAL_775 = _EVAL_2580 ? 8'h8 : _EVAL_2994;
  assign _EVAL_60 = _EVAL_494;
  assign _EVAL_973 = _EVAL_2163 | _EVAL_1961;
  assign _EVAL_296 = _EVAL_1117 ? _EVAL_3079 : _EVAL_417;
  assign _EVAL_903 = _EVAL_3186 | _EVAL_2569;
  assign _EVAL_1618 = _EVAL_776[72];
  assign _EVAL_953 = _EVAL_2848 ? 1'h0 : _EVAL_113;
  assign _EVAL_3119 = {{113'd0}, _EVAL_2342};
  assign _EVAL_1956 = _EVAL_1089 & _EVAL_2378;
  assign _EVAL_2934 = _EVAL_76 == 12'hb9a;
  assign _EVAL_1900 = _EVAL_776[4];
  assign _EVAL_749 = _EVAL_1813 | _EVAL_2095;
  assign _EVAL_52 = _EVAL_3052;
  assign _EVAL_3086 = _EVAL_162 ? 7'h5a : _EVAL_2662;
  assign _EVAL_2073 = _EVAL_76 == 12'hc89;
  assign _EVAL_883 = _EVAL_776[102];
  assign _EVAL_1199 = _EVAL_3 == 2'h3;
  assign _EVAL_2766 = _EVAL_2258[31:16];
  assign _EVAL_1541 = _EVAL_2013[63];
  assign _EVAL_159 = _EVAL_1525[11];
  assign _EVAL_631 = _EVAL_2013[123];
  assign _EVAL_1593 = _EVAL_3219 ? _EVAL_2258 : {{2'd0}, _EVAL_2799};
  assign _EVAL_1371 = ~_EVAL_2899;
  assign _EVAL_1305 = _EVAL_1209 | _EVAL_1928;
  assign _EVAL_1272 = _EVAL_2333 | _EVAL_1642;
  assign _EVAL_202 = _EVAL_1191 | _EVAL_2319;
  assign _EVAL_923 = _EVAL_1389 | _EVAL_2472;
  assign _EVAL_1074 = _EVAL_1056 ? 7'h76 : _EVAL_1381;
  assign _EVAL_1987 = _EVAL_1347 | _EVAL_855;
  assign _EVAL_306 = _EVAL_76 >= 12'hc80;
  assign _EVAL_2256 = _EVAL_2013[77];
  assign _EVAL_3051 = _EVAL_1877 ? 8'h6e : _EVAL_2056;
  assign _EVAL_3096 = _EVAL_316 ? 8'h83 : _EVAL_2279;
  assign _EVAL_717 = _EVAL_2105 | _EVAL_1289;
  assign _EVAL_876 = _EVAL_1858 | _EVAL_1367;
  assign _EVAL_1909 = _EVAL_2591 | _EVAL_254;
  assign _EVAL_1330 = _EVAL_305 | _EVAL_2876;
  assign _EVAL_1757 = _EVAL_1179 | _EVAL_2261;
  assign _EVAL_351 = _EVAL_776[20];
  assign _EVAL_2400 = _EVAL_2709 | _EVAL_901;
  assign _EVAL_1128 = _EVAL_1514 | _EVAL_584;
  assign _EVAL_1209 = _EVAL_2492 | _EVAL_962;
  assign _EVAL_473 = _EVAL_811 | _EVAL_1742;
  assign _EVAL_2937 = _EVAL_1294 ? _EVAL_3043 : {{33'd0}, _EVAL_2239};
  assign _EVAL_135 = _EVAL_2914;
  assign _EVAL_23 = _EVAL_1948;
  assign _EVAL_2994 = _EVAL_2495 ? 8'h0 : _EVAL_472;
  assign _EVAL_2838 = _EVAL_2013[9];
  assign _EVAL_1877 = _EVAL_2013[110];
  assign _EVAL_1671 = 32'h80000000 + _EVAL_3042;
  assign _EVAL_3044 = _EVAL_3239 + 58'h1;
  assign _EVAL_2986 = _EVAL_2716 | _EVAL_3156;
  assign _EVAL_1362 = _EVAL_2013[74];
  assign _EVAL_2135 = _EVAL_776[92];
  assign _EVAL_57 = _EVAL_699;
  assign _EVAL_862 = _EVAL_2909 ? _EVAL_3 : 2'h0;
  assign _EVAL_2834 = _EVAL_357 ? 8'h1 : _EVAL_911;
  assign _EVAL_1627 = _EVAL_2256 ? 8'h4d : _EVAL_278;
  assign _EVAL_2857 = _EVAL_646 | _EVAL_3014;
  assign _EVAL_34 = _EVAL_3026[31:0];
  assign _EVAL_3112 = {_EVAL_2867,2'h3};
  assign _EVAL_1952 = _EVAL_1308 | _EVAL_2138;
  assign _EVAL_336 = _EVAL_2013[13];
  assign _EVAL_2809 = _EVAL_1487[0];
  assign _EVAL_3102 = _EVAL_76 == 12'hc1e;
  assign _EVAL_698 = {{25'd0}, _EVAL_961};
  assign _EVAL_1825 = _EVAL_2567 ? _EVAL_2395 : _EVAL_1948;
  assign _EVAL_2411 = _EVAL_776[28];
  assign _EVAL_534 = _EVAL_76 == 12'hb1e;
  assign _EVAL_1515 = _EVAL_550 ? _EVAL_581 : 64'h0;
  assign _EVAL_901 = _EVAL_2013[136];
  assign _EVAL_2895 = _EVAL_3254[7:0];
  assign _EVAL_1275 = _EVAL_2013[91];
  assign _EVAL_379 = _EVAL_361 | _EVAL_1618;
  assign _EVAL_2092 = _EVAL_968 ? 8'h54 : _EVAL_224;
  assign _EVAL_2590 = _EVAL_1933 ? 8'h13 : _EVAL_2059;
  assign _EVAL_1730 = _EVAL_776[112];
  assign _EVAL_3164 = _EVAL_1783 | _EVAL_2130;
  assign _EVAL_597 = _EVAL_1121 ? 8'h19 : _EVAL_684;
  assign _EVAL_1079 = {_EVAL_850,_EVAL_1310};
  assign _EVAL_2098 = _EVAL_2013[75];
  assign _EVAL_244 = _EVAL_625 ? 8'h7d : _EVAL_420;
  assign _EVAL_1846 = _EVAL_2142 & _EVAL_1396;
  assign _EVAL_2366 = _EVAL_2848 ? 1'h0 : _EVAL_40;
  assign _EVAL_2047 = _EVAL_943 | _EVAL_2678;
  assign _EVAL_2168 = _EVAL_1079 + 31'h1;
  assign _EVAL_363 = _EVAL_2013[41];
  assign _EVAL_2527 = _EVAL_2305 ? _EVAL_862 : 2'h0;
  assign _EVAL_444 = _EVAL_1961 ? 6'h34 : _EVAL_1698;
  assign _EVAL_2344 = _EVAL_3245 ? 7'h4d : _EVAL_2833;
  assign _EVAL_2325 = _EVAL_1823 ? 7'h72 : _EVAL_3035;
  assign _EVAL_1454 = _EVAL_2281 | _EVAL_2908;
  assign _EVAL_2677 = _EVAL_1969 + 34'h1;
  assign _EVAL_2983 = _EVAL_2258[30];
  assign _EVAL_1462 = _EVAL_776[104];
  assign _EVAL_2666 = _EVAL_167 | _EVAL_1546;
  assign _EVAL_907 = _EVAL_824 ? 8'h8a : _EVAL_454;
  assign _EVAL_1424 = _EVAL_2001 & _EVAL_1384;
  assign _EVAL_1808 = _EVAL_3088 ? 11'h489 : 11'h0;
  assign _EVAL_2160 = _EVAL_1849 ? 8'h2a : _EVAL_2269;
  assign _EVAL_1416 = _EVAL_2511 | _EVAL_2256;
  assign _EVAL_1763 = _EVAL_2221 | _EVAL_2657;
  assign _EVAL_2815 = _EVAL_1098 & _EVAL_1790;
  assign _EVAL_2049 = 2'h2 == _EVAL_1512 ? _EVAL_845 : _EVAL_3209;
  assign _EVAL_916 = _EVAL_2677[33:0];
  assign _EVAL_2498 = _EVAL_1659 ? 12'h800 : 12'h808;
  assign _EVAL_2191 = _EVAL_1894 | _EVAL_941;
  assign _EVAL_2869 = _EVAL_76 == 12'hb99;
  assign _EVAL_1440 = _EVAL_1573 | _EVAL_2810;
  assign _EVAL_1979 = _EVAL_1799 | _EVAL_1235;
  assign _EVAL_2026 = _EVAL_415 ? 6'h32 : _EVAL_2173;
  assign _EVAL_3069 = _EVAL_1031 | _EVAL_1177;
  assign _EVAL_1428 = _EVAL_1812 ? 7'h64 : _EVAL_2338;
  assign _EVAL_2586 = _EVAL_2123 ? 8'h8e : _EVAL_2419;
  assign _EVAL_2159 = _EVAL_581[63:32];
  assign _EVAL_1104 = _EVAL_76 == 12'hb89;
  assign _EVAL_3021 = _EVAL_584 ? 8'h6b : _EVAL_2441;
  assign _EVAL_2229 = _EVAL_2713[27];
  assign _EVAL_119 = _EVAL_3217;
  assign _EVAL_1433 = _EVAL_170 ? 6'h3a : _EVAL_913;
  assign _EVAL_1457 = _EVAL_2717 | _EVAL_655;
  assign _EVAL_2736 = _EVAL_76 == 12'hb8b;
  assign _EVAL_515 = _EVAL_776[119];
  assign _EVAL_1553 = _EVAL_76 == 12'hc17;
  assign _EVAL_2101 = _EVAL_1681 ? _EVAL_1603 : {{2'd0}, _EVAL_850};
  assign _EVAL_1157 = _EVAL_2848 & _EVAL_3180;
  assign _EVAL_129 = _EVAL_2471;
  assign _EVAL_441 = _EVAL_892 | _EVAL_291;
  assign _EVAL_2748 = _EVAL_825 | _EVAL_2584;
  assign _EVAL_1651 = _EVAL_1044 | _EVAL_2817;
  assign _EVAL_2741 = _EVAL_2013[5];
  assign _EVAL_1384 = _EVAL_1742 | _EVAL_2647;
  assign _EVAL_2649 = {{5'd0}, _EVAL};
  assign _EVAL_543 = _EVAL_776[53];
  assign _EVAL_2989 = _EVAL_1208 ? 8'h5f : _EVAL_2090;
  assign _EVAL_2972 = _EVAL_76 == 12'hb8e;
  assign _EVAL_2727 = {4'h2,_EVAL_2842,14'h400,_EVAL_2784,_EVAL_3115,2'h0,_EVAL_2445,_EVAL_3168};
  assign _EVAL_1214 = _EVAL_402 | _EVAL_1207;
  assign _EVAL_53 = _EVAL_685;
  assign _EVAL_2222 = _EVAL_2157 ? 5'h1d : _EVAL_3087;
  assign _EVAL_1842 = _EVAL_350 | _EVAL_2658;
  assign _EVAL_1562 = _EVAL_76 == 12'hb09;
  assign _EVAL_3214 = _EVAL_1951 | _EVAL_2668;
  assign _EVAL_3095 = {{5'd0}, _EVAL_61};
  assign _EVAL_2455 = {_EVAL_1318,_EVAL_2205,_EVAL_1620,_EVAL_2949,_EVAL_728,_EVAL_2300,_EVAL_429,_EVAL_2479};
  assign _EVAL_828 = _EVAL_76 == 12'h336;
  assign _EVAL_3105 = _EVAL_1453 | _EVAL_2804;
  assign _EVAL_86 = _EVAL_1279;
  assign _EVAL_394 = _EVAL_76 == 12'hc8b;
  assign _EVAL_1174 = _EVAL_2013[73];
  assign _EVAL_1069 = _EVAL_2013[105];
  assign _EVAL_588 = _EVAL_2013[29];
  assign _EVAL_936 = {_EVAL_168, 2'h0};
  assign _EVAL_2462 = _EVAL_2013[71];
  assign _EVAL_2448 = _EVAL_182 ? 8'h2d : _EVAL_2322;
  assign _EVAL_1024 = _EVAL_76 == 12'h3b2;
  assign _EVAL_960 = _EVAL_1436 == 32'h20000000;
  assign _EVAL_1400 = _EVAL_76 == 12'h333;
  assign _EVAL_2487 = _EVAL_1853[7];
  assign _EVAL_1644 = _EVAL_1794 | _EVAL_815;
  assign _EVAL_979 = _EVAL_2076 ? 8'h42 : _EVAL_1631;
  assign _EVAL_2792 = _EVAL_2615 | _EVAL_1275;
  assign _EVAL_1986 = _EVAL_2314 | _EVAL_270;
  assign _EVAL_526 = ~_EVAL_2647;
  assign _EVAL_2489 = _EVAL_1916 | _EVAL_1793;
  assign _EVAL_2105 = _EVAL_1704 | _EVAL_2707;
  assign _EVAL_2317 = {_EVAL_1969,_EVAL_3070};
  assign _EVAL_2753 = _EVAL_2813 ? 7'h45 : _EVAL_1065;
  assign _EVAL_278 = _EVAL_702 ? 8'h4c : _EVAL_2652;
  assign _EVAL_2697 = _EVAL_1853[1];
  assign _EVAL_1482 = _EVAL_279[5:1];
  assign _EVAL_169 = _EVAL_2133 | _EVAL_2647;
  assign _EVAL_2805 = _EVAL_487 | _EVAL_832;
  assign _EVAL_2880 = _EVAL_581[63:32];
  assign _EVAL_299 = _EVAL_279[31:6];
  assign _EVAL_133 = _EVAL_1587[31:0];
  assign _EVAL_172 = _EVAL_810 ? 6'h38 : _EVAL_3162;
  assign _EVAL_1000 = _EVAL_2502 | _EVAL_1766;
  assign _EVAL_2725 = _EVAL_1853[2];
  assign _EVAL_2396 = _EVAL_795 | _EVAL_2145;
  assign _EVAL_2162 = _EVAL_3060 ? 7'h56 : _EVAL_2875;
  assign _EVAL_806 = _EVAL_1519 | _EVAL_404;
  assign _EVAL_1027 = _EVAL_2013[104];
  assign _EVAL_2546 = {{111'd0}, _EVAL_761};
  assign _EVAL_1508 = ~_EVAL_87;
  assign _EVAL_1007 = {_EVAL_612,1'h0,1'h0,_EVAL_1755,_EVAL_935,_EVAL_1268,_EVAL_920};
  assign _EVAL_1270 = _EVAL_2034 | _EVAL_1212;
  assign _EVAL_1790 = ~_EVAL_21;
  assign _EVAL_1805 = _EVAL_776[131];
  assign _EVAL_3254 = _EVAL_446 ? {{28'd0}, _EVAL_1800} : _EVAL_1395;
  assign _EVAL_2308 = _EVAL_2945 | _EVAL_181;
  assign _EVAL_2260 = _EVAL_2960 ? _EVAL_1032 : 32'h0;
  assign _EVAL_2150 = {{1'd0}, _EVAL_1265};
  assign _EVAL_2016 = _EVAL_2013[135];
  assign _EVAL_1778 = _EVAL_1940[12];
  assign _EVAL_350 = _EVAL_1199 & _EVAL_2927;
  assign _EVAL_187 = 2'h1 == _EVAL_1512 ? _EVAL_3058 : _EVAL_2784;
  assign _EVAL_2319 = _EVAL_776[55];
  assign _EVAL_1383 = _EVAL_3246 | _EVAL_1377;
  assign _EVAL_3088 = _EVAL_101 == 12'hf11;
  assign _EVAL_1492 = _EVAL_1215 | _EVAL_1205;
  assign _EVAL_466 = _EVAL_798 ? 8'h43 : _EVAL_979;
  assign _EVAL_2873 = {{6'd0}, _EVAL_694};
  assign _EVAL_1458 = _EVAL_76 == 12'h335;
  assign _EVAL_2100 = _EVAL_76 == 12'hf13;
  assign _EVAL_3035 = _EVAL_1012 ? 7'h71 : _EVAL_1984;
  assign _EVAL_2085 = _EVAL_2909 | _EVAL_509;
  assign _EVAL_1628 = _EVAL_1523 | _EVAL_2620;
  assign _EVAL_2309 = _EVAL_2730 | _EVAL_628;
  assign _EVAL_571 = _EVAL_3080 + _EVAL_2966;
  assign _EVAL_644 = _EVAL_944[30:0];
  assign _EVAL_1173 = _EVAL_776[97];
  assign _EVAL_2920 = _EVAL_101 == 12'h304;
  assign _EVAL_354 = {{111'd0}, _EVAL_1124};
  assign _EVAL_1908 = ~_EVAL_698;
  assign _EVAL_3064 = _EVAL_540 ? 7'h6d : _EVAL_1485;
  assign _EVAL_3140 = _EVAL_2381 | _EVAL_2276;
  assign _EVAL_2516 = {_EVAL_2258,_EVAL_1802};
  assign _EVAL_1480 = {_EVAL_1595,1'h0,1'h0,_EVAL_1450,_EVAL_1608,_EVAL_819,_EVAL_315};
  assign _EVAL_1584 = _EVAL_3193 ? 7'h6b : _EVAL_570;
  assign _EVAL_1185 = _EVAL_1282 | _EVAL_3250;
  assign _EVAL_1415 = _EVAL_776[41];
  assign _EVAL_974 = _EVAL_2571 ? 4'hd : _EVAL_3029;
  assign _EVAL_1704 = _EVAL_2458 | _EVAL_971;
  assign _EVAL_1306 = _EVAL_2013[97];
  assign _EVAL_598 = _EVAL_2013[108];
  assign _EVAL_2351 = _EVAL_776[65];
  assign _EVAL_2264 = _EVAL_76 == 12'hc07;
  assign _EVAL_1319 = _EVAL_2732[1];
  assign _EVAL_2663 = _EVAL_76 == 12'hc18;
  assign _EVAL_1884 = _EVAL_2500 | _EVAL_934;
  assign _EVAL_62 = _EVAL_2732;
  assign _EVAL_2849 = _EVAL_1559 | _EVAL_234;
  assign _EVAL_1813 = _EVAL_2295 | _EVAL_828;
  assign _EVAL_491 = {_EVAL_754, 2'h0};
  assign _EVAL_2053 = _EVAL_2670 ? _EVAL_2605 : 32'h0;
  assign _EVAL_2528 = _EVAL_2962 | _EVAL_2551;
  assign _EVAL_1720 = _EVAL_3170[0];
  assign _EVAL_1928 = _EVAL_2013[101];
  assign _EVAL_2808 = _EVAL_2629 | _EVAL_701;
  assign _EVAL_200 = _EVAL_1440 | _EVAL_791;
  assign _EVAL_1261 = _EVAL_996 ? 5'h16 : _EVAL_786;
  assign _EVAL_189 = _EVAL_76 == 12'hb19;
  assign _EVAL_1099 = _EVAL_76 == 12'h307;
  assign _EVAL_590 = _EVAL_655 ? 8'h44 : _EVAL_466;
  assign _EVAL_2369 = _EVAL_1229[31:0];
  assign _EVAL_241 = _EVAL_717 | _EVAL_808;
  assign _EVAL_1929 = _EVAL_776[40];
  assign _EVAL_1705 = _EVAL_1673 ? 8'h3 : _EVAL_1688;
  assign _EVAL_79 = _EVAL_2306;
  assign _EVAL_2171 = _EVAL_1925 ? 7'h5b : _EVAL_3086;
  assign _EVAL_573 = _EVAL_2830 | _EVAL_1749;
  assign _EVAL_1882 = {_EVAL_3239,_EVAL_3256};
  assign _EVAL_1382 = _EVAL_648 | _EVAL_1568;
  assign _EVAL_2322 = _EVAL_1212 ? 8'h2c : _EVAL_1313;
  assign _EVAL_1947 = _EVAL_2915 | _EVAL_1356;
  assign _EVAL_1525 = {_EVAL_43, 14'h0};
  assign _EVAL_2106 = _EVAL_76 == 12'hb17;
  assign _EVAL_2574 = _EVAL_2013[4];
  assign _EVAL_1782 = _EVAL_2013[122];
  assign _EVAL_1394 = _EVAL_36 == 2'h3;
  assign _EVAL_65 = _EVAL_1142;
  assign _EVAL_1010 = _EVAL_973 | _EVAL_1637;
  assign _EVAL_2903 = _EVAL_1418 | _EVAL_2589;
  assign _EVAL_2425 = _EVAL_776[85];
  assign _EVAL_1910 = _EVAL_2787[7];
  assign _EVAL_2184 = _EVAL_76 == 12'h3a1;
  assign _EVAL_2548 = _EVAL_218 | _EVAL_2345;
  assign _EVAL_1255 = _EVAL_2501 ? _EVAL_1882 : 64'h0;
  assign _EVAL_1984 = _EVAL_1730 ? 7'h70 : _EVAL_1964;
  assign _EVAL_2754 = _EVAL_776[38];
  assign _EVAL_2900 = _EVAL_2013[133];
  assign _EVAL_1924 = _EVAL_2510 & _EVAL_599;
  assign _EVAL_138 = _EVAL_920;
  assign _EVAL_691 = _EVAL_76 == 12'hb91;
  assign _EVAL_493 = _EVAL_2013[90];
  assign _EVAL_2323 = _EVAL_776[99];
  assign _EVAL_621 = _EVAL_765 | _EVAL_2089;
  assign _EVAL_1486 = _EVAL_1207 ? 5'h19 : _EVAL_1731;
  assign _EVAL_852 = {{113'd0}, _EVAL_1506};
  assign _EVAL_3075 = ~_EVAL_1850;
  assign _EVAL_932 = _EVAL_2088 | _EVAL_2217;
  assign _EVAL_778 = _EVAL_2060 ? 7'h49 : _EVAL_3120;
  assign _EVAL_2685 = _EVAL_1214 | _EVAL_1592;
  assign _EVAL_2509 = _EVAL_1767 | _EVAL_641;
  assign _EVAL_2968 = _EVAL_1095 & _EVAL_933;
  assign _EVAL_70 = _EVAL_2629 | _EVAL_3166;
  assign _EVAL_3210 = _EVAL_3063 & _EVAL_2848;
  assign _EVAL_2933 = _EVAL_776[123];
  assign _EVAL_3139 = _EVAL_704 | _EVAL_1835;
  assign _EVAL_808 = _EVAL_2013[115];
  assign _EVAL_826 = _EVAL_2808 | _EVAL_2606;
  assign _EVAL_1953 = _EVAL_1830 ? _EVAL_1279 : 30'h0;
  assign _EVAL_1885 = _EVAL_830 | _EVAL_515;
  assign _EVAL_2430 = _EVAL_76 == 12'h3b3;
  assign _EVAL_1097 = {_EVAL_2258,_EVAL_1998};
  assign _EVAL_2591 = _EVAL_1364 | _EVAL_1171;
  assign _EVAL_1937 = _EVAL_232 ? 8'h1 : _EVAL_2488;
  assign _EVAL_937 = _EVAL_2013[112];
  assign _EVAL_2535 = _EVAL_76 == 12'hb1c;
  assign _EVAL_2837 = _EVAL_1240[0];
  assign _EVAL_1265 = _EVAL_1278 ? _EVAL_3152 : 31'h0;
  assign _EVAL_946 = _EVAL_1525[9];
  assign _EVAL_2715 = _EVAL_76[4:0];
  assign _EVAL_795 = _EVAL_1006 | _EVAL_2592;
  assign _EVAL_624 = _EVAL_2482 ? 8'h82 : _EVAL_2691;
  assign _EVAL_817 = _EVAL_2699[0];
  assign _EVAL_854 = ~_EVAL_2510;
  assign _EVAL_3147 = _EVAL_101 == 12'h3b3;
  assign _EVAL_454 = _EVAL_730 ? 8'h89 : _EVAL_2821;
  assign _EVAL_2592 = _EVAL_76 == 12'h32b;
  assign _EVAL_914 = _EVAL_2107 ? 3'h0 : 3'h4;
  assign _EVAL_2215 = _EVAL_1460 + 4'h8;
  assign _EVAL_730 = _EVAL_2013[137];
  assign _EVAL_765 = _EVAL_771 | _EVAL_952;
  assign _EVAL_385 = _EVAL_2013[51];
  assign _EVAL_703 = _EVAL_1351[31:6];
  assign _EVAL_33 = _EVAL_2278 | _EVAL_1117;
  assign _EVAL_986 = _EVAL_2013[119];
  assign _EVAL_2297 = {{111'd0}, _EVAL_369};
  assign _EVAL_2113 = _EVAL_2013[78];
  assign _EVAL_399 = _EVAL_1240[2];
  assign _EVAL_267 = _EVAL_2258[31];
  assign _EVAL_1916 = _EVAL_1454 | _EVAL_2150;
  assign _EVAL_2193 = _EVAL_101 == 12'h7b2;
  assign _EVAL_232 = _EVAL_2013[1];
  assign _EVAL_554 = _EVAL_76 == 12'h32f;
  assign _EVAL_2310 = _EVAL_2013[59];
  assign _EVAL_1090 = _EVAL_2013[62];
  assign _EVAL_2209 = _EVAL_76 == 12'hb90;
  assign _EVAL_1376 = 2'h1 == _EVAL_1512 ? _EVAL_1507 : _EVAL_3217;
  assign _EVAL_137 = _EVAL_820;
  assign _EVAL_2175 = _EVAL_776[17];
  assign _EVAL_959 = _EVAL_1525[4];
  assign _EVAL_470 = _EVAL_2786 | _EVAL_2367;
  assign _EVAL_2787 = _EVAL_2766[7:0];
  assign _EVAL_2589 = _EVAL_76 == 12'hc8e;
  assign _EVAL_1040 = _EVAL_1391 ? 4'h8 : {{1'd0}, _EVAL_914};
  assign _EVAL_2119 = _EVAL_2960 ? _EVAL_2888 : 32'h0;
  assign _EVAL_2688 = _EVAL_776[49];
  assign _EVAL_2788 = _EVAL_2774 | _EVAL_2411;
  assign _EVAL_1475 = _EVAL_101 == 12'h340;
  assign _EVAL_562 = _EVAL_249 | _EVAL_3037;
  assign _EVAL_922 = _EVAL_169 ? {{20'd0}, _EVAL_2611} : _EVAL_1435;
  assign _EVAL_224 = _EVAL_1636 ? 8'h53 : _EVAL_2363;
  assign _EVAL_2970 = _EVAL_381 ? 8'h85 : _EVAL_1848;
  assign _EVAL_2107 = _EVAL_776[0];
  assign _EVAL_829 = _EVAL_76 == 12'hc9d;
  assign _EVAL_3018 = _EVAL_776[141];
  assign _EVAL_582 = _EVAL_2013[120];
  assign _EVAL_1710 = _EVAL_481 ? 8'h1e : _EVAL_2057;
  assign _EVAL_49 = _EVAL_3123 & _EVAL_526;
  assign _EVAL_3216 = _EVAL_2326 ? 8'h28 : _EVAL_670;
  assign _EVAL_1694 = _EVAL_2261 ? 4'hb : _EVAL_448;
  assign _EVAL_617 = _EVAL_3218 | _EVAL_2430;
  assign _EVAL_2729 = _EVAL_776[81];
  assign _EVAL_3249 = _EVAL_76 == 12'hc1f;
  assign _EVAL_3166 = _EVAL_1323 & _EVAL_526;
  assign _EVAL_1739 = {_EVAL_101, 20'h0};
  assign _EVAL_132 = _EVAL_261;
  assign _EVAL_1989 = 2'h1 == _EVAL_1512 ? _EVAL_3213 : _EVAL_2579;
  assign _EVAL_681 = _EVAL_2701 | _EVAL_2218;
  assign _EVAL_1537 = _EVAL_776[27];
  assign _EVAL_412 = _EVAL_2190;
  assign _EVAL_2722 = _EVAL_3000 ? 4'h9 : _EVAL_2770;
  assign _EVAL_2076 = _EVAL_2013[66];
  assign _EVAL_477 = _EVAL_1398 | _EVAL_1315;
  assign _EVAL_1591 = {{111'd0}, _EVAL_1349};
  assign _EVAL_1988 = _EVAL_412 >> _EVAL_2715;
  assign _EVAL_155 = _EVAL_197 ? 8'h1b : _EVAL_748;
  assign _EVAL_3168 = {_EVAL_1493,1'h0,1'h0,_EVAL_3217,_EVAL_2268,_EVAL_2579,_EVAL_2674};
  assign _EVAL_344 = _EVAL_3057 | _EVAL_1917;
  assign _EVAL_2029 = _EVAL_2013[46];
  assign _EVAL_45 = _EVAL_1595;
  assign _EVAL_539 = _EVAL_2013[99];
  assign _EVAL_2008 = _EVAL_500 | _EVAL_380;
  assign _EVAL_899 = _EVAL_1781 | _EVAL_1580;
  assign _EVAL_2965 = _EVAL_2794 & _EVAL_918;
  assign _EVAL_2636 = _EVAL_414 | _EVAL_2934;
  assign _EVAL_713 = {_EVAL_2673,2'h0,_EVAL_1246,_EVAL_699,_EVAL_3242,_EVAL_729};
  assign _EVAL_1802 = _EVAL_581[31:0];
  assign _EVAL_2507 = _EVAL_1841 ? _EVAL_1494 : _EVAL_922;
  assign _EVAL_2974 = _EVAL_2857 | _EVAL_2255;
  assign _EVAL_235 = {{113'd0}, _EVAL_504};
  assign _EVAL_211 = _EVAL_1176 | _EVAL_2655;
  assign _EVAL_207 = _EVAL_758 | _EVAL_653;
  assign _EVAL_15 = _EVAL_864;
  assign _EVAL_2095 = _EVAL_76 == 12'hb16;
  assign _EVAL_2408 = ~_EVAL_2990;
  assign _EVAL_2435 = _EVAL_76[9:8];
  assign _EVAL_2712 = _EVAL_76 == 12'hc19;
  assign _EVAL_601 = _EVAL_2848 & _EVAL_1771;
  assign _EVAL_2506 = _EVAL_2321 | _EVAL_320;
  assign _EVAL_212 = _EVAL_776[33];
  assign _EVAL_327 = _EVAL_2013[64];
  assign _EVAL_1934 = _EVAL_76 == 12'hc1c;
  assign _EVAL_2950 = _EVAL_3243 | _EVAL_2425;
  assign _EVAL_504 = _EVAL_3147 ? _EVAL_333 : 30'h0;
  assign _EVAL_708 = ~_EVAL_644;
  assign _EVAL_1734 = _EVAL_76 == 12'h341;
  assign _EVAL_1577 = _EVAL_76 == 12'h3b4;
  assign _EVAL_3002 = _EVAL_201 | _EVAL_631;
  assign _EVAL_2326 = _EVAL_2013[40];
  assign _EVAL_2658 = _EVAL_1037 & _EVAL_269;
  assign _EVAL_2102 = ~_EVAL_1447;
  assign _EVAL_547 = _EVAL_1217 & _EVAL_269;
  assign _EVAL_160 = _EVAL_1863 & _EVAL_708;
  assign _EVAL_715 = _EVAL_1681 ? _EVAL_1593 : {{2'd0}, _EVAL_2799};
  assign _EVAL_3089 = {_EVAL_76, 20'h0};
  assign _EVAL_596 = _EVAL_101 == 12'hf13;
  assign _EVAL_3173 = _EVAL_964 | _EVAL_520;
  assign _EVAL_2269 = _EVAL_363 ? 8'h29 : _EVAL_3216;
  assign _EVAL_2524 = ~_EVAL_2129;
  assign _EVAL_2908 = {{21'd0}, _EVAL_1808};
  assign _EVAL_1366 = _EVAL_776[103];
  assign _EVAL_1517 = _EVAL_2974 | _EVAL_822;
  assign _EVAL_2730 = _EVAL_2297 | _EVAL_2906;
  assign _EVAL_489 = _EVAL_2013[43];
  assign _EVAL_2865 = _EVAL_537 | _EVAL_1812;
  assign _EVAL_320 = _EVAL_776[80];
  assign _EVAL_167 = _EVAL_1911 | _EVAL_2650;
  assign _EVAL_5 = _EVAL_1332[31:0];
  assign _EVAL_1961 = _EVAL_776[52];
  assign _EVAL_944 = _EVAL_1863 + 31'h1;
  assign _EVAL_2019 = _EVAL_501 | _EVAL_582;
  assign _EVAL_72 = _EVAL_151 == 2'h3;
  assign _EVAL_298 = _EVAL_259 ? 6'h36 : _EVAL_364;
  assign _EVAL_134 = _EVAL_819;
  assign _EVAL_2480 = _EVAL_2274 ? 4'h7 : _EVAL_2722;
  assign _EVAL_1727 = _EVAL_1626 | _EVAL_2535;
  assign _EVAL_2284 = _EVAL_661 ? 8'h8b : _EVAL_3197;
  assign _EVAL_1960 = _EVAL_1071 ? _EVAL_1512 : 2'h0;
  assign _EVAL_1796 = _EVAL_2147[0];
  assign _EVAL_2141 = _EVAL_76 == 12'hb03;
  assign _EVAL_1940 = _EVAL_1751 & _EVAL_387;
  assign _EVAL_2728 = _EVAL_76 == 12'hf11;
  assign _EVAL_2428 = _EVAL_2013[49];
  assign _EVAL_1559 = _EVAL_2890 | _EVAL_2846;
  assign _EVAL_136 = _EVAL_1755;
  assign _EVAL_1348 = _EVAL_2848 & _EVAL_2983;
  assign _EVAL_609 = _EVAL_2013[128];
  assign _EVAL_1895 = _EVAL_1158 | _EVAL_2064;
  assign _EVAL_2362 = _EVAL_1564 | _EVAL_2688;
  assign _EVAL_896 = {{111'd0}, _EVAL_2413};
  assign _EVAL_2606 = _EVAL_1184 & _EVAL_2541;
  assign _EVAL_2267 = _EVAL_1878 ? _EVAL_1881 : 32'h0;
  assign _EVAL_2087 = _EVAL_2013[32];
  assign _EVAL_2495 = _EVAL_2013[0];
  assign _EVAL_1323 = _EVAL_1386 & _EVAL_469;
  assign _EVAL_1095 = _EVAL_101 == 12'h3a0;
  assign _EVAL_1215 = _EVAL_2054 | _EVAL_3102;
  assign _EVAL_209 = _EVAL_1843 | _EVAL_1945;
  assign _EVAL_557 = _EVAL_872 | _EVAL_2580;
  assign _EVAL_1030 = _EVAL_2013[34];
  assign _EVAL_2505 = _EVAL_2013[11];
  assign _EVAL_437 = _EVAL_2258[15];
  assign _EVAL_2420 = _EVAL_76 == 12'hb8c;
  assign _EVAL_1569 = _EVAL_145 | _EVAL_1856;
  assign _EVAL_1356 = _EVAL_2013[24];
  assign _EVAL_2206 = _EVAL_2013[69];
  assign _EVAL_3006 = _EVAL_2260 | _EVAL_18;
  assign _EVAL_788 = _EVAL_2093 | _EVAL_2141;
  assign _EVAL_266 = {{1'd0}, _EVAL_3052};
  assign _EVAL_2484 = _EVAL_76 == 12'hc14;
  assign _EVAL_252 = _EVAL_1502 | _EVAL_1586;
  assign _EVAL_95 = {_EVAL_2647,_EVAL_2147};
  assign _EVAL_1686 = {5'h0,_EVAL_273,1'h0,2'h0,_EVAL_2366,1'h0,2'h0,_EVAL_953,1'h0,2'h0};
  assign _EVAL_2661 = {{111'd0}, _EVAL_3113};
  assign _EVAL_1132 = _EVAL_609 ? 8'h80 : _EVAL_2508;
  assign _EVAL_2345 = _EVAL_98 == 3'h7;
  assign _EVAL_2627 = _EVAL_490 ? 8'h3c : _EVAL_482;
  assign _EVAL_1144 = _EVAL_2848 ? 16'h0 : _EVAL_2828;
  assign _EVAL_2608 = _EVAL_714 ? 6'h25 : _EVAL_2188;
  assign _EVAL_1743 = _EVAL_2933 ? 7'h7b : _EVAL_478;
  assign _EVAL_427 = _EVAL_2470 | _EVAL_1391;
  assign _EVAL_1423 = _EVAL_1476 | _EVAL_917;
  assign _EVAL_1325 = _EVAL_621 | _EVAL_3150;
  assign _EVAL_1269 = _EVAL_692 | _EVAL_2294;
  assign _EVAL_2557 = _EVAL_241 | _EVAL_2853;
  assign _EVAL_3246 = _EVAL_2165 | _EVAL_173;
  assign _EVAL_2127 = _EVAL_101 == 12'hc00;
  assign _EVAL_130 = _EVAL_774;
  assign _EVAL_251 = _EVAL_3256 + _EVAL_2649;
  assign _EVAL_173 = _EVAL_76 == 12'h332;
  assign _EVAL_3042 = {{24'd0}, _EVAL_853};
  assign _EVAL_1235 = _EVAL_776[21];
  assign _EVAL_995 = _EVAL_76 == 12'hc86;
  assign _EVAL_1913 = {4'h2,_EVAL_1080,14'h400,_EVAL_608,_EVAL_845,2'h0,_EVAL_2914,_EVAL_1007};
  assign _EVAL_319 = _EVAL_169 ? _EVAL_2251 : _EVAL_859;
  assign _EVAL_82 = _EVAL_2673;
  assign _EVAL_36 = _EVAL_440;
  assign _EVAL_2602 = _EVAL_601 & _EVAL_2394;
  assign _EVAL_722 = _EVAL_306 & _EVAL_3179;
  assign _EVAL_1716 = _EVAL_776[78];
  assign _EVAL_1291 = _EVAL_1557 | _EVAL_2462;
  assign _EVAL_1252 = _EVAL_1387 & _EVAL_59;
  assign _EVAL_1736 = _EVAL_250 | _EVAL_2712;
  assign _EVAL_2954 = _EVAL_1532 == 12'h410;
  assign _EVAL_481 = _EVAL_2013[30];
  assign _EVAL_421 = _EVAL_2013[36];
  assign _EVAL_2702 = ~_EVAL_1971;
  assign _EVAL_558 = _EVAL_1474 | _EVAL_568;
  assign _EVAL_1777 = _EVAL_1884 | _EVAL_1446;
  assign _EVAL_2298 = _EVAL_1534 | _EVAL_3167;
  assign _EVAL_2379 = _EVAL_515 ? 7'h77 : _EVAL_1074;
  assign _EVAL_1329 = _EVAL_1246[1];
  assign _EVAL_1788 = _EVAL_76 == 12'h3b1;
  assign _EVAL_2442 = _EVAL_76 == 12'h327;
  assign _EVAL_745 = ~_EVAL_1080;
  assign _EVAL_611 = _EVAL_2651 | 32'h1;
  assign _EVAL_2013 = _EVAL_2452 ? _EVAL_2408 : 143'h0;
  assign _EVAL_139 = _EVAL_753;
  assign _EVAL_802 = _EVAL_1550 != 5'h1;
  assign _EVAL_2540 = _EVAL_2805 | _EVAL_1004;
  assign _EVAL_3031 = _EVAL_1763 | _EVAL_385;
  assign _EVAL_414 = _EVAL_1169 | _EVAL_1643;
  assign _EVAL_2681 = _EVAL_76 == 12'hb97;
  assign _EVAL_1851 = _EVAL_1224 | _EVAL_787;
  assign _EVAL_811 = _EVAL_1949 & _EVAL_2647;
  assign _EVAL_1892 = _EVAL_776[68];
  assign _EVAL_1278 = _EVAL_101 == 12'h301;
  assign _EVAL_164 = _EVAL_776[94];
  assign _EVAL_2563 = _EVAL_2258[31:6];
  assign _EVAL_1205 = _EVAL_76 == 12'hb9e;
  assign _EVAL_102 = _EVAL_2349;
  assign _EVAL_782 = _EVAL_194 ? 6'h3b : _EVAL_1433;
  assign _EVAL_3062 = {{79'd0}, _EVAL_1515};
  assign _EVAL_382 = _EVAL_493 ? 8'h5a : _EVAL_2296;
  assign _EVAL_1396 = ~_EVAL_192;
  assign _EVAL_2848 = _EVAL_1482 == 5'h1;
  assign _EVAL_1911 = _EVAL_1750 | _EVAL_2409;
  assign _EVAL_3084 = _EVAL_2567 ? _EVAL_879 : _EVAL_820;
  assign _EVAL_2056 = _EVAL_184 ? 8'h6d : _EVAL_887;
  assign _EVAL_1176 = _EVAL_1518 | _EVAL_1857;
  assign _EVAL_790 = _EVAL_294 | _EVAL_460;
  assign _EVAL_952 = _EVAL_76 == 12'h301;
  assign _EVAL_2204 = _EVAL_1739 & 32'h20200000;
  assign _EVAL_2772 = _EVAL_2013[111];
  assign _EVAL_3000 = _EVAL_776[9];
  assign _EVAL_2451 = _EVAL_320 ? 7'h50 : _EVAL_492;
  assign _EVAL_1299 = _EVAL_467 ? 7'h4a : _EVAL_778;
  assign _EVAL_754 = _EVAL_3254[4:0];
  assign _EVAL_2372 = _EVAL_2986 | _EVAL_2196;
  assign _EVAL_2130 = _EVAL_76 == 12'hc8f;
  assign _EVAL_198 = _EVAL_1118 ? 8'h46 : _EVAL_2023;
  assign _EVAL_1939 = _EVAL_101 == 12'hc03;
  assign _EVAL_726 = _EVAL_1127 ? _EVAL_880 : 32'h0;
  assign _EVAL_2280 = _EVAL_55 * 8'h4;
  assign _EVAL_2315 = _EVAL_1935[63:6];
  assign _EVAL_882 = {{30'd0}, _EVAL_2699};
  assign _EVAL_2054 = _EVAL_2250 | _EVAL_534;
  assign _EVAL_1397 = _EVAL_2013[35];
  assign _EVAL_286 = _EVAL_252 | _EVAL_1099;
  assign _EVAL_1379 = _EVAL_841 ? _EVAL_2011 : 8'h0;
  assign _EVAL_3057 = _EVAL_1915 | _EVAL_1673;
  assign _EVAL_2128 = _EVAL_1919 ? 8'hd : _EVAL_1283;
  assign _EVAL_2117 = _EVAL_800 & _EVAL_1110;
  assign _EVAL_2872 = _EVAL_3129 & _EVAL_387;
  assign _EVAL_578 = _EVAL_1146 ? _EVAL_780 : 32'h0;
  assign _EVAL_890 = _EVAL_2285 | _EVAL_1805;
  assign _EVAL_586 = _EVAL_2009 ? 8'h36 : _EVAL_2622;
  assign _EVAL_861 = _EVAL_76 == 12'hb9d;
  assign _EVAL_1673 = _EVAL_1525[3];
  assign _EVAL_404 = _EVAL_2013[79];
  assign _EVAL_1753 = _EVAL_2202 | _EVAL_2861;
  assign _EVAL_2878 = _EVAL_2539 | _EVAL_3125;
  assign _EVAL_748 = _EVAL_1367 ? 8'h1a : _EVAL_597;
  assign _EVAL_1964 = _EVAL_1596 ? 7'h6f : _EVAL_564;
  assign _EVAL_2699 = _EVAL_2258[1:0];
  assign _EVAL_2583 = _EVAL_1397 ? 8'h23 : _EVAL_330;
  assign _EVAL_2422 = _EVAL_891 | _EVAL_1995;
  assign _EVAL_2295 = _EVAL_3214 | _EVAL_1029;
  assign _EVAL_88 = _EVAL_495;
  assign _EVAL_2409 = _EVAL_76 == 12'h306;
  assign _EVAL_1333 = _EVAL_1137 ? 7'h46 : _EVAL_2753;
  assign _EVAL_1017 = _EVAL_3199 | _EVAL_481;
  assign _EVAL_2343 = _EVAL_1987 | _EVAL_1978;
  assign _EVAL_1967 = 143'h0;
  assign _EVAL_700 = _EVAL_101 == 12'hc82;
  assign _EVAL_1578 = _EVAL_3254[31];
  assign _EVAL_370 = _EVAL_76 == 12'h7b1;
  assign _EVAL_1016 = _EVAL_2653 | _EVAL_1976;
  assign _EVAL_1037 = _EVAL_3 == 2'h1;
  assign _EVAL_2667 = _EVAL_789 ? _EVAL_3144 : 32'h0;
  assign _EVAL_1204 = _EVAL_1666 ? 8'h25 : _EVAL_356;
  assign _EVAL_210 = _EVAL_718 | _EVAL_2219;
  assign _EVAL_1062 = _EVAL_313 & _EVAL_1404;
  assign _EVAL_2219 = _EVAL_2013[132];
  assign _EVAL_2097 = _EVAL_1952 | _EVAL_1458;
  assign _EVAL_2843 = _EVAL_2567 ? _EVAL_2031 : {{1'd0}, _EVAL_3052};
  assign _EVAL_228 = _EVAL_1815 & _EVAL_1778;
  assign _EVAL_2464 = {_EVAL_53,_EVAL_132,_EVAL_128,_EVAL_130,_EVAL_137,_EVAL_36,_EVAL_52,_EVAL_23,_EVAL_2752};
  assign _EVAL_2678 = _EVAL_776[76];
  assign _EVAL_1819 = _EVAL_711 & _EVAL_2003;
  assign _EVAL_2717 = _EVAL_662 | _EVAL_2206;
  assign _EVAL_672 = _EVAL_2581 | _EVAL_1012;
  assign _EVAL_2755 = _EVAL_380 ? 8'h7 : _EVAL_1756;
  assign _EVAL_925 = _EVAL_76 == 12'h331;
  assign _EVAL_3179 = _EVAL_76 < 12'hca0;
  assign _EVAL_777 = _EVAL_2308 | _EVAL_3157;
  assign _EVAL_1899 = _EVAL_1274 | _EVAL_2778;
  assign _EVAL_1737 = _EVAL_2182 ? _EVAL_1882 : 64'h0;
  assign _EVAL_2466 = _EVAL_551 | _EVAL_2410;
  assign _EVAL_2813 = _EVAL_776[69];
  assign _EVAL_1292 = _EVAL_2605[0];
  assign _EVAL_81 = _EVAL_446 ? {{28'd0}, _EVAL_1800} : _EVAL_1395;
  assign _EVAL_1958 = {72'h0,36'h0,18'h0,_EVAL_1686};
  assign _EVAL_1543 = _EVAL_2013[113];
  assign _EVAL_2737 = _EVAL_76 == 12'hb8d;
  assign _EVAL_1388 = _EVAL_76 == 12'hffc;
  assign _EVAL_875 = _EVAL_1240[4:3];
  assign _EVAL_3012 = _EVAL_1083 ? _EVAL_1821 : _EVAL_780;
  assign _EVAL_632 = _EVAL_776[48];
  assign _EVAL_508 = _EVAL_1993 | _EVAL_1985;
  assign _EVAL_3005 = _EVAL_76 == 12'hb0e;
  assign _EVAL_1122 = 2'h3 == _EVAL_1512 ? _EVAL_1608 : _EVAL_743;
  assign _EVAL_2588 = _EVAL_1678 | _EVAL_370;
  assign _EVAL_117 = _EVAL_1493;
  assign _EVAL_1194 = _EVAL_1270 | _EVAL_489;
  assign _EVAL_274 = _EVAL_2423 ? _EVAL_2011 : 8'h0;
  assign _EVAL_2468 = _EVAL_1128 | _EVAL_277;
  assign _EVAL_1240 = _EVAL_2258[7:0];
  assign _EVAL_1666 = _EVAL_2013[37];
  assign _EVAL_1125 = _EVAL_1335 | _EVAL_972;
  assign _EVAL_1476 = _EVAL_2248 | _EVAL_2073;
  assign _EVAL_627 = 32'h0;
  assign _EVAL_818 = _EVAL_2013[127];
  assign _EVAL_1116 = _EVAL_1420 | _EVAL_206;
  assign _EVAL_1533 = _EVAL_279[1:0];
  assign _EVAL_297 = _EVAL_2235 & _EVAL_2837;
  assign _EVAL_2224 = _EVAL_2016 ? 8'h87 : _EVAL_2525;
  assign _EVAL_2327 = _EVAL_903 | _EVAL_1189;
  assign _EVAL_7 = _EVAL_673;
  assign _EVAL_408 = _EVAL_1297 | _EVAL_547;
  assign _EVAL_3160 = _EVAL_2920 ? _EVAL_1495 : 32'h0;
  assign _EVAL_2510 = _EVAL_1563 & _EVAL_1077;
  assign _EVAL_2884 = _EVAL_76 == 12'h33d;
  assign _EVAL_1064 = _EVAL_76 == 12'h3a2;
  assign _EVAL_1031 = _EVAL_2898 | _EVAL_3018;
  assign _EVAL_2492 = _EVAL_2941 | _EVAL_423;
  assign _EVAL_1326 = {{111'd0}, _EVAL_2667};
  assign _EVAL_2694 = _EVAL_76 == 12'h330;
  assign _EVAL_559 = _EVAL_1095 & _EVAL_2561;
  assign _EVAL_2806 = _EVAL_353 | _EVAL_2496;
  assign _EVAL_1635 = _EVAL_856 | _EVAL_1137;
  assign _EVAL_2296 = _EVAL_2568 ? 8'h59 : _EVAL_542;
  assign _EVAL_3022 = _EVAL_2998 | _EVAL_407;
  assign _EVAL_1218 = _EVAL_1929 ? 6'h28 : _EVAL_3055;
  assign _EVAL_2711 = _EVAL_776[71];
  assign _EVAL_2889 = _EVAL_617 | _EVAL_1577;
  assign _EVAL_1085 = _EVAL_2087 ? 8'h20 : _EVAL_1033;
  assign _EVAL_2652 = _EVAL_2098 ? 8'h4b : _EVAL_1544;
  assign _EVAL_217 = _EVAL_1213 | _EVAL_2326;
  assign _EVAL_32 = _EVAL_2764;
  assign _EVAL_2703 = {{111'd0}, _EVAL_578};
  assign _EVAL_2255 = _EVAL_76 == 12'hb04;
  assign _EVAL_2030 = _EVAL_776[64];
  assign _EVAL_1380 = _EVAL_2204 == 32'h20000000;
  assign _EVAL_423 = _EVAL_2013[103];
  assign _EVAL_312 = _EVAL_2382 | _EVAL_3229;
  assign _EVAL_71 = _EVAL_315;
  assign _EVAL_3225 = {{111'd0}, _EVAL_3110};
  assign _EVAL_2822 = _EVAL_1011 | _EVAL_354;
  assign _EVAL_2241 = {_EVAL_160,2'h3};
  assign _EVAL_2958 = _EVAL_76 >= 12'hc00;
  assign _EVAL_961 = _EVAL_1464 ? 7'h7e : {{1'd0}, _EVAL_1403};
  assign _EVAL_1015 = _EVAL_202 | _EVAL_259;
  assign _EVAL_873 = _EVAL_3002 | _EVAL_1782;
  assign _EVAL_260 = _EVAL_2013[12];
  assign _EVAL_449 = _EVAL_2953 | _EVAL_2669;
  assign _EVAL_3097 = ~_EVAL_1578;
  assign _EVAL_3101 = _EVAL_281 ? 6'h2b : _EVAL_237;
  assign _EVAL_1563 = _EVAL_1958 & 143'h7fffffffffffffffffffffffffffffff0888;
  assign _EVAL_2913 = _EVAL_2258 & 32'h7ff01;
  assign _EVAL_2122 = _EVAL_256 ? 6'h20 : {{1'd0}, _EVAL_2775};
  assign _EVAL_909 = _EVAL_2013[80];
  assign _EVAL_2731 = _EVAL_776[128];
  assign _EVAL_1 = _EVAL_1353 ? _EVAL_3231 : _EVAL_2527;
  assign _EVAL_1213 = _EVAL_2234 | _EVAL_363;
  assign _EVAL_522 = ~_EVAL_3100;
  assign _EVAL_3153 = _EVAL_76 == 12'h346;
  assign _EVAL_2338 = _EVAL_2323 ? 7'h63 : _EVAL_1021;
  assign _EVAL_514 = ~_EVAL_3115;
  assign _EVAL_141 = _EVAL_1451;
  assign _EVAL_705 = _EVAL_1723 | _EVAL_411;
  assign _EVAL_1011 = _EVAL_2528 | _EVAL_1500;
  assign _EVAL_1364 = _EVAL_1334 | _EVAL_157;
  assign _EVAL_666 = _EVAL_1885 | _EVAL_1056;
  assign _EVAL_1344 = _EVAL_76 == 12'hc9f;
  assign _EVAL_1312 = _EVAL_2594 ? 8'h48 : _EVAL_1276;
  assign _EVAL_2733 = _EVAL_2013[23];
  assign _EVAL_2493 = _EVAL_2950 | _EVAL_1119;
  assign _EVAL_2543 = _EVAL_2014 | _EVAL_2100;
  assign _EVAL_1847 = _EVAL_2013[100];
  assign _EVAL_620 = _EVAL_337 ? _EVAL_2880 : 32'h0;
  assign _EVAL_2881 = _EVAL_776[134];
  assign _EVAL_1738 = _EVAL_2013[33];
  assign _EVAL_763 = _EVAL_2013[17];
  assign _EVAL_591 = _EVAL_776[98];
  assign _EVAL_1609 = _EVAL_2977 | _EVAL_521;
  assign _EVAL_734 = _EVAL_1739 & 32'h30000000;
  assign _EVAL_568 = _EVAL_2013[96];
  assign _EVAL_1873 = _EVAL_2013[124];
  assign _EVAL_3196 = _EVAL_76 == 12'hc90;
  assign _EVAL_659 = _EVAL_108 > _EVAL_2251;
  assign _EVAL_264 = ~_EVAL_1303;
  assign _EVAL_2960 = _EVAL_98[1];
  assign _EVAL_2444 = _EVAL_254 ? 8'h56 : _EVAL_2046;
  assign _EVAL_77 = _EVAL_1467;
  assign _EVAL_1617 = _EVAL_885 | _EVAL_1929;
  assign _EVAL_1982 = _EVAL_2134 | _EVAL_2736;
  assign _EVAL_707 = _EVAL_76 == 12'hb18;
  assign _EVAL_1815 = _EVAL_1513 & _EVAL_1526;
  assign _EVAL_950 = _EVAL_1856 ? 7'h58 : _EVAL_2114;
  assign _EVAL_2536 = _EVAL_101 == 12'h344;
  assign _EVAL_2750 = _EVAL_2362 | _EVAL_632;
  assign _EVAL_2998 = _EVAL_1492 | _EVAL_2461;
  assign _EVAL_1505 = _EVAL_2467 | _EVAL_1672;
  assign _EVAL_1970 = _EVAL_967 ? 6'h3c : _EVAL_782;
  assign _EVAL_2210 = _EVAL_2748 | _EVAL_1666;
  assign _EVAL_821 = 2'h3 == _EVAL_1512 ? _EVAL_495 : _EVAL_1223;
  assign _EVAL_1124 = _EVAL_1700 ? _EVAL_2880 : 32'h0;
  assign _EVAL_535 = _EVAL_1609 | _EVAL_227;
  assign _EVAL_2760 = _EVAL_1292 & _EVAL_1578;
  assign _EVAL_2169 = _EVAL_2346 ? 8'h8c : _EVAL_857;
  assign _EVAL_2940 = _EVAL_2822 | _EVAL_3175;
  assign _EVAL_3197 = _EVAL_832 ? 8'h8a : _EVAL_419;
  assign _EVAL_2277 = _EVAL_1305 | _EVAL_1847;
  assign _EVAL_314 = _EVAL_776[105];
  assign _EVAL_733 = _EVAL > 1'h0;
  assign _EVAL_1136 = _EVAL_2960 ? _EVAL_2727 : 32'h0;
  assign _EVAL_340 = _EVAL_397[6];
  assign _EVAL_2065 = _EVAL_2147 <= 2'h1;
  assign _EVAL_64 = _EVAL_1047;
  assign _EVAL_583 = _EVAL_2005 & _EVAL_2809;
  assign _EVAL_2000 = _EVAL_1423 | _EVAL_1660;
  assign _EVAL_1896 = _EVAL_2258[8:7];
  assign _EVAL_1281 = _EVAL_253 | _EVAL_805;
  assign _EVAL_1225 = _EVAL_1541 ? 8'h3f : _EVAL_2790;
  assign _EVAL_1391 = _EVAL_776[8];
  assign _EVAL_2002 = _EVAL_101 == 12'h343;
  assign _EVAL_2645 = _EVAL_606 ? 7'h7c : _EVAL_1743;
  assign _EVAL_2250 = _EVAL_287 | _EVAL_1944;
  assign _EVAL_2172 = _EVAL_1815 | _EVAL_3075;
  assign _EVAL_1073 = _EVAL_2115 | _EVAL_2094;
  assign _EVAL_3194 = _EVAL_851 | _EVAL_2647;
  assign _EVAL_316 = _EVAL_2013[131];
  assign _EVAL_1303 = _EVAL_2258[1];
  assign _EVAL_461 = _EVAL_2389 | _EVAL_1772;
  assign _EVAL_2427 = _EVAL_76 == 12'hb11;
  assign _EVAL_2823 = _EVAL_128 == 2'h3;
  assign _EVAL_877 = _EVAL_76 == 12'hb1f;
  assign _EVAL_789 = _EVAL_101 == 12'h7b0;
  assign _EVAL_1744 = _EVAL_977 ? 5'h17 : _EVAL_1261;
  assign _EVAL_1141 = _EVAL_2744 & _EVAL_3207;
  assign _EVAL_1273 = _EVAL_535 | _EVAL_1788;
  assign _EVAL_1226 = _EVAL_2257 | _EVAL_2737;
  assign _EVAL_1405 = _EVAL_1119 ? 7'h54 : _EVAL_2595;
  assign _EVAL_2063 = _EVAL_2013[31];
  assign _EVAL_221 = _EVAL_1201 | _EVAL_467;
  assign _EVAL_1039 = _EVAL_1758 | _EVAL_2265;
  assign _EVAL_856 = _EVAL_379 | _EVAL_2711;
  assign _EVAL_1823 = _EVAL_776[114];
  assign _EVAL_1983 = _EVAL_76 == 12'hc03;
  assign _EVAL_2719 = _EVAL_1681 ? _EVAL_1530 : {{2'd0}, _EVAL_1279};
  assign _EVAL_1203 = _EVAL_776[30];
  assign _EVAL_2311 = _EVAL_1154 ? 8'he : _EVAL_2128;
  assign _EVAL_1494 = {_EVAL_2185, 1'h0};
  assign _EVAL_2001 = 2'h1 == _EVAL_1512;
  assign _EVAL_1534 = _EVAL_2660 | _EVAL_2320;
  assign _EVAL_3121 = _EVAL_76 == 12'hb98;
  assign _EVAL_824 = _EVAL_2013[138];
  assign _EVAL_1677 = _EVAL_2481 ? 4'he : _EVAL_974;
  assign _EVAL_2139 = _EVAL_742 | _EVAL_391;
  assign _EVAL_2573 = ~_EVAL_156;
  assign _EVAL_373 = _EVAL_1610 & _EVAL_3169;
  assign _EVAL_1749 = _EVAL_2013[134];
  assign _EVAL_1243 = 10'h0;
  assign _EVAL_66 = _EVAL_331;
  assign _EVAL_2810 = _EVAL_76 == 12'hc88;
  assign _EVAL_1295 = _EVAL_1940[27];
  assign _EVAL_1759 = {_EVAL_2907,1'h0,1'h0,_EVAL_1507,_EVAL_2764,_EVAL_3213,_EVAL_753};
  assign _EVAL_2075 = _EVAL_776[93];
  assign _EVAL_1094 = _EVAL_351 ? 5'h14 : _EVAL_814;
  assign _EVAL_553 = _EVAL_3043[39:6];
  assign _EVAL_460 = _EVAL_776[96];
  assign _EVAL_719 = _EVAL_146 | _EVAL_591;
  assign _EVAL_2050 = _EVAL_2081 ? 32'h80000002 : 32'h0;
  assign _EVAL_2631 = _EVAL_3167 ? 5'h12 : _EVAL_1832;
  assign _EVAL_3014 = _EVAL_76 == 12'h324;
  assign _EVAL_50 = _EVAL_171 & _EVAL_3248;
  assign _EVAL_339 = _EVAL_1976 ? 8'h2f : _EVAL_1719;
  assign _EVAL_3090 = _EVAL_2557 | _EVAL_1543;
  assign _EVAL_176 = {_EVAL_2563, 6'h0};
  assign _EVAL_693 = _EVAL_76 == 12'hf12;
  assign _EVAL_1089 = _EVAL_2858[1];
  assign _EVAL_1081 = 2'h1 == _EVAL_1512 ? _EVAL_975 : _EVAL_2842;
  assign _EVAL_2156 = _EVAL_631 ? 8'h7b : _EVAL_1163;
  assign _EVAL_3250 = _EVAL_776[16];
  assign _EVAL_2086 = _EVAL_2872[12];
  assign _EVAL_2235 = _EVAL_1240[1];
  assign _EVAL_1545 = _EVAL_375 | _EVAL_2030;
  assign _EVAL_996 = _EVAL_776[22];
  assign _EVAL_2077 = _EVAL_2960 ? _EVAL_1913 : 32'h0;
  assign _EVAL_1435 = _EVAL_322 ? _EVAL_2517 : _EVAL_1131;
  assign _EVAL_1514 = _EVAL_1920 | _EVAL_598;
  assign _EVAL_10 = _EVAL_192;
  assign _EVAL_3251 = _EVAL_2496 ? 7'h73 : _EVAL_2325;
  assign _EVAL_1794 = _EVAL_1736 | _EVAL_2869;
  assign _EVAL_193 = _EVAL_2013[92];
  assign _EVAL_928 = _EVAL_642 | _EVAL_2571;
  assign _EVAL_2746 = _EVAL_2510 != 143'h0;
  assign _EVAL_688 = _EVAL_1408 & _EVAL_2647;
  assign _EVAL_993 = _EVAL_329 | _EVAL_968;
  assign _EVAL_1719 = _EVAL_2029 ? 8'h2e : _EVAL_2448;
  assign _EVAL_2231 = 2'h3 == _EVAL_1512 ? 1'h0 : _EVAL_2049;
  assign _EVAL_89 = _EVAL_3068;
  assign _EVAL_2376 = _EVAL_76 == 12'hb94;
  assign _EVAL_2057 = _EVAL_588 ? 8'h1d : _EVAL_1327;
  assign _EVAL_2279 = _EVAL_3229 ? 8'h82 : _EVAL_840;
  assign _EVAL_2152 = {{111'd0}, _EVAL_1600};
  assign _EVAL_492 = _EVAL_3165 ? 7'h4f : _EVAL_1181;
  assign _EVAL_1634 = _EVAL_2848 & _EVAL_1353;
  assign _EVAL_2429 = _EVAL_555 | _EVAL_3063;
  assign _EVAL_1338 = _EVAL_552 ? 7'h74 : _EVAL_3251;
  assign _EVAL_2595 = _EVAL_2917 ? 7'h53 : _EVAL_1965;
  assign _EVAL_1110 = _EVAL_745 | _EVAL_2647;
  assign _EVAL_800 = 2'h2 == _EVAL_1512;
  assign _EVAL_2817 = _EVAL_76 == 12'h326;
  assign _EVAL_519 = _EVAL_1882[63:32];
  assign _EVAL_2648 = _EVAL_2804 ? 7'h7e : _EVAL_1866;
  assign _EVAL_886 = _EVAL_2374 & _EVAL_387;
  assign _EVAL_2165 = _EVAL_2796 | _EVAL_523;
  assign _EVAL_954 = _EVAL_776[120];
  assign _EVAL_3229 = _EVAL_2013[130];
  assign _EVAL_1936 = _EVAL_1599 ? 2'h2 : 2'h1;
  assign _EVAL_892 = _EVAL_1407 | _EVAL_818;
  assign _EVAL_1878 = _EVAL_101 == 12'hb82;
  assign _EVAL_75 = _EVAL_2567;
  assign _EVAL_2804 = _EVAL_776[126];
  assign _EVAL_280 = _EVAL_76 == 12'hb88;
  assign _EVAL_1013 = _EVAL_404 ? 8'h4f : _EVAL_741;
  assign _EVAL_524 = _EVAL_2628 | _EVAL_606;
  assign _EVAL_452 = ~_EVAL_660;
  assign _EVAL_814 = _EVAL_2320 ? 5'h13 : _EVAL_2631;
  assign _EVAL_1993 = _EVAL_325 | _EVAL_572;
  assign _EVAL_1963 = _EVAL_905 | _EVAL_381;
  assign _EVAL_3181 = _EVAL_853 * 8'h4;
  assign _EVAL_111 = _EVAL_826 | _EVAL_3025;
  assign _EVAL_1735 = _EVAL_262 & _EVAL_526;
  assign _EVAL_19 = _EVAL_2689;
  assign _EVAL_366 = _EVAL_1294 ? _EVAL_2317 : 40'h0;
  assign _EVAL_1549 = _EVAL_776[47];
  assign _EVAL_2482 = _EVAL_776[130];
  assign _EVAL_2875 = _EVAL_2425 ? 7'h55 : _EVAL_1405;
  assign _EVAL_2348 = _EVAL_2354 | _EVAL_3249;
  assign _EVAL_84 = _EVAL_733 | _EVAL_75;
  assign _EVAL_335 = _EVAL_2533 | _EVAL_1890;
  assign _EVAL_2397 = _EVAL_2330 & _EVAL_1680;
  assign _EVAL_2020 = _EVAL_2129 | _EVAL_1685;
  assign _EVAL_2713 = _EVAL_980 & _EVAL_387;
  assign _EVAL_2853 = _EVAL_2013[114];
  assign _EVAL_3008 = 2'h2 == _EVAL_1512 ? _EVAL_920 : _EVAL_3172;
  assign _EVAL_2561 = ~_EVAL_1466;
  assign _EVAL_2163 = _EVAL_1015 | _EVAL_543;
  assign _EVAL_1812 = _EVAL_776[100];
  assign _EVAL_1693 = _EVAL_76 == 12'hc0a;
  assign _EVAL_1999 = _EVAL_2102 | _EVAL_2616;
  assign _EVAL_1619 = _EVAL_101 == 12'h7a1;
  assign _EVAL_397 = _EVAL_2644 + 6'h1;
  assign _EVAL_1332 = {_EVAL_1372,2'h3};
  assign _EVAL_917 = _EVAL_76 == 12'h32a;
  assign _EVAL_1818 = _EVAL_776[136];
  assign _EVAL_2868 = _EVAL_3099 | _EVAL_2574;
  assign _EVAL_706 = _EVAL_1275 ? 8'h5b : _EVAL_382;
  assign _EVAL_1683 = _EVAL_2258[9:0];
  assign _EVAL_1127 = _EVAL_101 == 12'h323;
  assign _EVAL_375 = _EVAL_143 | _EVAL_2351;
  assign _EVAL_3078 = _EVAL_275[30:0];
  assign _EVAL_2262 = _EVAL_76 < 12'hc20;
  assign _EVAL_2234 = _EVAL_1194 | _EVAL_1849;
  assign _EVAL_313 = _EVAL_688 & _EVAL_1930;
  assign _EVAL_1557 = _EVAL_1601 | _EVAL_2594;
  assign _EVAL_1006 = _EVAL_1817 | _EVAL_1682;
  assign _EVAL_2179 = _EVAL_3187 | _EVAL_2149;
  assign _EVAL_8 = _EVAL_2380;
  assign _EVAL_325 = _EVAL_1073 | _EVAL_896;
  assign _EVAL_2496 = _EVAL_776[115];
  assign _EVAL_1510 = _EVAL_934 ? 8'hf : _EVAL_1413;
  assign _EVAL_1179 = _EVAL_928 | _EVAL_1665;
  assign _EVAL_3013 = _EVAL_2318 | _EVAL_2442;
  assign _EVAL_704 = _EVAL_1269 | _EVAL_2460;
  assign _EVAL_855 = _EVAL_76 == 12'h3b6;
  assign _EVAL_3026 = _EVAL_1290 | _EVAL_235;
  assign _EVAL_2469 = _EVAL_2746 | _EVAL_43;
  assign _EVAL_2173 = _EVAL_2688 ? 6'h31 : _EVAL_3066;
  assign _EVAL_1231 = _EVAL_1193 | _EVAL_357;
  assign _EVAL_3079 = _EVAL_1083 ? _EVAL_2609 : _EVAL_820;
  assign _EVAL_2467 = _EVAL_220 | _EVAL_3007;
  assign _EVAL_1601 = _EVAL_179 | _EVAL_1174;
  assign _EVAL_1972 = _EVAL_571[31:0];
  assign _EVAL_2354 = _EVAL_3022 | _EVAL_877;
  assign _EVAL_2350 = _EVAL_2148 | _EVAL_1528;
  assign _EVAL_967 = _EVAL_776[60];
  assign _EVAL_3149 = _EVAL_2013[121];
  assign _EVAL_467 = _EVAL_776[74];
  assign _EVAL_365 = _EVAL_76 == 12'hb9b;
  assign _EVAL_1410 = _EVAL_1287 | _EVAL_736;
  assign _EVAL_2060 = _EVAL_776[73];
  assign _EVAL_841 = _EVAL_101 == 12'hb83;
  assign _EVAL_1245 = _EVAL_3139 | _EVAL_3046;
  assign _EVAL_859 = _EVAL_1258 ? _EVAL_108 : _EVAL_2251;
  assign _EVAL_1056 = _EVAL_776[118];
  assign _EVAL_2508 = _EVAL_818 ? 8'h7f : _EVAL_1401;
  assign _EVAL_386 = _EVAL_59 & _EVAL_525;
  assign _EVAL_2213 = _EVAL_1192 | _EVAL_3225;
  assign _EVAL_741 = _EVAL_2113 ? 8'h4e : _EVAL_1627;
  assign _EVAL_391 = _EVAL_776[108];
  assign _EVAL_220 = _EVAL_1165 | _EVAL_2632;
  assign _EVAL_106 = _EVAL_3254[31];
  assign _EVAL_1894 = _EVAL_2195 | _EVAL_616;
  assign _EVAL_1586 = _EVAL_76 == 12'hf14;
  assign _EVAL_787 = _EVAL_776[35];
  assign _EVAL_1830 = _EVAL_101 == 12'h3b0;
  assign _EVAL_2962 = _EVAL_1078 | _EVAL_2152;
  assign _EVAL_2942 = _EVAL_1681 ? _EVAL_2549 : {{127'd0}, _EVAL_2828};
  assign _EVAL_1860 = _EVAL_2787[4:3];
  assign _EVAL_2081 = _EVAL_101 == 12'hf12;
  assign _EVAL_1721 = {_EVAL_1240,_EVAL_2769};
  assign _EVAL_860 = _EVAL_1537 ? 5'h1b : _EVAL_1197;
  assign _EVAL_1585 = _EVAL_666 | _EVAL_486;
  assign _EVAL_1117 = _EVAL_2330 & _EVAL_960;
  assign _EVAL_2247 = _EVAL_906 | _EVAL_332;
  assign _EVAL_2111 = _EVAL_2713[11];
  assign _EVAL_2584 = _EVAL_2013[38];
  assign _EVAL_2955 = _EVAL_470 | _EVAL_1375;
  assign _EVAL_2088 = _EVAL_2391 | _EVAL_3163;
  assign _EVAL_648 = _EVAL_2277 | _EVAL_539;
  assign _EVAL_242 = _EVAL_2239[6];
  assign _EVAL_1907 = _EVAL_98[1:0];
  assign _EVAL_1920 = _EVAL_3206 | _EVAL_184;
  assign _EVAL_2597 = _EVAL_2569 ? 6'h3e : _EVAL_3201;
  assign _EVAL_2568 = _EVAL_2013[89];
  assign _EVAL_1869 = _EVAL_772[7];
  assign _EVAL_1965 = _EVAL_1469 ? 7'h52 : _EVAL_1715;
  assign _EVAL_2887 = _EVAL_2258[2];
  assign _EVAL_2195 = {{30'd0}, _EVAL_1960};
  assign _EVAL_502 = _EVAL_2247 | _EVAL_763;
  assign _EVAL_1484 = _EVAL_460 ? 7'h60 : _EVAL_3082;
  assign _EVAL_2500 = _EVAL_502 | _EVAL_1455;
  assign _EVAL_498 = _EVAL_260 ? 8'hc : _EVAL_1164;
  assign _EVAL_2867 = _EVAL_303 & _EVAL_480;
  assign _EVAL_1197 = _EVAL_2607 ? 5'h1a : _EVAL_1486;
  assign _EVAL_1803 = _EVAL_1681 ? _EVAL_2999 : _EVAL_1277;
  assign _EVAL_1455 = _EVAL_2013[16];
  assign _EVAL_442 = _EVAL_1071 ? _EVAL_2258 : {{30'd0}, _EVAL_1512};
  assign _EVAL_1248 = _EVAL_2258[29:28];
  assign _EVAL_2064 = _EVAL_76 == 12'hc9c;
  assign _EVAL_2189 = _EVAL_790 | _EVAL_2364;
  assign _EVAL_2374 = _EVAL_560 | _EVAL_18;
  assign _EVAL_1009 = _EVAL_2815 & _EVAL_2443;
  assign _EVAL_308 = _EVAL_3011 == 3'h0;
  assign _EVAL_31 = _EVAL_2252 | _EVAL_1394;
  assign _EVAL_292 = _EVAL_3152[2];
  assign _EVAL_2146 = _EVAL_2534 | _EVAL_2264;
  assign _EVAL_2347 = _EVAL_1419 | _EVAL_3196;
  assign _EVAL_1126 = _EVAL_2731 ? 8'h80 : {{1'd0}, _EVAL_2178};
  assign _EVAL_1681 = _EVAL_2548 | _EVAL_2421;
  assign _EVAL_1098 = _EVAL_2848 & _EVAL_2659;
  assign _EVAL_694 = _EVAL_596 ? 26'h2200826 : 26'h0;
  assign _EVAL_918 = _EVAL_1246[0];
  assign _EVAL_1473 = _EVAL_1069 ? 8'h69 : _EVAL_2447;
  assign _EVAL_2611 = _EVAL_2647 ? _EVAL_2498 : 12'h800;
  assign _EVAL_3171 = _EVAL_2217 ? 8'h51 : _EVAL_2624;
  assign _EVAL_1453 = _EVAL_1298 | _EVAL_263;
  assign _EVAL_2384 = _EVAL_2219 ? 8'h84 : _EVAL_3096;
  assign _EVAL_277 = _EVAL_2013[106];
  assign _EVAL_1347 = _EVAL_2889 | _EVAL_669;
  assign _EVAL_1078 = _EVAL_668 | _EVAL_2638;
  assign _EVAL_670 = _EVAL_1392 ? 8'h27 : _EVAL_3015;
  assign _EVAL_2971 = _EVAL_1116 | _EVAL_3119;
  assign _EVAL_1129 = _EVAL_76 == 12'hb05;
  assign _EVAL_721 = _EVAL_130 == 2'h3;
  assign _EVAL_2740 = ~_EVAL_611;
  assign _EVAL_190 = _EVAL_169 ? _EVAL_731 : 2'h3;
  assign _EVAL_727 = _EVAL_1422 == 32'h0;
  assign _EVAL_2164 = _EVAL_76 == 12'h33c;
  assign _EVAL_1949 = _EVAL_2872[27];
  assign _EVAL_356 = _EVAL_421 ? 8'h24 : _EVAL_2583;
  assign _EVAL_3016 = _EVAL_776[110];
  assign _EVAL_2472 = _EVAL_2013[65];
  assign _EVAL_2640 = _EVAL_1681 ? _EVAL_442 : {{30'd0}, _EVAL_1512};
  assign _EVAL_105 = _EVAL_2654;
  assign _EVAL_1864 = _EVAL_76 == 12'h7a2;
  assign _EVAL_962 = _EVAL_2013[102];
  assign _EVAL_2841 = _EVAL_2516[63:6];
  assign _EVAL_1054 = 2'h1 == _EVAL_1512 ? _EVAL_1142 : _EVAL_2445;
  assign _EVAL_143 = _EVAL_610 | _EVAL_3074;
  assign _EVAL_971 = _EVAL_2013[118];
  assign _EVAL_857 = _EVAL_499 ? 8'h8b : _EVAL_907;
  assign _EVAL_206 = {{113'd0}, _EVAL_1953};
  assign _EVAL_1944 = _EVAL_76 == 12'h33e;
  assign _EVAL_1906 = _EVAL_2317[39:32];
  assign _EVAL_732 = _EVAL_1306 ? 8'h61 : _EVAL_1112;
  assign _EVAL_1849 = _EVAL_2013[42];
  assign _EVAL_3113 = _EVAL_3063 ? _EVAL_2108 : 32'h0;
  assign _EVAL_1714 = _EVAL_76 == 12'h323;
  assign _EVAL_472 = _EVAL_2574 ? 8'h4 : _EVAL_2586;
  assign _EVAL_1123 = _EVAL_2521 | _EVAL_1925;
  assign _EVAL_610 = _EVAL_1488 | _EVAL_2203;
  assign _EVAL_2070 = _EVAL_76 == 12'h337;
  assign _EVAL_1274 = _EVAL_3 > _EVAL_2147;
  assign _EVAL_2324 = _EVAL_1982 | _EVAL_394;
  assign _EVAL_381 = _EVAL_776[133];
  assign _EVAL_968 = _EVAL_2013[84];
  assign _EVAL_2990 = _EVAL_854 | _EVAL_599;
  assign _EVAL_2413 = _EVAL_368 ? _EVAL_2455 : 32'h0;
  assign _EVAL_317 = _EVAL_1185 | _EVAL_690;
  assign _EVAL_1837 = _EVAL_76 == 12'h342;
  assign _EVAL_1349 = _EVAL_1807 ? _EVAL_1821 : 32'h0;
  assign _EVAL_1159 = _EVAL_1240[7];
  assign _EVAL_1792 = _EVAL_2637 | _EVAL_2271;
  assign _EVAL_194 = _EVAL_776[59];
  assign _EVAL_613 = _EVAL_776[44];
  assign _EVAL_1807 = _EVAL_101 == 12'h7b1;
  assign _EVAL_853 = _EVAL_2305 ? _EVAL_897 : _EVAL_2311;
  assign _EVAL_683 = _EVAL_2707 ? 8'h75 : _EVAL_1656;
  assign _EVAL_934 = _EVAL_2013[15];
  assign _EVAL_263 = _EVAL_776[127];
  assign _EVAL_1114 = _EVAL_101 == 12'h306;
  assign _EVAL_1614 = _EVAL_76 == 12'hb86;
  assign _EVAL_1115 = _EVAL_422 ? 8'h39 : _EVAL_2286;
  assign _EVAL_650 = _EVAL_1200 | _EVAL_2754;
  assign _EVAL_1725 = _EVAL_2216 & _EVAL_1790;
  assign _EVAL_2671 = {_EVAL_891,2'h0,_EVAL_3170,_EVAL_406,_EVAL_507,_EVAL_2349};
  assign _EVAL_2286 = _EVAL_781 ? 8'h38 : _EVAL_737;
  assign _EVAL_913 = _EVAL_2236 ? 6'h39 : _EVAL_172;
  assign _EVAL_199 = _EVAL_962 ? 8'h66 : _EVAL_1724;
  assign _EVAL_405 = _EVAL_76 == 12'hc16;
  assign _EVAL_661 = _EVAL_776[139];
  assign _EVAL_2227 = _EVAL_2895 == 8'he;
  assign _EVAL_2090 = _EVAL_2096 ? 8'h5e : _EVAL_409;
  assign _EVAL_390 = _EVAL_776[101];
  assign _EVAL_3049 = ~_EVAL_51;
  assign _EVAL_1529 = _EVAL_776[39];
  assign _EVAL_1152 = _EVAL_456 ? 8'h0 : _EVAL_2893;
  assign _EVAL_2657 = _EVAL_2013[52];
  assign _EVAL_2096 = _EVAL_2013[94];
  assign _EVAL_1119 = _EVAL_776[84];
  assign _EVAL_1375 = _EVAL_76 == 12'hb0d;
  assign _EVAL_2447 = _EVAL_1027 ? 8'h68 : _EVAL_1087;
  assign _EVAL_2690 = _EVAL_1568 ? 8'h62 : _EVAL_732;
  assign _EVAL_1331 = _EVAL_2170 & _EVAL_463;
  assign _EVAL_85 = _EVAL_1117 ? _EVAL_3012 : _EVAL_2507;
  assign _EVAL_2182 = _EVAL_101 == 12'hc02;
  assign _EVAL_73 = _EVAL_3112[31:0];
  assign _EVAL_2964 = 2'h2 == _EVAL_1512 ? _EVAL_1755 : _EVAL_1376;
  assign _EVAL_2263 = _EVAL_2062 | _EVAL_212;
  assign _EVAL_2562 = 2'h3 == _EVAL_1512 ? _EVAL_1451 : _EVAL_3116;
  assign _EVAL_2342 = _EVAL_2789 ? _EVAL_850 : 30'h0;
  assign _EVAL_2836 = {{103'd0}, _EVAL_366};
  assign _EVAL_1105 = _EVAL_2118 | _EVAL_2772;
  assign _EVAL_2394 = ~_EVAL_42;
  assign _EVAL_3106 = _EVAL_76 == 12'h7a0;
  assign _EVAL_341 = _EVAL_2111 & _EVAL_2582;
  assign _EVAL_83 = _EVAL_581[31:0];
  assign _EVAL_943 = _EVAL_2199 | _EVAL_3245;
  assign _EVAL_2902 = _EVAL_1805 ? 8'h83 : _EVAL_624;
  assign _EVAL_1886 = _EVAL_1108 | _EVAL_1738;
  assign _EVAL_616 = _EVAL_1619 ? _EVAL_3053 : 32'h0;
  assign _EVAL_436 = _EVAL_776[1];
  assign _EVAL_122 = _EVAL_3058;
  assign _EVAL_1523 = _EVAL_749 | _EVAL_405;
  assign _EVAL_302 = _EVAL_76 == 12'hb1a;
  assign _EVAL_1945 = _EVAL_76 == 12'h345;
  assign _EVAL_1893 = _EVAL_1330 | _EVAL_2484;
  assign _EVAL_2069 = _EVAL_2711 ? 7'h47 : _EVAL_1333;
  assign _EVAL_69 = _EVAL_1019;
  assign _EVAL_2660 = _EVAL_1979 | _EVAL_351;
  assign _EVAL_1905 = 2'h3 == _EVAL_1512 ? _EVAL_1239 : _EVAL_204;
  assign _EVAL_2669 = _EVAL_76 == 12'hb0f;
  assign _EVAL_906 = _EVAL_2360 | _EVAL_1933;
  assign _EVAL_2265 = _EVAL_76 == 12'hc97;
  assign _EVAL_1700 = _EVAL_101 == 12'hb80;
  assign _EVAL_871 = _EVAL_76 == 12'h3bd;
  assign _EVAL_843 = _EVAL_2685 | _EVAL_977;
  assign _EVAL_124 = _EVAL_2380 | _EVAL_103;
  assign _EVAL_546 = _EVAL_3164 | _EVAL_2694;
  assign _EVAL_445 = _EVAL_76 == 12'hb8f;
  assign _EVAL_731 = _EVAL_526 ? 2'h3 : _EVAL_2147;
  assign _EVAL_2463 = _EVAL_1226 | _EVAL_3081;
  assign _EVAL_253 = _EVAL_1149 | _EVAL_2485;
  assign _EVAL_2378 = _EVAL_2858[0];
  assign _EVAL_1689 = {{111'd0}, _EVAL_304};
  assign _EVAL_1931 = _EVAL_471 | _EVAL_2184;
  assign _EVAL_1501 = _EVAL_1738 ? 8'h21 : _EVAL_1085;
  assign _EVAL_2637 = _EVAL_740 | _EVAL_895;
  assign _EVAL_29 = _EVAL_2241[31:0];
  assign _EVAL_388 = {_EVAL_2129,2'h0,_EVAL_2732,_EVAL_3183,_EVAL_1491,_EVAL_1467,_EVAL_713,_EVAL_1399};
  assign _EVAL_2037 = _EVAL_1681 ? _EVAL_215 : {{33'd0}, _EVAL_2239};
  assign _EVAL_1856 = _EVAL_776[88];
  assign _EVAL_1389 = _EVAL_183 | _EVAL_2076;
  assign _EVAL_1859 = _EVAL_2191 | _EVAL_2873;
  assign _EVAL_2023 = _EVAL_2206 ? 8'h45 : _EVAL_590;
  assign _EVAL_2423 = _EVAL_101 == 12'hc83;
  assign _EVAL_1766 = _EVAL_776[106];
  assign _EVAL_3133 = _EVAL_835 | _EVAL_2406;
  assign _EVAL_2747 = _EVAL_243[0];
  assign _EVAL_2538 = _EVAL_3 == _EVAL_2147;
  assign _EVAL_1589 = _EVAL_3114 | _EVAL_284;
  assign _EVAL_2186 = 2'h1 == _EVAL_1512 ? _EVAL_2764 : _EVAL_2268;
  assign _EVAL_2582 = ~_EVAL_1697;
  assign _EVAL_3134 = _EVAL_1830 & _EVAL_1247;
  assign _EVAL_1150 = _EVAL_1095 & _EVAL_675;
  assign _EVAL_2211 = {_EVAL_38,_EVAL_104,_EVAL_96,_EVAL_15,_EVAL_120,_EVAL_112,_EVAL_11,_EVAL_105};
  assign _EVAL_692 = _EVAL_2343 | _EVAL_513;
  assign _EVAL_1238 = {4'h2,_EVAL_1850,14'h400,_EVAL_495,1'h0,2'h0,_EVAL_1451,_EVAL_1480};
  assign _EVAL_2458 = _EVAL_2019 | _EVAL_986;
  assign _EVAL_304 = _EVAL_1475 ? _EVAL_1271 : 32'h0;
  assign _EVAL_2569 = _EVAL_776[62];
  assign _EVAL_250 = _EVAL_2372 | _EVAL_189;
  assign _EVAL_197 = _EVAL_2013[27];
  assign _EVAL_904 = _EVAL_159 ? 8'hb : _EVAL_1705;
  assign _EVAL_1631 = _EVAL_2472 ? 8'h41 : _EVAL_1337;
  assign _EVAL_2504 = _EVAL_283 | _EVAL_2075;
  assign _EVAL_2034 = _EVAL_3237 | _EVAL_182;
  assign _EVAL_3109 = _EVAL_811 & _EVAL_2086;
  assign _EVAL_499 = _EVAL_2013[139];
  assign _EVAL_1390 = _EVAL_3059 | _EVAL_1596;
  assign _EVAL_1568 = _EVAL_2013[98];
  assign _EVAL_439 = _EVAL_2258[12];
  assign _EVAL_866 = _EVAL_76 == 12'hb1d;
  assign _EVAL_551 = _EVAL_890 | _EVAL_2482;
  assign _EVAL_3080 = {_EVAL_703, 6'h0};
  assign _EVAL_285 = _EVAL_2013[141];
  assign _EVAL_887 = _EVAL_598 ? 8'h6c : _EVAL_3021;
  assign _EVAL_1321 = _EVAL_776[132];
  assign _EVAL_671 = _EVAL_76 == 12'hc0b;
  assign _EVAL_2059 = _EVAL_332 ? 8'h12 : _EVAL_657;
  assign _EVAL_1392 = _EVAL_2013[39];
  assign _EVAL_1029 = _EVAL_76 == 12'hc95;
  assign _EVAL_1033 = _EVAL_2063 ? 8'h1f : _EVAL_1710;
  assign _EVAL_2695 = _EVAL_3033 & _EVAL_3194;
  assign _EVAL_184 = _EVAL_2013[109];
  assign _EVAL_2330 = _EVAL_98 == 3'h4;
  assign _EVAL_669 = _EVAL_76 == 12'h3b5;
  assign _EVAL_1258 = _EVAL_2449 & _EVAL_3207;
  assign _EVAL_2539 = _EVAL_1410 | _EVAL_1129;
  assign _EVAL_1985 = {{111'd0}, _EVAL_739};
  assign _EVAL_2287 = _EVAL_976 | _EVAL_2290;
  assign _EVAL_2770 = _EVAL_436 ? 4'h1 : _EVAL_214;
  assign _EVAL_1610 = _EVAL_2617 == 6'h2;
  assign _EVAL_469 = _EVAL_76[10];
  assign _EVAL_368 = _EVAL_101 == 12'h342;
  assign _EVAL_2453 = _EVAL_1947 | _EVAL_2733;
  assign _EVAL_361 = _EVAL_221 | _EVAL_2060;
  assign _EVAL_1146 = _EVAL_101 == 12'h341;
  assign _EVAL_1377 = _EVAL_76 == 12'hb12;
  assign _EVAL_1832 = _EVAL_2175 ? 5'h11 : _EVAL_667;
  assign _EVAL_933 = ~_EVAL_2673;
  assign _EVAL_2605 = _EVAL_279 & _EVAL_1908;
  assign _EVAL_1603 = _EVAL_413 ? _EVAL_2258 : {{2'd0}, _EVAL_850};
  assign _EVAL_1297 = _EVAL_2147 < 2'h1;
  assign _EVAL_1971 = _EVAL_2168[30:0];
  assign _EVAL_2786 = _EVAL_809 | _EVAL_208;
  assign _EVAL_2391 = _EVAL_993 | _EVAL_1636;
  assign _EVAL_30 = _EVAL_1353 ? _EVAL_3184 : _EVAL_1972;
  assign _EVAL_3015 = _EVAL_2584 ? 8'h26 : _EVAL_1204;
  assign _EVAL_1592 = _EVAL_776[24];
  assign _EVAL_1247 = ~_EVAL_2422;
  assign _EVAL_2819 = _EVAL_2537 | _EVAL_1695;
  assign _EVAL_218 = _EVAL_98 == 3'h6;
  assign _EVAL_1581 = _EVAL_1988[0];
  assign _EVAL_1169 = _EVAL_1241 | _EVAL_302;
  assign _EVAL_1762 = _EVAL_76 == 12'hb9f;
  assign _EVAL_1539 = _EVAL_76 == 12'hb85;
  assign _EVAL_131 = 1'h0;
  assign _EVAL_1675 = _EVAL_618 | _EVAL_490;
  assign _EVAL_311 = _EVAL_1000 | _EVAL_314;
  assign _EVAL_2761 = _EVAL_2013[61];
  assign _EVAL_2624 = _EVAL_909 ? 8'h50 : _EVAL_1013;
  assign _EVAL_532 = _EVAL_2713[12];
  assign _EVAL_879 = _EVAL_169 ? _EVAL_820 : _EVAL_1887;
  assign _EVAL_668 = _EVAL_1753 | _EVAL_948;
  assign _EVAL_3027 = _EVAL_772[3];
  assign _EVAL_2364 = _EVAL_776[95];
  assign _EVAL_1487 = _EVAL_1868 >> _EVAL_2147;
  assign _EVAL_1566 = _EVAL_1175 | _EVAL_2663;
  assign _EVAL_490 = _EVAL_2013[60];
  assign _EVAL_1588 = _EVAL_1416 | _EVAL_702;
  assign _EVAL_3228 = _EVAL_2258[27];
  assign _EVAL_1560 = _EVAL_76 == 12'hc85;
  assign _EVAL_37 = _EVAL_1671[31:0];
  assign _EVAL_710 = _EVAL_2985 | _EVAL_436;
  assign _EVAL_2604 = _EVAL_76 == 12'hc11;
  assign _EVAL_1770 = _EVAL_2192 & _EVAL_2172;
  assign _EVAL_2999 = _EVAL_3210 ? _EVAL_2545 : _EVAL_2405;
  assign _EVAL_480 = ~_EVAL_3078;
  assign _EVAL_2859 = _EVAL_2754 ? 6'h26 : _EVAL_2608;
  assign _EVAL_2692 = _EVAL_1604 ? 6'h22 : _EVAL_2440;
  assign _EVAL_770 = {{21'd0}, _EVAL_2280};
  assign _EVAL_2818 = _EVAL_1489 | _EVAL_1366;
  assign _EVAL_1192 = _EVAL_2613 | _EVAL_1591;
  assign _EVAL_1217 = _EVAL_2147 == 2'h1;
  assign _EVAL_1315 = _EVAL_776[46];
  assign _EVAL_322 = ~_EVAL_2848;
  assign _EVAL_780 = ~_EVAL_1045;
  assign _EVAL_1018 = _EVAL_2351 ? 7'h41 : _EVAL_919;
  assign _EVAL_2155 = _EVAL_954 ? 7'h78 : _EVAL_2379;
  assign _EVAL_275 = _EVAL_303 + 31'h1;
  assign _EVAL_2701 = _EVAL_200 | _EVAL_1562;
  assign _EVAL_3182 = _EVAL_1761 | _EVAL_2604;
  assign _EVAL_1308 = _EVAL_1893 | _EVAL_2376;
  assign _EVAL_2620 = _EVAL_76 == 12'hb96;
  assign _EVAL_506 = _EVAL_1123 | _EVAL_162;
  assign _EVAL_411 = _EVAL_76 == 12'hc9b;
  assign _EVAL_2494 = _EVAL_2271 ? 7'h79 : _EVAL_2155;
  assign _EVAL_284 = _EVAL_76 == 12'hc0e;
  assign _EVAL_1343 = _EVAL_937 ? 8'h70 : _EVAL_1571;
  assign _EVAL_1051 = _EVAL_1853[4:3];
  assign _EVAL_1087 = _EVAL_423 ? 8'h67 : _EVAL_199;
  assign _EVAL_1407 = _EVAL_2827 | _EVAL_609;
  assign _EVAL_2858 = _EVAL_1465[7:0];
  assign _EVAL_142 = 2'h3 == _EVAL_1512;
  assign _EVAL_2558 = _EVAL_76 == 12'h33b;
  assign _EVAL_2778 = _EVAL_1740 & _EVAL_659;
  assign _EVAL_332 = _EVAL_2013[18];
  assign _EVAL_1419 = _EVAL_2851 | _EVAL_2209;
  assign _EVAL_326 = _EVAL_1505 | _EVAL_1684;
  assign _EVAL_1290 = _EVAL_2971 | _EVAL_852;
  assign _EVAL_2446 = _EVAL_972 ? 8'h3a : _EVAL_1115;
  assign _EVAL_791 = _EVAL_76 == 12'h329;
  assign _EVAL_3207 = ~_EVAL_43;
  assign _EVAL_2395 = _EVAL_169 ? _EVAL_1948 : _EVAL_2927;
  assign _EVAL_642 = _EVAL_317 | _EVAL_2481;
  assign _EVAL_2551 = {{79'd0}, _EVAL_3020};
  assign _EVAL_3150 = _EVAL_76 == 12'h305;
  assign _EVAL_1995 = _EVAL_1466 & _EVAL_677;
  assign _EVAL_99 = _EVAL_612;
  assign _EVAL_1228 = _EVAL_2792 | _EVAL_493;
  assign _EVAL_1414 = _EVAL_1533 == 2'h0;
  assign _EVAL_2906 = _EVAL_2536 ? _EVAL_1563 : 143'h0;
  assign _EVAL_2067 = _EVAL_2881 ? 8'h86 : _EVAL_2970;
  assign _EVAL_1502 = _EVAL_1871 | _EVAL_1837;
  assign _EVAL_1506 = _EVAL_1717 ? _EVAL_2799 : 30'h0;
  assign _EVAL_2537 = _EVAL_1651 | _EVAL_2407;
  assign _EVAL_3218 = _EVAL_1273 | _EVAL_1024;
  assign _EVAL_1692 = _EVAL_292 ? 2'h1 : 2'h3;
  assign _EVAL_2533 = _EVAL_874 | _EVAL_2096;
  assign _EVAL_431 = _EVAL_2042 | _EVAL_959;
  assign _EVAL_1767 = _EVAL_2540 | _EVAL_1818;
  assign _EVAL_1233 = _EVAL_76 == 12'h7b0;
  assign _EVAL_3199 = _EVAL_759 | _EVAL_2063;
  assign _EVAL_127 = _EVAL_1246;
  assign _EVAL_2367 = _EVAL_76 == 12'h32d;
  assign _EVAL_1811 = _EVAL_76 == 12'hb92;
  assign _EVAL_3175 = {{111'd0}, _EVAL_2267};
  assign _EVAL_3055 = _EVAL_1529 ? 6'h27 : _EVAL_2859;
  assign _EVAL_2946 = _EVAL_2831 ? 8'h30 : _EVAL_339;
  assign _EVAL_1499 = _EVAL_76 == 12'hc0c;
  assign _EVAL_1658 = _EVAL_142 & _EVAL_1831;
  assign _EVAL_1171 = _EVAL_2013[87];
  assign _EVAL_3243 = _EVAL_2121 | _EVAL_3060;
  assign _EVAL_201 = _EVAL_428 | _EVAL_1873;
  assign _EVAL_2771 = _EVAL_776[87];
  assign _EVAL_3209 = 2'h1 == _EVAL_1512 ? _EVAL_192 : _EVAL_3115;
  assign _EVAL_701 = ~_EVAL_1281;
  assign _EVAL_1465 = _EVAL_2258[31:8];
  assign _EVAL_1642 = _EVAL_2013[28];
  assign _EVAL_453 = _EVAL_787 ? 6'h23 : _EVAL_2692;
  assign _EVAL_468 = _EVAL_1727 | _EVAL_1934;
  assign _EVAL_3206 = _EVAL_1105 | _EVAL_1877;
  assign _EVAL_96 = _EVAL_31;
  assign _EVAL_482 = _EVAL_2310 ? 8'h3b : _EVAL_2446;
  assign _EVAL_1485 = _EVAL_391 ? 7'h6c : _EVAL_1584;
  assign _EVAL_501 = _EVAL_873 | _EVAL_3149;
  assign _EVAL_2774 = _EVAL_435 | _EVAL_2157;
  assign _EVAL_809 = _EVAL_3198 | _EVAL_2420;
  assign _EVAL_2142 = _EVAL_2872[11];
  assign _EVAL_422 = _EVAL_2013[57];
  assign _EVAL_424 = _EVAL_2501 ? _EVAL_1187 : {{57'd0}, _EVAL_251};
  assign _EVAL_3158 = _EVAL_76 == 12'hc0f;
  assign _EVAL_825 = _EVAL_217 | _EVAL_1392;
  assign _EVAL_2517 = _EVAL_1479 ? _EVAL_3233 : _EVAL_936;
  assign _EVAL_521 = _EVAL_76 == 12'h3a3;
  assign _EVAL_576 = _EVAL_1939 ? _EVAL_2317 : 40'h0;
  assign _EVAL_1259 = _EVAL_2146 | _EVAL_1752;
  assign _EVAL_3020 = _EVAL_2127 ? _EVAL_581 : 64'h0;
  assign _EVAL_2915 = _EVAL_876 | _EVAL_1121;
  assign _EVAL_649 = _EVAL_385 ? 8'h33 : _EVAL_2529;
  assign _EVAL_1761 = _EVAL_483 | _EVAL_2427;
  assign _EVAL_1439 = _EVAL_76 == 12'hc12;
  assign _EVAL_2281 = _EVAL_1859 | _EVAL_2050;
  assign _EVAL_20 = _EVAL_2907;
  assign _EVAL_2421 = _EVAL_98 == 3'h5;
  assign _EVAL_259 = _EVAL_776[54];
  assign _EVAL_2346 = _EVAL_2013[140];
  assign _EVAL_3034 = _EVAL_2468 | _EVAL_1069;
  assign _EVAL_2389 = _EVAL_1113 | _EVAL_281;
  assign _EVAL_3046 = _EVAL_76 == 12'h3bc;
  assign _EVAL_2196 = _EVAL_76 == 12'h339;
  assign _EVAL_1399 = {_EVAL_1466,2'h0,_EVAL_3068,_EVAL_331,_EVAL_494,_EVAL_673,_EVAL_2671};
  assign _EVAL_100 = _EVAL_2579;
  assign _EVAL_3233 = {_EVAL_865,_EVAL_491};
  assign _EVAL_13 = _EVAL_1608;
  assign _EVAL_520 = _EVAL_76 == 12'hb1b;
  assign _EVAL_1551 = _EVAL_2213 | _EVAL_3062;
  assign _EVAL_739 = _EVAL_3148 ? _EVAL_3080 : 32'h0;
  assign _EVAL_223 = _EVAL_322 ? _EVAL_751 : {{127'd0}, _EVAL_2828};
  assign _EVAL_1359 = _EVAL_1174 ? 8'h49 : _EVAL_1312;
  assign _EVAL_2293 = ~_EVAL_39;
  assign _EVAL_2461 = _EVAL_76 == 12'hc9e;
  assign _EVAL_2918 = _EVAL_3044[57:0];
  assign _EVAL_110 = _EVAL_1491;
  assign _EVAL_2192 = _EVAL_1621 & _EVAL_1396;
  assign _EVAL_759 = _EVAL_1886 | _EVAL_2087;
  assign _EVAL_657 = _EVAL_763 ? 8'h11 : _EVAL_1035;
  assign _EVAL_234 = _EVAL_76 == 12'hb02;
  assign _EVAL_1685 = _EVAL_2129 & _EVAL_1819;
  assign _EVAL_2821 = _EVAL_901 ? 8'h88 : _EVAL_2224;
  assign _EVAL_290 = _EVAL_2002 ? _EVAL_2931 : 32'h0;
  assign _EVAL_2909 = _EVAL_2454 & _EVAL_1899;
  assign _EVAL_815 = _EVAL_76 == 12'hc99;
  assign _EVAL_2851 = _EVAL_870 | _EVAL_902;
  assign _EVAL_3169 = _EVAL_2305 & _EVAL_2302;
  assign _EVAL_1871 = _EVAL_2179 | _EVAL_3202;
  assign _EVAL_2571 = _EVAL_776[13];
  assign _EVAL_2216 = _EVAL_1141 | _EVAL_1634;
  assign _EVAL_919 = _EVAL_2030 ? 7'h40 : {{1'd0}, _EVAL_2803};
  assign _EVAL_487 = _EVAL_3069 | _EVAL_661;
  assign _EVAL_2236 = _EVAL_776[57];
  assign _EVAL_2460 = _EVAL_76 == 12'h3ba;
  assign _EVAL_3172 = 2'h1 == _EVAL_1512 ? _EVAL_753 : _EVAL_2674;
  assign _EVAL_1841 = _EVAL_1252 & _EVAL_1508;
  assign _EVAL_1679 = _EVAL_804 | _EVAL_2944;
  assign _EVAL_1193 = _EVAL_344 | _EVAL_946;
  assign _EVAL_645 = _EVAL_883 ? 7'h66 : _EVAL_2564;
  assign _EVAL_145 = _EVAL_506 | _EVAL_2225;
  assign _EVAL_3224 = _EVAL_293 | _EVAL_1581;
  assign _EVAL_2252 = _EVAL_721 | _EVAL_2823;
  assign _EVAL_2457 = _EVAL_474 | _EVAL_194;
  assign _EVAL_640 = _EVAL_2928 | _EVAL_2505;
  assign _EVAL_865 = _EVAL_2605[31:7];
  assign _EVAL_1594 = _EVAL_2878 | _EVAL_1539;
  assign _EVAL_3193 = _EVAL_776[107];
  assign _EVAL_2607 = _EVAL_776[26];
  assign _EVAL_2951 = _EVAL_1898 ? _EVAL_663 : 32'h0;
  assign _EVAL_2831 = _EVAL_2013[48];
  assign _EVAL_3066 = _EVAL_632 ? 6'h30 : _EVAL_1746;
  assign _EVAL_2386 = _EVAL_76 == 12'hc08;
  assign _EVAL_1165 = _EVAL_2287 | _EVAL_1400;
  assign _EVAL_3144 = {_EVAL_908,_EVAL_2987,_EVAL_619,_EVAL_2387,_EVAL_153,_EVAL_2158,_EVAL_2356,_EVAL_834};
  assign _EVAL_2613 = _EVAL_2901 | _EVAL_1326;
  assign _EVAL_2320 = _EVAL_776[19];
  assign _EVAL_2431 = _EVAL_449 | _EVAL_3158;
  assign _EVAL_2966 = {{21'd0}, _EVAL_3181};
  assign _EVAL_3060 = _EVAL_776[86];
  assign _EVAL_1187 = {_EVAL_519,_EVAL_2258};
  assign _EVAL_1665 = _EVAL_776[12];
  assign _EVAL_2481 = _EVAL_776[14];
  assign _EVAL_475 = _EVAL_2097 | _EVAL_1646;
  assign _EVAL_2846 = _EVAL_76 == 12'hb00;
  assign _EVAL_771 = _EVAL_2720 | _EVAL_1388;
  assign _EVAL_2299 = _EVAL_3068[1];
  assign _EVAL_3114 = _EVAL_236 | _EVAL_3005;
  assign _EVAL_2594 = _EVAL_2013[72];
  assign _EVAL_243 = _EVAL_772[12:11];
  assign _EVAL_2617 = _EVAL_279[5:0];
  assign _EVAL_1643 = _EVAL_76 == 12'hc1a;
  assign _EVAL_1843 = _EVAL_286 | _EVAL_3153;
  assign _EVAL_2443 = ~_EVAL_2148;
  assign _EVAL_2638 = {{135'd0}, _EVAL_274};
  assign _EVAL_1881 = _EVAL_1882[63:32];
  assign _EVAL_112 = _EVAL_762;
  assign _EVAL_2567 = _EVAL_2278 | _EVAL_93;
  assign _EVAL_245 = _EVAL_2203 ? 7'h43 : _EVAL_912;
  assign _EVAL_1195 = _EVAL_2258[6];
  assign _EVAL_1751 = _EVAL_2077 | _EVAL_18;
  assign _EVAL_56 = _EVAL_2445;
  assign _EVAL_1717 = _EVAL_101 == 12'h3b2;
  assign _EVAL_3036 = _EVAL_2787[0];
  assign _EVAL_2257 = _EVAL_2955 | _EVAL_716;
  assign _EVAL_2628 = _EVAL_3105 | _EVAL_2418;
  assign _EVAL_1746 = _EVAL_1549 ? 6'h2f : _EVAL_1020;
  assign _EVAL_2289 = _EVAL_776[75];
  assign _EVAL_799 = _EVAL_2958 & _EVAL_2262;
  assign _EVAL_417 = _EVAL_2567 ? _EVAL_190 : _EVAL_2147;
  assign _EVAL_24 = _EVAL_608;
  assign _EVAL_3099 = _EVAL_557 | _EVAL_2495;
  assign _EVAL_2944 = _EVAL_776[31];
  assign _EVAL_836 = _EVAL_177 | _EVAL_2070;
  assign _EVAL_804 = _EVAL_2263 | _EVAL_256;
  assign _EVAL_2285 = _EVAL_1963 | _EVAL_1321;
  assign _EVAL_1688 = _EVAL_1917 ? 8'h7 : _EVAL_1061;
  assign _EVAL_3165 = _EVAL_776[79];
  assign _EVAL_976 = _EVAL_1130 | _EVAL_1811;
  assign _EVAL_977 = _EVAL_776[23];
  assign _EVAL_294 = _EVAL_719 | _EVAL_1173;
  assign _EVAL_249 = _EVAL_2324 | _EVAL_2863;
  assign _EVAL_2866 = _EVAL_1517 | _EVAL_2058;
  assign _EVAL_27 = _EVAL_3183;
  assign _EVAL_2271 = _EVAL_776[121];
  assign _EVAL_2830 = _EVAL_2400 | _EVAL_2016;
  assign _EVAL_68 = _EVAL_333;
  assign _EVAL_1021 = _EVAL_591 ? 7'h62 : _EVAL_801;
  assign _EVAL_972 = _EVAL_2013[58];
  assign _EVAL_2803 = _EVAL_813 ? 6'h3f : _EVAL_2597;
  assign _EVAL_2511 = _EVAL_806 | _EVAL_2113;
  assign _EVAL_1404 = _EVAL_886[12];
  assign _EVAL_1957 = _EVAL_169 ? {{22'd0}, _EVAL_2479} : _EVAL_3254;
  assign _EVAL_2939 = _EVAL_2013[21];
  assign _EVAL_262 = _EVAL_1630 & _EVAL_2443;
  assign _EVAL_555 = _EVAL_101 == 12'h300;
  assign _EVAL_2668 = _EVAL_76 == 12'hb95;
  assign _EVAL_3136 = _EVAL_2858[7];
  assign _EVAL_2743 = 2'h3 == _EVAL_1512 ? _EVAL_819 : _EVAL_2767;
  assign _EVAL_911 = _EVAL_769 ? 8'h5 : _EVAL_2856;
  assign _EVAL_1107 = _EVAL_2469 | _EVAL_2567;
  assign _EVAL_237 = _EVAL_1772 ? 6'h2a : _EVAL_1190;
  assign _EVAL_3116 = 2'h2 == _EVAL_1512 ? _EVAL_2914 : _EVAL_1054;
  assign _EVAL_840 = _EVAL_1918 ? 8'h81 : _EVAL_1132;
  assign _EVAL_48 = _EVAL_935;
  assign _EVAL_1750 = _EVAL_3208 | _EVAL_1344;
  assign _EVAL_2042 = _EVAL_1852 | _EVAL_456;
  assign _EVAL_1395 = _EVAL_1659 ? 32'h3 : _EVAL_107;
  assign _EVAL_1992 = _EVAL_788 | _EVAL_1983;
  assign _EVAL_3037 = _EVAL_76 == 12'hb0c;
  assign _EVAL_956 = _EVAL_1543 ? 8'h71 : _EVAL_1343;
  assign _EVAL_2228 = _EVAL_776[3];
  assign _EVAL_1427 = _EVAL_169 & _EVAL_2927;
  assign _EVAL_2302 = _EVAL_2909 & _EVAL_42;
  assign _EVAL_1276 = _EVAL_2462 ? 8'h47 : _EVAL_198;
  assign _EVAL_1184 = _EVAL_799 | _EVAL_722;
  assign _EVAL_1469 = _EVAL_776[82];
  assign _EVAL_1020 = _EVAL_1315 ? 6'h2e : _EVAL_2656;
  assign _EVAL_743 = 2'h2 == _EVAL_1512 ? _EVAL_935 : _EVAL_2186;
  assign _EVAL_2208 = _EVAL_1331 & _EVAL_532;
  assign _EVAL_2977 = _EVAL_1931 | _EVAL_1064;
  assign _EVAL_114 = _EVAL_406;
  assign _EVAL_291 = _EVAL_2013[126];
  assign _EVAL_1283 = _EVAL_2975 ? 8'hc : _EVAL_904;
  assign _EVAL_402 = _EVAL_2779 | _EVAL_2607;
  assign _EVAL_1564 = _EVAL_1010 | _EVAL_415;
  assign _EVAL_889 = _EVAL_2617 == 6'h3;
  assign _EVAL_1181 = _EVAL_1716 ? 7'h4e : _EVAL_2344;
  assign _EVAL_2202 = _EVAL_899 | _EVAL_2836;
  assign _EVAL_982 = _EVAL_2587 | _EVAL_285;
  assign _EVAL_2199 = _EVAL_2698 | _EVAL_1716;
  assign _EVAL_2985 = _EVAL_544 | _EVAL_3000;
  assign _EVAL_714 = _EVAL_776[37];
  assign _EVAL_2814 = _EVAL_1528 ? 2'h3 : _EVAL_1936;
  assign _EVAL_2599 = _EVAL_341 & _EVAL_1280;
  assign _EVAL_2333 = _EVAL_1017 | _EVAL_588;
  assign _EVAL_2145 = _EVAL_76 == 12'hb0b;
  assign _EVAL_183 = _EVAL_1457 | _EVAL_798;
  assign _EVAL_226 = _EVAL_776[5];
  assign _EVAL_2876 = _EVAL_76 == 12'hb14;
  assign _EVAL_606 = _EVAL_776[124];
  assign _EVAL_3128 = _EVAL_2404 | _EVAL_2148;
  assign _EVAL_1202 = _EVAL_2787[1];
  assign _EVAL_3074 = _EVAL_776[66];
  assign _EVAL_1200 = _EVAL_1617 | _EVAL_1529;
  assign _EVAL_3065 = _EVAL_1729 & _EVAL_1508;
  assign _EVAL_94 = _EVAL_3213;
  assign _EVAL_2358 = {{111'd0}, _EVAL_620};
  assign _EVAL_2716 = _EVAL_1566 | _EVAL_3121;
  assign _EVAL_2185 = _EVAL_6[31:1];
  assign _EVAL_254 = _EVAL_2013[86];
  assign _EVAL_2318 = _EVAL_1996 | _EVAL_995;
  assign _EVAL_1106 = _EVAL_1525[8];
  assign _EVAL_1740 = _EVAL_1842 & _EVAL_2538;
  assign _EVAL_2704 = _EVAL_2124 | _EVAL_1469;
  assign _EVAL_2003 = _EVAL_2732[0];
  assign _EVAL_1742 = ~_EVAL_975;
  assign _EVAL_9 = _EVAL_1268;
  assign _EVAL_1464 = _EVAL_1533 == 2'h1;
  assign _EVAL_2519 = _EVAL_296[0];
  assign _EVAL_570 = _EVAL_1766 ? 7'h6a : _EVAL_567;
  assign _EVAL_157 = _EVAL_2013[88];
  assign _EVAL_2454 = _EVAL_2848 & _EVAL_3207;
  assign _EVAL_2928 = _EVAL_512 | _EVAL_260;
  assign _EVAL_1793 = _EVAL_555 ? _EVAL_1816 : 32'h0;
  assign _EVAL_1241 = _EVAL_1644 | _EVAL_196;
  assign _EVAL_2975 = _EVAL_1525[12];
  assign _EVAL_3007 = _EVAL_76 == 12'hc13;
  assign _EVAL_3091 = ~_EVAL_2020;
  assign _EVAL_179 = _EVAL_1463 | _EVAL_1362;
  assign _EVAL_1413 = _EVAL_1446 ? 8'he : _EVAL_3122;
  assign _EVAL_1974 = _EVAL_772[17];
  assign _EVAL_2470 = _EVAL_710 | _EVAL_226;
  assign _EVAL_1287 = _EVAL_2866 | _EVAL_910;
  assign _EVAL_2388 = {{111'd0}, _EVAL_2258};
  assign _EVAL_629 = _EVAL_1462 ? 7'h68 : _EVAL_1975;
  assign _EVAL_1277 = _EVAL_2567 ? _EVAL_1957 : {{22'd0}, _EVAL_2479};
  assign _EVAL_2653 = _EVAL_1393 | _EVAL_2831;
  assign _EVAL_1868 = {_EVAL_2387,_EVAL_153,_EVAL_2158,_EVAL_2356};
  assign _EVAL_387 = ~_EVAL_2614;
  assign _EVAL_1866 = _EVAL_2418 ? 7'h7d : _EVAL_2645;
  assign _EVAL_563 = _EVAL_1847 ? 8'h64 : _EVAL_3131;
  assign _EVAL_3033 = 2'h0 == _EVAL_1512;
  assign _EVAL_675 = ~_EVAL_891;
  assign _EVAL_2978 = _EVAL_1942 | _EVAL_1397;
  assign _EVAL_2898 = _EVAL_2868 | _EVAL_2123;
  assign _EVAL_1530 = _EVAL_3134 ? _EVAL_2258 : {{2'd0}, _EVAL_1279};
  assign _EVAL_2072 = _EVAL_3048 | _EVAL_824;
  assign _EVAL_1966 = _EVAL_1771 & _EVAL_2394;
  assign _EVAL_781 = _EVAL_2013[56];
  assign _EVAL_740 = _EVAL_524 | _EVAL_2933;
  assign _EVAL_2133 = _EVAL_362 | _EVAL_583;
  assign _EVAL_2659 = _EVAL_2305 ? _EVAL_2085 : _EVAL_509;
  assign _EVAL_3082 = _EVAL_2364 ? 7'h5f : _EVAL_2340;
  assign _EVAL_1901 = _EVAL_1681 ? _EVAL_1244 : {{57'd0}, _EVAL_251};
  assign _EVAL_2767 = 2'h2 == _EVAL_1512 ? _EVAL_1268 : _EVAL_1989;
  assign _EVAL_409 = _EVAL_1890 ? 8'h5d : _EVAL_2048;
  assign _EVAL_1783 = _EVAL_2431 | _EVAL_445;
  assign _EVAL_1224 = _EVAL_1063 | _EVAL_970;
  assign _EVAL_1519 = _EVAL_932 | _EVAL_909;
  assign _EVAL_448 = _EVAL_2228 ? 4'h3 : _EVAL_2480;
  assign _EVAL_948 = {{135'd0}, _EVAL_1379};
  assign _EVAL_2048 = _EVAL_193 ? 8'h5c : _EVAL_706;
  assign _EVAL_1676 = _EVAL_2858[4:3];
  assign _EVAL_2188 = _EVAL_970 ? 6'h24 : _EVAL_453;
  assign _EVAL_1927 = _EVAL_3173 | _EVAL_594;
  assign _EVAL_1596 = _EVAL_776[111];
  assign _EVAL_474 = _EVAL_2327 | _EVAL_967;
  assign _EVAL_1479 = _EVAL_2760 & _EVAL_308;
  assign _EVAL_420 = _EVAL_1873 ? 8'h7c : _EVAL_2156;
  assign _EVAL_181 = _EVAL_76 == 12'h328;
  assign _EVAL_1887 = _EVAL_1796 ? 2'h3 : 2'h0;
  assign _EVAL_2115 = _EVAL_969 | _EVAL_2703;
  assign _EVAL_3117 = _EVAL_2013[50];
  assign _EVAL_2340 = _EVAL_164 ? 7'h5e : _EVAL_773;
  assign _EVAL_3157 = _EVAL_76 == 12'hb08;
  assign _EVAL_2953 = _EVAL_2903 | _EVAL_554;
  assign _EVAL_684 = _EVAL_1356 ? 8'h18 : _EVAL_301;
  assign _EVAL_751 = _EVAL_2388 & 143'h7fffffffffffffffffffffffffffffff0888;
  assign _EVAL_54 = _EVAL_3242;
  assign _EVAL_589 = {_EVAL_2799,_EVAL_918};
  assign _EVAL_1724 = _EVAL_1928 ? 8'h65 : _EVAL_563;
  assign _EVAL_2705 = _EVAL_1097[63:6];
  assign _EVAL_978 = _EVAL_2818 | _EVAL_883;
  assign _EVAL_2233 = _EVAL_776[45];
  assign _EVAL_1293 = _EVAL_2428 ? 8'h31 : _EVAL_2946;
  assign _EVAL_1587 = {_EVAL_531,2'h3};
  assign _EVAL_2414 = _EVAL_3040 == 32'h100000;
  assign _EVAL_1636 = _EVAL_2013[83];
  assign _EVAL_2614 = _EVAL_2824 ? _EVAL_18 : 32'h0;
  assign _EVAL_2381 = _EVAL_2166 | _EVAL_866;
  assign _EVAL_2877 = _EVAL_836 | _EVAL_2106;
  assign _EVAL_2407 = _EVAL_76 == 12'hb06;
  assign _EVAL_103 = _EVAL_2406;
  assign _EVAL_1298 = _EVAL_2466 | _EVAL_2731;
  assign _EVAL_3208 = _EVAL_2348 | _EVAL_1762;
  assign _EVAL_2360 = _EVAL_1412 | _EVAL_1429;
  assign _EVAL_2294 = _EVAL_76 == 12'h3b9;
  assign _EVAL_1474 = _EVAL_1382 | _EVAL_1306;
  assign _EVAL_798 = _EVAL_2013[67];
  assign _EVAL_1611 = _EVAL_477 | _EVAL_2233;
  assign _EVAL_2833 = _EVAL_2678 ? 7'h4c : _EVAL_938;
  assign _EVAL_1071 = _EVAL_101 == 12'h7a0;
  assign _EVAL_2274 = _EVAL_776[7];
  assign _EVAL_560 = _EVAL_2960 ? _EVAL_1238 : 32'h0;
  assign _EVAL_926 = 2'h3 == _EVAL_1512 ? _EVAL_1595 : _EVAL_2151;
  assign _EVAL_126 = _EVAL_2542;
  assign _EVAL_1472 = _EVAL_1700 ? _EVAL_2516 : _EVAL_2993;
  assign _EVAL_1660 = _EVAL_76 == 12'hb0a;
  assign _EVAL_957 = _EVAL_690 ? 4'hf : _EVAL_1677;
  assign _EVAL_970 = _EVAL_776[36];
  assign _EVAL_1799 = _EVAL_843 | _EVAL_996;
  assign _EVAL_2108 = _EVAL_2602 ? _EVAL_2369 : 32'h0;
  assign _EVAL_1579 = 2'h2 == _EVAL_1512 ? _EVAL_1080 : _EVAL_1081;
  assign _EVAL_1387 = _EVAL_2848 & _EVAL_525;
  assign _EVAL_2525 = _EVAL_1749 ? 8'h86 : _EVAL_565;
  assign _EVAL_1659 = _EVAL_2330 & _EVAL_2414;
  assign _EVAL_11 = _EVAL_484;
  assign _EVAL_2529 = _EVAL_3117 ? 8'h32 : _EVAL_1293;
  assign _EVAL_1446 = _EVAL_2013[14];
  assign _EVAL_330 = _EVAL_1030 ? 8'h22 : _EVAL_1501;
  assign _EVAL_2258 = _EVAL_3006 & _EVAL_387;
  assign _EVAL_2501 = _EVAL_101 == 12'hb02;
  assign _EVAL_1621 = _EVAL_1940[11];
  assign _EVAL_457 = _EVAL_2013[53];
  assign _EVAL_3059 = _EVAL_672 | _EVAL_1730;
  assign _EVAL_653 = _EVAL_386 ? 1'h0 : _EVAL_525;
  assign _EVAL_1646 = _EVAL_76 == 12'hb15;
  assign _EVAL_2615 = _EVAL_335 | _EVAL_193;
  assign _EVAL_2452 = _EVAL_2065 | _EVAL_2927;
  assign _EVAL_47 = {{1'd0}, _EVAL_3152};
  assign _EVAL_2904 = _EVAL_2647 | _EVAL_103;
  assign _EVAL_1175 = _EVAL_966 | _EVAL_707;
  assign _EVAL_3040 = _EVAL_1739 & 32'h10100000;
  assign _EVAL_1925 = _EVAL_776[91];
  assign _EVAL_801 = _EVAL_1173 ? 7'h61 : _EVAL_1484;
  assign _EVAL_2696 = _EVAL_76 == 12'hc15;
  assign _EVAL_851 = ~_EVAL_2842;
  assign _EVAL_2410 = _EVAL_776[129];
  assign _EVAL_905 = _EVAL_2509 | _EVAL_2881;
  assign _EVAL_667 = _EVAL_3250 ? 5'h10 : {{1'd0}, _EVAL_957};
  assign _EVAL_1919 = _EVAL_1525[13];
  assign _EVAL_2622 = _EVAL_457 ? 8'h35 : _EVAL_2201;
  assign _EVAL_2580 = _EVAL_2013[8];
  assign _EVAL_1678 = _EVAL_209 | _EVAL_1233;
  assign _EVAL_2385 = _EVAL_2988 | _EVAL_232;
  assign _EVAL_1941 = _EVAL_746 + 58'h1;
  assign _EVAL_3245 = _EVAL_776[77];
  assign _EVAL_3063 = _EVAL_101 == 12'h345;
  assign _EVAL_21 = _EVAL_1172 & _EVAL_526;
  assign _EVAL_2218 = _EVAL_76 == 12'hc09;
  assign _EVAL_446 = _EVAL_2330 & _EVAL_727;
  assign _EVAL_2166 = _EVAL_1895 | _EVAL_2884;
  assign _EVAL_1600 = _EVAL_1114 ? _EVAL_412 : 32'h0;
  assign _EVAL_1212 = _EVAL_2013[44];
  assign _EVAL_2988 = _EVAL_2008 | _EVAL_2838;
  assign _EVAL_1459 = _EVAL_3140 | _EVAL_861;
  assign _EVAL_1764 = _EVAL_3106 | _EVAL_328;
  assign _EVAL_1637 = _EVAL_776[51];
  assign _EVAL_1580 = {{111'd0}, _EVAL_726};
  assign _EVAL_2752 = {_EVAL_12,_EVAL_58,_EVAL_28,_EVAL_2,_EVAL_126,_EVAL_118,_EVAL_69};
  assign _EVAL_716 = _EVAL_76 == 12'hc0d;
  assign _EVAL_1367 = _EVAL_2013[26];
  assign _EVAL_1381 = _EVAL_486 ? 7'h75 : _EVAL_1338;
  assign _EVAL_1513 = _EVAL_1295 & _EVAL_2647;
  assign _EVAL_2134 = _EVAL_2396 | _EVAL_671;
  assign _EVAL_3029 = _EVAL_1665 ? 4'hc : _EVAL_1694;
  assign _EVAL_1130 = _EVAL_1383 | _EVAL_1439;
  assign _EVAL_870 = _EVAL_546 | _EVAL_1844;
  assign _EVAL_1045 = _EVAL_2573 | _EVAL_2616;
  assign _EVAL_985 = _EVAL_101 == 12'h7a2;
  assign _EVAL_1223 = 2'h2 == _EVAL_1512 ? _EVAL_608 : _EVAL_187;
  assign _EVAL_910 = _EVAL_76 == 12'hc84;
  assign _EVAL_737 = _EVAL_270 ? 8'h37 : _EVAL_586;
  assign _EVAL_1418 = _EVAL_1589 | _EVAL_2972;
  assign _EVAL_2304 = _EVAL_1941[57:0];
  assign _EVAL_1365 = _EVAL_76 == 12'hc96;
  assign _EVAL_2058 = _EVAL_76 == 12'hb84;
  assign _EVAL_3076 = _EVAL_3089 & 32'h20400000;
  assign _EVAL_1001 = _EVAL_2223 | _EVAL_3127;
  assign _EVAL_2433 = _EVAL_2666 | _EVAL_2490;
  assign _EVAL_2896 = _EVAL_1095 ? _EVAL_388 : 32'h0;
  assign _EVAL_208 = _EVAL_76 == 12'hc8c;
  assign _EVAL_1935 = {_EVAL_2159,_EVAL_2258};
  assign _EVAL_2305 = _EVAL_108 != 8'h0;
  assign _EVAL_1327 = _EVAL_1642 ? 8'h1c : _EVAL_155;
  assign _EVAL_1546 = _EVAL_76 == 12'hc02;
  assign _EVAL_966 = _EVAL_1039 | _EVAL_1133;
  assign _EVAL_1862 = _EVAL_2258[3];
  assign _EVAL_2440 = _EVAL_212 ? 6'h21 : _EVAL_2122;
  assign _EVAL_230 = _EVAL_76 == 12'hb82;
  assign _EVAL_2416 = _EVAL_76 == 12'hc9a;
  assign _EVAL_1715 = _EVAL_2729 ? 7'h51 : _EVAL_2451;
  assign _EVAL_1360 = _EVAL_808 ? 8'h73 : _EVAL_1093;
  assign _EVAL_1795 = _EVAL_1125 | _EVAL_422;
  assign _EVAL_1070 = {{79'd0}, _EVAL_1255};
  assign _EVAL_227 = _EVAL_76 == 12'h3b0;
  assign _EVAL_35 = _EVAL_2784;
  assign _EVAL_1300 = _EVAL_982 | _EVAL_2346;
  assign _EVAL_1393 = _EVAL_2544 | _EVAL_2428;
  assign _EVAL_902 = _EVAL_76 == 12'hc10;
  assign _EVAL_599 = 143'h0;
  assign _EVAL_26 = _EVAL_51;
  assign _EVAL_2738 = _EVAL_1177 ? 8'h8c : _EVAL_2284;
  assign _EVAL_1411 = _EVAL_1350 | _EVAL_1090;
  assign _EVAL_2434 = 2'h3 == _EVAL_1512 ? _EVAL_1850 : _EVAL_1579;
  assign _EVAL_1422 = _EVAL_1739 & 32'h20100000;
  assign _EVAL_1350 = _EVAL_430 | _EVAL_1541;
  assign _EVAL_2735 = _EVAL_285 ? 8'h8d : _EVAL_2169;
  assign _EVAL_2993 = _EVAL_550 ? _EVAL_1935 : {{57'd0}, _EVAL_397};
  assign _EVAL_1154 = _EVAL_1525[14];
  assign _EVAL_1158 = _EVAL_468 | _EVAL_639;
  assign _EVAL_1421 = ~_EVAL_2550;
  assign _EVAL_364 = _EVAL_543 ? 6'h35 : _EVAL_444;
  assign _EVAL_1772 = _EVAL_776[42];
  assign _EVAL_1208 = _EVAL_2013[95];
  assign _EVAL_2178 = _EVAL_263 ? 7'h7f : _EVAL_2648;
  assign _EVAL_3011 = _EVAL_2895[7:5];
  assign _EVAL_380 = _EVAL_2013[7];
  assign _EVAL_711 = ~_EVAL_1319;
  assign _EVAL_981 = _EVAL_2761 ? 8'h3d : _EVAL_2627;
  assign _EVAL_273 = _EVAL_2848 ? 1'h0 : _EVAL_0;
  assign _EVAL_1121 = _EVAL_2013[25];
  assign _EVAL_1488 = _EVAL_447 | _EVAL_1892;
  assign _EVAL_2757 = _EVAL_76 == 12'h32e;
  assign _EVAL_2581 = _EVAL_2806 | _EVAL_1823;
  assign _EVAL_497 = _EVAL_1681 ? _EVAL_1558 : {{2'd0}, _EVAL_333};
  assign _EVAL_2201 = _EVAL_2657 ? 8'h34 : _EVAL_649;
  assign _EVAL_97 = _EVAL_845;
  assign _EVAL_256 = _EVAL_776[32];
  assign _EVAL_2441 = _EVAL_277 ? 8'h6a : _EVAL_1473;
  assign _EVAL_1781 = _EVAL_1551 | _EVAL_1070;
  assign _EVAL_92 = _EVAL_729;
  assign _EVAL_550 = _EVAL_101 == 12'hb00;
  assign _EVAL_1372 = _EVAL_1079 & _EVAL_2702;
  assign _EVAL_2276 = _EVAL_76 == 12'hc1d;
  assign _EVAL_435 = _EVAL_1679 | _EVAL_1203;
  assign _EVAL_2170 = _EVAL_2229 & _EVAL_2647;
  assign _EVAL_1955 = _EVAL_1707 ? 8'h3 : _EVAL_2755;
  assign _EVAL_483 = _EVAL_2347 | _EVAL_925;
  assign _EVAL_2161 = _EVAL_2433 | _EVAL_230;
  assign _EVAL_1189 = _EVAL_776[61];
  assign _EVAL_2061 = _EVAL_2013[85];
  assign _EVAL_1548 = _EVAL_1616 ? 8'h8e : _EVAL_2735;
  assign _EVAL_964 = _EVAL_686 | _EVAL_2558;
  assign _EVAL_2769 = _EVAL_2317[31:0];
  assign _EVAL_2124 = _EVAL_2493 | _EVAL_2917;
  assign _EVAL_1571 = _EVAL_2772 ? 8'h6f : _EVAL_3051;
  assign _EVAL_1848 = _EVAL_1321 ? 8'h84 : _EVAL_2902;
  assign _EVAL_152 = _EVAL_1721[39:6];
  assign _EVAL_1951 = _EVAL_475 | _EVAL_2696;
  assign _EVAL_3167 = _EVAL_776[18];
  assign _EVAL_2488 = _EVAL_2741 ? 8'h5 : _EVAL_775;
  assign _EVAL_3156 = _EVAL_76 == 12'hc98;
  assign _EVAL_486 = _EVAL_776[117];
  assign _EVAL_941 = _EVAL_985 ? _EVAL_1905 : 32'h0;
  assign _EVAL_1335 = _EVAL_1675 | _EVAL_2310;
  assign _EVAL_542 = _EVAL_157 ? 8'h58 : _EVAL_1058;
  assign _EVAL_567 = _EVAL_314 ? 7'h69 : _EVAL_629;
  assign _EVAL_786 = _EVAL_1235 ? 5'h15 : _EVAL_1094;
  assign _EVAL_1201 = _EVAL_2047 | _EVAL_2289;
  assign _EVAL_38 = 2'h0;
  assign _EVAL_1682 = _EVAL_76 == 12'hc8a;
  assign _EVAL_776 = _EVAL_408 ? _EVAL_1924 : 143'h0;
  assign _EVAL_1520 = _EVAL_2940 | _EVAL_2358;
  assign _EVAL_2094 = {{111'd0}, _EVAL_290};
  assign _EVAL_1063 = _EVAL_650 | _EVAL_714;
  assign _EVAL_1829 = _EVAL_2802 | _EVAL_2975;
  assign _EVAL_1978 = _EVAL_76 == 12'h3b7;
  assign _EVAL_822 = _EVAL_76 == 12'hc04;
  assign _EVAL_702 = _EVAL_2013[76];
  assign _EVAL_531 = _EVAL_589 & _EVAL_522;
  assign _EVAL_2062 = _EVAL_1851 | _EVAL_1604;
  assign _EVAL_78 = _EVAL_3115;
  assign _EVAL_2890 = _EVAL_2588 | _EVAL_1385;
  assign _EVAL_2861 = {{103'd0}, _EVAL_576};
  assign _EVAL_3129 = _EVAL_1136 | _EVAL_18;
  assign _EVAL_3110 = _EVAL_2193 ? _EVAL_459 : 32'h0;
  assign _EVAL_1065 = _EVAL_1892 ? 7'h44 : _EVAL_245;
  assign _EVAL_2419 = _EVAL_3018 ? 8'h8d : _EVAL_2738;
  assign _EVAL_3148 = _EVAL_101 == 12'h307;
  assign _EVAL_1408 = _EVAL_886[27];
  assign _EVAL_1773 = _EVAL_2858[2];
  assign _EVAL_1337 = _EVAL_327 ? 8'h40 : _EVAL_1225;
  assign _EVAL_1500 = {{79'd0}, _EVAL_1737};
  assign _EVAL_1800 = _EVAL_2215[3:0];
  assign _EVAL_2217 = _EVAL_2013[81];
  assign _EVAL_1697 = _EVAL_3115 | _EVAL_845;
  assign _EVAL_425 = _EVAL_49 & _EVAL_2293;
  assign _EVAL_785 = _EVAL_2543 | _EVAL_693;
  assign _EVAL_28 = _EVAL_2375;
  assign _EVAL_1998 = _EVAL_1882[31:0];
  assign _EVAL_2796 = _EVAL_3182 | _EVAL_691;
  assign _EVAL_1863 = {_EVAL_1279,_EVAL_1720};
  assign _EVAL_1429 = _EVAL_2013[20];
  assign _EVAL_236 = _EVAL_2463 | _EVAL_2757;
  assign _EVAL_1838 = _EVAL_971 ? 8'h76 : _EVAL_683;
  assign _EVAL_2123 = _EVAL_776[142];
  assign _EVAL_1463 = _EVAL_1588 | _EVAL_2098;
  assign _EVAL_2793 = _EVAL_76 == 12'hb07;
  assign _EVAL_3180 = _EVAL_853 != 8'he;
  assign _EVAL_1604 = _EVAL_776[34];
  assign _EVAL_196 = _EVAL_76 == 12'h33a;
  assign _EVAL_1032 = _EVAL_3063 ? _EVAL_1816 : _EVAL_34;
  assign _EVAL_2789 = _EVAL_101 == 12'h3b1;
  assign _EVAL_581 = {_EVAL_746,_EVAL_2644};
  assign _EVAL_2046 = _EVAL_2061 ? 8'h55 : _EVAL_2092;
  assign _EVAL_2827 = _EVAL_312 | _EVAL_1918;
  assign _EVAL_912 = _EVAL_3074 ? 7'h42 : _EVAL_1018;
  assign _EVAL_1403 = _EVAL_1414 ? 6'h2 : 6'h3c;
  assign _EVAL_835 = _EVAL_2330 & _EVAL_1380;
  assign _EVAL_897 = _EVAL_2909 ? _EVAL_55 : _EVAL_2311;
  assign _EVAL_1898 = _EVAL_101 == 12'h346;
  assign _EVAL_1573 = _EVAL_1478 | _EVAL_280;
  assign _EVAL_2941 = _EVAL_3034 | _EVAL_1027;
  assign _EVAL_2662 = _EVAL_2225 ? 7'h59 : _EVAL_950;
  assign _EVAL_428 = _EVAL_441 | _EVAL_625;
  assign _EVAL_537 = _EVAL_978 | _EVAL_390;
  assign _EVAL_1620 = _EVAL_2848 ? _EVAL_820 : 2'h0;
  assign _EVAL_1518 = _EVAL_1325 | _EVAL_265;
  assign _EVAL_1532 = _EVAL_76 & 12'hc10;
  assign _EVAL_104 = 2'h1;
  assign _EVAL_2899 = _EVAL_1466 | _EVAL_345;
  assign _EVAL_2239 = _EVAL_3070 + _EVAL_3095;
  assign _EVAL_2014 = _EVAL_1764 | _EVAL_1864;
  assign _EVAL_301 = _EVAL_2733 ? 8'h17 : _EVAL_2996;
  assign _EVAL_1996 = _EVAL_2819 | _EVAL_1614;
  assign _EVAL_2382 = _EVAL_210 | _EVAL_316;
  assign _EVAL_2698 = _EVAL_2506 | _EVAL_3165;
  assign _EVAL_849 = _EVAL_2135 ? 7'h5c : _EVAL_2171;
  assign _EVAL_125 = _EVAL_924;
  assign _EVAL_2845 = ~_EVAL_845;
  assign _EVAL_605 = _EVAL_641 ? 8'h87 : _EVAL_2067;
  assign _EVAL_2513 = _EVAL_76 == 12'hc87;
  assign _EVAL_1061 = _EVAL_946 ? 8'h9 : _EVAL_2834;
  assign _EVAL_1672 = _EVAL_76 == 12'hb93;
  assign _EVAL_2405 = _EVAL_368 ? {{22'd0}, _EVAL_1683} : _EVAL_1277;
  assign _EVAL_3198 = _EVAL_562 | _EVAL_1499;
  assign _EVAL_357 = _EVAL_1525[1];
  assign _EVAL_2359 = _EVAL_1735 & _EVAL_3207;
  assign _EVAL_215 = _EVAL_841 ? _EVAL_1721 : _EVAL_2937;
  assign _EVAL_1035 = _EVAL_1455 ? 8'h10 : _EVAL_1510;
  assign _EVAL_305 = _EVAL_326 | _EVAL_779;
  assign _EVAL_2888 = {4'h2,_EVAL_975,14'h400,_EVAL_3058,_EVAL_192,2'h0,_EVAL_1142,_EVAL_1759};
  assign _EVAL_3203 = _EVAL_2258[0];
  assign _EVAL_1177 = _EVAL_776[140];
  assign _EVAL_2651 = ~_EVAL_2258;
  assign _EVAL_1190 = _EVAL_1415 ? 6'h29 : _EVAL_1218;
  assign _EVAL_2991 = _EVAL_3147 & _EVAL_3091;
  assign _EVAL_2485 = _EVAL_76 == 12'h3be;
  assign _EVAL_895 = _EVAL_776[122];
  assign _EVAL_1108 = _EVAL_2978 | _EVAL_1030;
  assign _EVAL_1758 = _EVAL_884 | _EVAL_2681;
  assign _EVAL_2709 = _EVAL_2072 | _EVAL_730;
  assign _EVAL_2744 = _EVAL_2929 & _EVAL_2659;
  assign _EVAL_1412 = _EVAL_505 | _EVAL_2939;
  assign _EVAL_2352 = 2'h1 == _EVAL_1512 ? _EVAL_1047 : _EVAL_2689;
  assign _EVAL_1975 = _EVAL_1366 ? 7'h67 : _EVAL_645;
  assign _EVAL_2949 = _EVAL_2848 & _EVAL_1948;
  assign _EVAL_690 = _EVAL_776[15];
  assign _EVAL_1280 = _EVAL_1331 | _EVAL_745;
  assign _EVAL_646 = _EVAL_1286 | _EVAL_947;
  assign _EVAL_4 = _EVAL_880;
  assign _EVAL_3201 = _EVAL_1189 ? 6'h3d : _EVAL_1970;
  assign _EVAL_641 = _EVAL_776[135];
  assign _EVAL_25 = _EVAL_2799;
  assign _EVAL_3235 = _EVAL_758 ? 1'h0 : _EVAL_1353;
  assign _EVAL_3236 = _EVAL_2039 | _EVAL_2380;
  assign _EVAL_1322 = _EVAL_2929 | _EVAL_2041;
  assign _EVAL_329 = _EVAL_1909 | _EVAL_2061;
  assign _EVAL_2335 = 2'h1 == _EVAL_1512 ? _EVAL_2907 : _EVAL_1493;
  assign _EVAL_1816 = _EVAL_1814[31:0];
  assign _EVAL_14 = _EVAL_1466;
  assign _EVAL_1229 = _EVAL_3080 + _EVAL_770;
  assign _EVAL_639 = _EVAL_76 == 12'hb9c;
  assign _EVAL_768 = _EVAL_1203 ? 5'h1e : _EVAL_2222;
  assign _EVAL_1707 = _EVAL_2013[3];
  assign _EVAL_2221 = _EVAL_1264 | _EVAL_457;
  assign _EVAL_1401 = _EVAL_291 ? 8'h7e : _EVAL_244;
  assign _EVAL_1112 = _EVAL_568 ? 8'h60 : _EVAL_2989;
  assign _EVAL_162 = _EVAL_776[90];
  assign _EVAL_1310 = _EVAL_3068[0];
  assign _EVAL_2545 = _EVAL_1966 ? {{24'd0}, _EVAL_55} : _EVAL_2405;
  assign _EVAL_2477 = _EVAL_724 | _EVAL_2236;
  assign _EVAL_2031 = _EVAL_169 ? {{1'd0}, _EVAL_3052} : _EVAL_266;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_153 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_156 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_163 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_178 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_192 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_261 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_269 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_272 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_279 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_315 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_331 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_333 = _RAND_11[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_334 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_406 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_429 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_438 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_440 = _RAND_16[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_459 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_484 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_494 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_495 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_507 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_525 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_608 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_612 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_619 = _RAND_25[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_673 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_685 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_699 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_728 = _RAND_29[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_729 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  _EVAL_746 = _RAND_31[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_753 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_762 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_767 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_774 = _RAND_35[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_819 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_820 = _RAND_37[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _EVAL_845 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _EVAL_850 = _RAND_39[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _EVAL_864 = _RAND_40[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _EVAL_880 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _EVAL_891 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _EVAL_908 = _RAND_43[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _EVAL_920 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _EVAL_924 = _RAND_45[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _EVAL_935 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _EVAL_975 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _EVAL_1019 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _EVAL_1047 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _EVAL_1080 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _EVAL_1142 = _RAND_51[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _EVAL_1172 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _EVAL_1239 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _EVAL_1246 = _RAND_54[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _EVAL_1267 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _EVAL_1268 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _EVAL_1271 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _EVAL_1279 = _RAND_58[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _EVAL_1318 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _EVAL_1351 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _EVAL_1353 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _EVAL_1447 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _EVAL_1450 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _EVAL_1451 = _RAND_64[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _EVAL_1466 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _EVAL_1467 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _EVAL_1491 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _EVAL_1493 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _EVAL_1507 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _EVAL_1512 = _RAND_70[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _EVAL_1595 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _EVAL_1608 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _EVAL_1722 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _EVAL_1755 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _EVAL_1850 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _EVAL_1888 = _RAND_76[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _EVAL_1948 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {2{`RANDOM}};
  _EVAL_1969 = _RAND_78[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _EVAL_2083 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _EVAL_2129 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _EVAL_2147 = _RAND_81[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _EVAL_2148 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _EVAL_2158 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _EVAL_2251 = _RAND_84[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _EVAL_2268 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _EVAL_2306 = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _EVAL_2349 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _EVAL_2355 = _RAND_88[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _EVAL_2356 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _EVAL_2375 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _EVAL_2380 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _EVAL_2387 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _EVAL_2392 = _RAND_93[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _EVAL_2406 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _EVAL_2445 = _RAND_95[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _EVAL_2471 = _RAND_96[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _EVAL_2479 = _RAND_97[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _EVAL_2486 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _EVAL_2542 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _EVAL_2579 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _EVAL_2593 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _EVAL_2609 = _RAND_102[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _EVAL_2644 = _RAND_103[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _EVAL_2647 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _EVAL_2654 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _EVAL_2665 = _RAND_106[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _EVAL_2673 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _EVAL_2674 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _EVAL_2676 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _EVAL_2689 = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _EVAL_2708 = _RAND_111[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _EVAL_2732 = _RAND_112[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _EVAL_2764 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _EVAL_2784 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _EVAL_2791 = _RAND_115[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _EVAL_2799 = _RAND_116[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _EVAL_2828 = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _EVAL_2842 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _EVAL_2844 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _EVAL_2870 = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _EVAL_2907 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _EVAL_2914 = _RAND_122[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _EVAL_2927 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _EVAL_2931 = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _EVAL_2987 = _RAND_125[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _EVAL_3052 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _EVAL_3058 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _EVAL_3068 = _RAND_128[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _EVAL_3070 = _RAND_129[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _EVAL_3115 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _EVAL_3143 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _EVAL_3152 = _RAND_132[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _EVAL_3170 = _RAND_133[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _EVAL_3183 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _EVAL_3184 = _RAND_135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _EVAL_3195 = _RAND_136[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _EVAL_3213 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _EVAL_3217 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _EVAL_3231 = _RAND_139[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {2{`RANDOM}};
  _EVAL_3239 = _RAND_140[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _EVAL_3242 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _EVAL_3256 = _RAND_142[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_16) begin
    if (_EVAL_63) begin
      _EVAL_153 <= 1'h0;
    end
    if (_EVAL_1681) begin
      if (_EVAL_1146) begin
        _EVAL_156 <= _EVAL_2740;
      end else if (_EVAL_2567) begin
        if (!(_EVAL_169)) begin
          _EVAL_156 <= _EVAL_1421;
        end
      end
    end else if (_EVAL_2567) begin
      if (!(_EVAL_169)) begin
        _EVAL_156 <= _EVAL_1421;
      end
    end
    if (_EVAL_63) begin
      _EVAL_163 <= 1'h0;
    end
    if (_EVAL_63) begin
      _EVAL_178 <= 32'h0;
    end
    if (_EVAL_63) begin
      _EVAL_192 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1424) begin
        if (_EVAL_1619) begin
          _EVAL_192 <= _EVAL_2599;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_261 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2429) begin
        _EVAL_261 <= _EVAL_1974;
      end
    end
    if (_EVAL_63) begin
      _EVAL_269 <= 1'h0;
    end
    if (_EVAL_63) begin
      _EVAL_272 <= 1'h0;
    end
    if (_EVAL_63) begin
      _EVAL_279 <= 32'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2670) begin
        if (_EVAL_264) begin
          _EVAL_279 <= _EVAL_2258;
        end else begin
          _EVAL_279 <= _EVAL_432;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_315 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1658) begin
        if (_EVAL_1619) begin
          _EVAL_315 <= _EVAL_3203;
        end
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_559) begin
        _EVAL_331 <= _EVAL_1773;
      end
    end
    _EVAL_333 <= _EVAL_497[29:0];
    if (_EVAL_63) begin
      _EVAL_334 <= 1'h0;
    end
    if (_EVAL_1681) begin
      if (_EVAL_1150) begin
        _EVAL_406 <= _EVAL_399;
      end
    end
    if (_EVAL_63) begin
      _EVAL_429 <= 6'h0;
    end
    if (_EVAL_63) begin
      _EVAL_438 <= 2'h0;
    end
    if (_EVAL_63) begin
      _EVAL_440 <= 2'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2429) begin
        _EVAL_440 <= 2'h0;
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_2193) begin
        _EVAL_459 <= _EVAL_2258;
      end
    end
    if (_EVAL_63) begin
      _EVAL_484 <= 1'h0;
    end
    if (_EVAL_1681) begin
      if (_EVAL_559) begin
        _EVAL_494 <= _EVAL_1956;
      end
    end
    if (_EVAL_63) begin
      _EVAL_495 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1658) begin
        if (_EVAL_1619) begin
          _EVAL_495 <= _EVAL_1062;
        end
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_1150) begin
        _EVAL_507 <= _EVAL_297;
      end
    end
    if (_EVAL_63) begin
      _EVAL_525 <= 1'h0;
    end else begin
      _EVAL_525 <= _EVAL_207;
    end
    if (_EVAL_63) begin
      _EVAL_608 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2117) begin
        if (_EVAL_1619) begin
          _EVAL_608 <= _EVAL_228;
        end
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_2117) begin
        if (_EVAL_1619) begin
          _EVAL_612 <= _EVAL_1195;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_619 <= 12'h0;
    end
    if (_EVAL_1681) begin
      if (_EVAL_559) begin
        _EVAL_673 <= _EVAL_2378;
      end
    end
    if (_EVAL_63) begin
      _EVAL_685 <= 1'h0;
    end
    if (_EVAL_1681) begin
      if (_EVAL_2968) begin
        _EVAL_699 <= _EVAL_2621;
      end
    end
    if (_EVAL_63) begin
      _EVAL_728 <= 3'h0;
    end
    if (_EVAL_1681) begin
      if (_EVAL_2968) begin
        _EVAL_729 <= _EVAL_3036;
      end
    end
    if (_EVAL_63) begin
      _EVAL_746 <= 58'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1700) begin
        _EVAL_746 <= _EVAL_2841;
      end else if (_EVAL_550) begin
        _EVAL_746 <= _EVAL_2315;
      end else if (_EVAL_340) begin
        _EVAL_746 <= _EVAL_2304;
      end
    end else if (_EVAL_340) begin
      _EVAL_746 <= _EVAL_2304;
    end
    if (_EVAL_63) begin
      _EVAL_753 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1424) begin
        if (_EVAL_1619) begin
          _EVAL_753 <= _EVAL_3203;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_762 <= 1'h0;
    end
    if (_EVAL_1681) begin
      if (_EVAL_1114) begin
        _EVAL_767 <= _EVAL_2258;
      end
    end
    if (_EVAL_63) begin
      _EVAL_774 <= 2'h0;
    end
    if (_EVAL_63) begin
      _EVAL_819 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1658) begin
        if (_EVAL_1619) begin
          _EVAL_819 <= _EVAL_1303;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_820 <= 2'h3;
    end else if (_EVAL_1681) begin
      if (_EVAL_368) begin
        if (_EVAL_2848) begin
          _EVAL_820 <= _EVAL_1248;
        end else if (_EVAL_2429) begin
          if (_EVAL_2747) begin
            _EVAL_820 <= 2'h3;
          end else begin
            _EVAL_820 <= 2'h0;
          end
        end else if (_EVAL_1117) begin
          if (_EVAL_1083) begin
            if (_EVAL_2567) begin
              if (!(_EVAL_169)) begin
                if (_EVAL_1796) begin
                  _EVAL_820 <= 2'h3;
                end else begin
                  _EVAL_820 <= 2'h0;
                end
              end
            end
          end else begin
            _EVAL_820 <= 2'h0;
          end
        end else if (_EVAL_2567) begin
          if (!(_EVAL_169)) begin
            if (_EVAL_1796) begin
              _EVAL_820 <= 2'h3;
            end else begin
              _EVAL_820 <= 2'h0;
            end
          end
        end
      end else if (_EVAL_2429) begin
        if (_EVAL_2747) begin
          _EVAL_820 <= 2'h3;
        end else begin
          _EVAL_820 <= 2'h0;
        end
      end else if (_EVAL_1117) begin
        if (_EVAL_1083) begin
          if (_EVAL_2567) begin
            if (!(_EVAL_169)) begin
              if (_EVAL_1796) begin
                _EVAL_820 <= 2'h3;
              end else begin
                _EVAL_820 <= 2'h0;
              end
            end
          end
        end else begin
          _EVAL_820 <= 2'h0;
        end
      end else if (_EVAL_2567) begin
        if (!(_EVAL_169)) begin
          if (_EVAL_1796) begin
            _EVAL_820 <= 2'h3;
          end else begin
            _EVAL_820 <= 2'h0;
          end
        end
      end
    end else if (_EVAL_1117) begin
      if (_EVAL_1083) begin
        _EVAL_820 <= _EVAL_3084;
      end else begin
        _EVAL_820 <= 2'h0;
      end
    end else begin
      _EVAL_820 <= _EVAL_3084;
    end
    if (_EVAL_63) begin
      _EVAL_845 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2117) begin
        if (_EVAL_1619) begin
          _EVAL_845 <= _EVAL_1770;
        end
      end
    end
    _EVAL_850 <= _EVAL_2101[29:0];
    if (_EVAL_63) begin
      _EVAL_864 <= 8'h0;
    end
    if (_EVAL_63) begin
      _EVAL_880 <= 32'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1127) begin
        _EVAL_880 <= _EVAL_2913;
      end
    end
    if (_EVAL_63) begin
      _EVAL_891 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1150) begin
        _EVAL_891 <= _EVAL_1159;
      end
    end
    if (_EVAL_63) begin
      _EVAL_908 <= 2'h1;
    end
    if (_EVAL_63) begin
      _EVAL_920 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2117) begin
        if (_EVAL_1619) begin
          _EVAL_920 <= _EVAL_3203;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_924 <= 27'h0;
    end
    if (_EVAL_63) begin
      _EVAL_935 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2117) begin
        if (_EVAL_1619) begin
          _EVAL_935 <= _EVAL_2887;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_975 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1424) begin
        if (_EVAL_1619) begin
          _EVAL_975 <= _EVAL_1331;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_1019 <= 1'h0;
    end
    if (_EVAL_1681) begin
      if (_EVAL_1424) begin
        if (_EVAL_985) begin
          _EVAL_1047 <= _EVAL_2258;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_1080 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2117) begin
        if (_EVAL_1619) begin
          _EVAL_1080 <= _EVAL_1815;
        end
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_1424) begin
        if (_EVAL_1619) begin
          _EVAL_1142 <= _EVAL_1896;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_1172 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_789) begin
        _EVAL_1172 <= _EVAL_2887;
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_1658) begin
        if (_EVAL_985) begin
          _EVAL_1239 <= _EVAL_2258;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_1246 <= 2'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2968) begin
        _EVAL_1246 <= _EVAL_1860;
      end
    end
    if (_EVAL_63) begin
      _EVAL_1267 <= 8'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_368) begin
        if (_EVAL_2848) begin
          _EVAL_1267 <= _EVAL_1088;
        end else begin
          _EVAL_1267 <= 8'h0;
        end
      end else if (_EVAL_2670) begin
        if (_EVAL_802) begin
          _EVAL_1267 <= 8'h0;
        end else if (_EVAL_2567) begin
          if (!(_EVAL_169)) begin
            if (_EVAL_1258) begin
              _EVAL_1267 <= _EVAL_2251;
            end
          end
        end
      end else if (_EVAL_2567) begin
        if (!(_EVAL_169)) begin
          if (_EVAL_1258) begin
            _EVAL_1267 <= _EVAL_2251;
          end
        end
      end
    end else if (_EVAL_2567) begin
      if (!(_EVAL_169)) begin
        if (_EVAL_1258) begin
          _EVAL_1267 <= _EVAL_2251;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_1268 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2117) begin
        if (_EVAL_1619) begin
          _EVAL_1268 <= _EVAL_1303;
        end
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_1475) begin
        _EVAL_1271 <= _EVAL_2258;
      end
    end
    _EVAL_1279 <= _EVAL_2719[29:0];
    if (_EVAL_63) begin
      _EVAL_1318 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_368) begin
        _EVAL_1318 <= _EVAL_267;
      end else if (_EVAL_2567) begin
        if (!(_EVAL_169)) begin
          _EVAL_1318 <= _EVAL_1578;
        end
      end
    end else if (_EVAL_2567) begin
      if (!(_EVAL_169)) begin
        _EVAL_1318 <= _EVAL_1578;
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_3148) begin
        _EVAL_1351 <= _EVAL_176;
      end
    end
    if (_EVAL_63) begin
      _EVAL_1353 <= 1'h0;
    end else begin
      _EVAL_1353 <= _EVAL_258;
    end
    if (_EVAL_1681) begin
      if (_EVAL_1807) begin
        _EVAL_1447 <= _EVAL_2740;
      end else if (_EVAL_2567) begin
        if (_EVAL_169) begin
          if (_EVAL_526) begin
            _EVAL_1447 <= _EVAL_1421;
          end
        end
      end
    end else if (_EVAL_2567) begin
      if (_EVAL_169) begin
        if (_EVAL_526) begin
          _EVAL_1447 <= _EVAL_1421;
        end
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_1658) begin
        if (_EVAL_1619) begin
          _EVAL_1450 <= _EVAL_1862;
        end
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_1658) begin
        if (_EVAL_1619) begin
          _EVAL_1451 <= _EVAL_1896;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_1466 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_559) begin
        _EVAL_1466 <= _EVAL_3136;
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_1706) begin
        _EVAL_1467 <= _EVAL_1050;
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_1706) begin
        _EVAL_1491 <= _EVAL_1026;
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_2695) begin
        if (_EVAL_1619) begin
          _EVAL_1493 <= _EVAL_1195;
        end
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_1424) begin
        if (_EVAL_1619) begin
          _EVAL_1507 <= _EVAL_1862;
        end
      end
    end
    _EVAL_1512 <= _EVAL_2640[1:0];
    if (_EVAL_1681) begin
      if (_EVAL_1658) begin
        if (_EVAL_1619) begin
          _EVAL_1595 <= _EVAL_1195;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_1608 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1658) begin
        if (_EVAL_1619) begin
          _EVAL_1608 <= _EVAL_2887;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_1722 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_368) begin
        _EVAL_1722 <= _EVAL_1348;
      end else if (_EVAL_2670) begin
        if (_EVAL_802) begin
          _EVAL_1722 <= 1'h0;
        end else if (_EVAL_3065) begin
          _EVAL_1722 <= 1'h0;
        end else if (_EVAL_2359) begin
          _EVAL_1722 <= _EVAL_1322;
        end
      end else if (_EVAL_3065) begin
        _EVAL_1722 <= 1'h0;
      end else if (_EVAL_2359) begin
        _EVAL_1722 <= _EVAL_1322;
      end
    end else if (_EVAL_3065) begin
      _EVAL_1722 <= 1'h0;
    end else if (_EVAL_2359) begin
      _EVAL_1722 <= _EVAL_1322;
    end
    if (_EVAL_1681) begin
      if (_EVAL_2117) begin
        if (_EVAL_1619) begin
          _EVAL_1755 <= _EVAL_1862;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_1850 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1658) begin
        if (_EVAL_1619) begin
          _EVAL_1850 <= _EVAL_313;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_1888 <= 3'h0;
    end
    if (_EVAL_63) begin
      _EVAL_1948 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_368) begin
        if (_EVAL_2848) begin
          _EVAL_1948 <= _EVAL_3228;
        end else if (_EVAL_2429) begin
          _EVAL_1948 <= _EVAL_1869;
        end else if (_EVAL_1117) begin
          if (_EVAL_1083) begin
            if (_EVAL_2567) begin
              if (!(_EVAL_169)) begin
                _EVAL_1948 <= _EVAL_2927;
              end
            end
          end else begin
            _EVAL_1948 <= 1'h1;
          end
        end else if (_EVAL_2567) begin
          if (!(_EVAL_169)) begin
            _EVAL_1948 <= _EVAL_2927;
          end
        end
      end else if (_EVAL_2429) begin
        _EVAL_1948 <= _EVAL_1869;
      end else if (_EVAL_1117) begin
        if (_EVAL_1083) begin
          if (_EVAL_2567) begin
            if (!(_EVAL_169)) begin
              _EVAL_1948 <= _EVAL_2927;
            end
          end
        end else begin
          _EVAL_1948 <= 1'h1;
        end
      end else if (_EVAL_2567) begin
        if (!(_EVAL_169)) begin
          _EVAL_1948 <= _EVAL_2927;
        end
      end
    end else if (_EVAL_1117) begin
      if (_EVAL_1083) begin
        _EVAL_1948 <= _EVAL_1825;
      end else begin
        _EVAL_1948 <= 1'h1;
      end
    end else begin
      _EVAL_1948 <= _EVAL_1825;
    end
    if (_EVAL_1681) begin
      if (_EVAL_841) begin
        _EVAL_1969 <= _EVAL_152;
      end else if (_EVAL_1294) begin
        _EVAL_1969 <= _EVAL_553;
      end else if (_EVAL_242) begin
        _EVAL_1969 <= _EVAL_916;
      end
    end else if (_EVAL_242) begin
      _EVAL_1969 <= _EVAL_916;
    end
    if (_EVAL_63) begin
      _EVAL_2083 <= 1'h0;
    end
    if (_EVAL_63) begin
      _EVAL_2129 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1706) begin
        _EVAL_2129 <= _EVAL_2487;
      end
    end
    if (_EVAL_63) begin
      _EVAL_2147 <= 2'h3;
    end else if (_EVAL_2519) begin
      _EVAL_2147 <= 2'h3;
    end else begin
      _EVAL_2147 <= 2'h0;
    end
    if (_EVAL_1790) begin
      _EVAL_2148 <= 1'h0;
    end else begin
      _EVAL_2148 <= _EVAL_3128;
    end
    if (_EVAL_63) begin
      _EVAL_2158 <= 1'h0;
    end
    if (_EVAL_63) begin
      _EVAL_2251 <= 8'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_3210) begin
        if (_EVAL_1966) begin
          _EVAL_2251 <= _EVAL_108;
        end else if (_EVAL_1117) begin
          if (_EVAL_1083) begin
            if (_EVAL_2567) begin
              if (!(_EVAL_169)) begin
                if (_EVAL_1258) begin
                  _EVAL_2251 <= _EVAL_108;
                end
              end
            end
          end else if (_EVAL_2848) begin
            _EVAL_2251 <= _EVAL_1267;
          end else if (_EVAL_2567) begin
            if (!(_EVAL_169)) begin
              if (_EVAL_1258) begin
                _EVAL_2251 <= _EVAL_108;
              end
            end
          end
        end else if (_EVAL_2567) begin
          if (!(_EVAL_169)) begin
            if (_EVAL_1258) begin
              _EVAL_2251 <= _EVAL_108;
            end
          end
        end
      end else if (_EVAL_1117) begin
        if (_EVAL_1083) begin
          if (_EVAL_2567) begin
            if (!(_EVAL_169)) begin
              if (_EVAL_1258) begin
                _EVAL_2251 <= _EVAL_108;
              end
            end
          end
        end else if (_EVAL_2848) begin
          _EVAL_2251 <= _EVAL_1267;
        end else begin
          _EVAL_2251 <= _EVAL_674;
        end
      end else begin
        _EVAL_2251 <= _EVAL_674;
      end
    end else if (_EVAL_1117) begin
      if (_EVAL_1083) begin
        _EVAL_2251 <= _EVAL_674;
      end else if (_EVAL_2848) begin
        _EVAL_2251 <= _EVAL_1267;
      end else begin
        _EVAL_2251 <= _EVAL_674;
      end
    end else begin
      _EVAL_2251 <= _EVAL_674;
    end
    if (_EVAL_63) begin
      _EVAL_2268 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2695) begin
        if (_EVAL_1619) begin
          _EVAL_2268 <= _EVAL_2887;
        end
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_2117) begin
        if (_EVAL_985) begin
          _EVAL_2306 <= _EVAL_2258;
        end
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_1150) begin
        _EVAL_2349 <= _EVAL_2837;
      end
    end
    if (_EVAL_63) begin
      _EVAL_2355 <= 3'h0;
    end else if (_EVAL_2567) begin
      if (_EVAL_169) begin
        if (_EVAL_526) begin
          if (_EVAL_2148) begin
            _EVAL_2355 <= 3'h4;
          end else begin
            _EVAL_2355 <= {{1'd0}, _EVAL_2814};
          end
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_2356 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_789) begin
        _EVAL_2356 <= _EVAL_439;
      end
    end
    if (_EVAL_63) begin
      _EVAL_2375 <= 1'h0;
    end
    if (_EVAL_63) begin
      _EVAL_2380 <= 1'h0;
    end else if (_EVAL_2305) begin
      _EVAL_2380 <= 1'h0;
    end else if (_EVAL_1107) begin
      _EVAL_2380 <= 1'h0;
    end else begin
      _EVAL_2380 <= _EVAL_3236;
    end
    if (_EVAL_63) begin
      _EVAL_2387 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_789) begin
        _EVAL_2387 <= _EVAL_437;
      end
    end
    if (_EVAL_63) begin
      _EVAL_2392 <= 2'h0;
    end
    if (_EVAL_63) begin
      _EVAL_2406 <= 1'h0;
    end else begin
      _EVAL_2406 <= _EVAL_3133;
    end
    if (_EVAL_1681) begin
      if (_EVAL_2695) begin
        if (_EVAL_1619) begin
          _EVAL_2445 <= _EVAL_1896;
        end
      end
    end
    if (_EVAL_1452) begin
      _EVAL_2471 <= _EVAL_820;
    end else begin
      _EVAL_2471 <= _EVAL_2147;
    end
    if (_EVAL_63) begin
      _EVAL_2479 <= 10'h0;
    end else begin
      _EVAL_2479 <= _EVAL_1803[9:0];
    end
    if (_EVAL_63) begin
      _EVAL_2486 <= 1'h0;
    end
    if (_EVAL_63) begin
      _EVAL_2542 <= 1'h0;
    end
    if (_EVAL_63) begin
      _EVAL_2579 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2695) begin
        if (_EVAL_1619) begin
          _EVAL_2579 <= _EVAL_1303;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_2593 <= 1'h0;
    end
    if (_EVAL_63) begin
      _EVAL_2609 <= 2'h3;
    end else if (_EVAL_1681) begin
      if (_EVAL_789) begin
        if (_EVAL_817) begin
          _EVAL_2609 <= 2'h3;
        end else begin
          _EVAL_2609 <= 2'h0;
        end
      end else if (_EVAL_2567) begin
        if (_EVAL_169) begin
          if (_EVAL_526) begin
            _EVAL_2609 <= _EVAL_1887;
          end
        end
      end
    end else if (_EVAL_2567) begin
      if (_EVAL_169) begin
        if (_EVAL_526) begin
          _EVAL_2609 <= _EVAL_1887;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_2644 <= 6'h0;
    end else begin
      _EVAL_2644 <= _EVAL_2956[5:0];
    end
    if (_EVAL_63) begin
      _EVAL_2647 <= 1'h0;
    end else if (_EVAL_1117) begin
      if (_EVAL_1083) begin
        _EVAL_2647 <= 1'h0;
      end else if (_EVAL_2567) begin
        if (_EVAL_169) begin
          _EVAL_2647 <= _EVAL_927;
        end
      end
    end else if (_EVAL_2567) begin
      if (_EVAL_169) begin
        _EVAL_2647 <= _EVAL_927;
      end
    end
    if (_EVAL_63) begin
      _EVAL_2654 <= 1'h0;
    end
    if (_EVAL_63) begin
      _EVAL_2665 <= 24'h0;
    end
    if (_EVAL_63) begin
      _EVAL_2673 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2968) begin
        _EVAL_2673 <= _EVAL_1910;
      end
    end
    if (_EVAL_63) begin
      _EVAL_2674 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2695) begin
        if (_EVAL_1619) begin
          _EVAL_2674 <= _EVAL_3203;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_2676 <= 1'h0;
    end
    if (_EVAL_1681) begin
      if (_EVAL_2695) begin
        if (_EVAL_985) begin
          _EVAL_2689 <= _EVAL_2258;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_2708 <= 2'h0;
    end
    if (_EVAL_63) begin
      _EVAL_2732 <= 2'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1706) begin
        _EVAL_2732 <= _EVAL_1051;
      end
    end
    if (_EVAL_63) begin
      _EVAL_2764 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1424) begin
        if (_EVAL_1619) begin
          _EVAL_2764 <= _EVAL_2887;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_2784 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2695) begin
        if (_EVAL_1619) begin
          _EVAL_2784 <= _EVAL_3109;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_2791 <= 2'h0;
    end
    _EVAL_2799 <= _EVAL_715[29:0];
    _EVAL_2828 <= _EVAL_2942[15:0];
    if (_EVAL_63) begin
      _EVAL_2842 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2695) begin
        if (_EVAL_1619) begin
          _EVAL_2842 <= _EVAL_811;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_2844 <= 1'h0;
    end
    _EVAL_2870 <= _EVAL_2870;
    if (_EVAL_1681) begin
      if (_EVAL_1424) begin
        if (_EVAL_1619) begin
          _EVAL_2907 <= _EVAL_1195;
        end
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_2117) begin
        if (_EVAL_1619) begin
          _EVAL_2914 <= _EVAL_1896;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_2927 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2429) begin
        _EVAL_2927 <= _EVAL_3027;
      end else if (_EVAL_1117) begin
        if (_EVAL_1083) begin
          if (_EVAL_2567) begin
            _EVAL_2927 <= _EVAL_1427;
          end
        end else begin
          _EVAL_2927 <= _EVAL_1948;
        end
      end else if (_EVAL_2567) begin
        _EVAL_2927 <= _EVAL_1427;
      end
    end else if (_EVAL_1117) begin
      if (_EVAL_1083) begin
        if (_EVAL_2567) begin
          _EVAL_2927 <= _EVAL_1427;
        end
      end else begin
        _EVAL_2927 <= _EVAL_1948;
      end
    end else if (_EVAL_2567) begin
      _EVAL_2927 <= _EVAL_1427;
    end
    if (_EVAL_1681) begin
      if (_EVAL_2002) begin
        _EVAL_2931 <= _EVAL_2258;
      end else if (_EVAL_2567) begin
        if (!(_EVAL_169)) begin
          _EVAL_2931 <= _EVAL_109;
        end
      end
    end else if (_EVAL_2567) begin
      if (!(_EVAL_169)) begin
        _EVAL_2931 <= _EVAL_109;
      end
    end
    if (_EVAL_63) begin
      _EVAL_2987 <= 2'h0;
    end
    if (_EVAL_63) begin
      _EVAL_3052 <= 1'h0;
    end else begin
      _EVAL_3052 <= _EVAL_2843[0];
    end
    if (_EVAL_63) begin
      _EVAL_3058 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1424) begin
        if (_EVAL_1619) begin
          _EVAL_3058 <= _EVAL_2208;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_3068 <= 2'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_559) begin
        _EVAL_3068 <= _EVAL_1676;
      end
    end
    _EVAL_3070 <= _EVAL_2037[5:0];
    if (_EVAL_63) begin
      _EVAL_3115 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_2695) begin
        if (_EVAL_1619) begin
          _EVAL_3115 <= _EVAL_1236;
        end
      end
    end
    if (_EVAL_63) begin
      _EVAL_3143 <= 1'h0;
    end
    if (_EVAL_63) begin
      _EVAL_3152 <= 31'h40901105;
    end
    if (_EVAL_63) begin
      _EVAL_3170 <= 2'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1150) begin
        _EVAL_3170 <= _EVAL_875;
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_1706) begin
        _EVAL_3183 <= _EVAL_2725;
      end
    end
    if (_EVAL_49) begin
      _EVAL_3184 <= _EVAL_30;
    end
    if (_EVAL_63) begin
      _EVAL_3195 <= 2'h0;
    end
    if (_EVAL_63) begin
      _EVAL_3213 <= 1'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1424) begin
        if (_EVAL_1619) begin
          _EVAL_3213 <= _EVAL_1303;
        end
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_2695) begin
        if (_EVAL_1619) begin
          _EVAL_3217 <= _EVAL_1862;
        end
      end
    end
    if (_EVAL_49) begin
      _EVAL_3231 <= _EVAL_1;
    end
    if (_EVAL_63) begin
      _EVAL_3239 <= 58'h0;
    end else if (_EVAL_1681) begin
      if (_EVAL_1878) begin
        _EVAL_3239 <= _EVAL_2705;
      end else if (_EVAL_2501) begin
        _EVAL_3239 <= _EVAL_282;
      end else if (_EVAL_1148) begin
        _EVAL_3239 <= _EVAL_2918;
      end
    end else if (_EVAL_1148) begin
      _EVAL_3239 <= _EVAL_2918;
    end
    if (_EVAL_1681) begin
      if (_EVAL_2968) begin
        _EVAL_3242 <= _EVAL_1302;
      end
    end
    if (_EVAL_63) begin
      _EVAL_3256 <= 6'h0;
    end else begin
      _EVAL_3256 <= _EVAL_1901[5:0];
    end
  end
endmodule
