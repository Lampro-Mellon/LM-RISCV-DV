//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_61(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  output        _EVAL_1,
  input  [31:0] _EVAL_2,
  output        _EVAL_3,
  input  [31:0] _EVAL_4,
  output [31:0] _EVAL_5,
  input  [29:0] _EVAL_6,
  input  [3:0]  _EVAL_7,
  output        _EVAL_8,
  output        _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  output        _EVAL_12,
  output        _EVAL_13,
  input         _EVAL_14,
  output [2:0]  _EVAL_15,
  input         _EVAL_16,
  input  [2:0]  _EVAL_17,
  output [1:0]  _EVAL_18,
  input         _EVAL_19,
  input         _EVAL_20,
  output        _EVAL_21,
  input  [2:0]  _EVAL_22,
  output [3:0]  _EVAL_23,
  output        _EVAL_24,
  input         _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  output [2:0]  _EVAL_30,
  output [29:0] _EVAL_31,
  output [2:0]  _EVAL_32,
  output [2:0]  _EVAL_33,
  output        _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  input  [3:0]  _EVAL_38,
  input         _EVAL_39,
  input         _EVAL_40,
  output [3:0]  _EVAL_41,
  input  [3:0]  _EVAL_42,
  output        _EVAL_43,
  output [3:0]  _EVAL_44,
  output [2:0]  _EVAL_45,
  output        _EVAL_46,
  input  [2:0]  _EVAL_47,
  input  [2:0]  _EVAL_48,
  output [31:0] _EVAL_49,
  output        _EVAL_50,
  output        _EVAL_51,
  output        _EVAL_52,
  output        _EVAL_53,
  input  [1:0]  _EVAL_54
);
  assign _EVAL_12 = _EVAL_37;
  assign _EVAL_50 = _EVAL_16;
  assign _EVAL_3 = _EVAL_27;
  assign _EVAL_51 = _EVAL_20;
  assign _EVAL_52 = _EVAL_10;
  assign _EVAL_9 = _EVAL_14;
  assign _EVAL_31 = _EVAL_6;
  assign _EVAL_24 = _EVAL_26;
  assign _EVAL_5 = _EVAL_4;
  assign _EVAL_15 = _EVAL_48;
  assign _EVAL_45 = _EVAL_17;
  assign _EVAL_30 = _EVAL;
  assign _EVAL_32 = _EVAL_22;
  assign _EVAL_13 = _EVAL_0;
  assign _EVAL_23 = _EVAL_42;
  assign _EVAL_46 = _EVAL_39;
  assign _EVAL_44 = _EVAL_38;
  assign _EVAL_33 = _EVAL_47;
  assign _EVAL_53 = _EVAL_36;
  assign _EVAL_41 = _EVAL_7;
  assign _EVAL_34 = _EVAL_40;
  assign _EVAL_8 = _EVAL_29;
  assign _EVAL_49 = _EVAL_2;
  assign _EVAL_1 = _EVAL_25;
  assign _EVAL_18 = _EVAL_54;
  assign _EVAL_21 = _EVAL_19;
  assign _EVAL_43 = _EVAL_35;
endmodule
