//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_8(
  output [2:0]  _EVAL,
  input  [1:0]  _EVAL_0,
  input         _EVAL_1,
  output [2:0]  _EVAL_2,
  input         _EVAL_3,
  output        _EVAL_4,
  output        _EVAL_5,
  input         _EVAL_6,
  input  [1:0]  _EVAL_7,
  output        _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  output [2:0]  _EVAL_11,
  input  [3:0]  _EVAL_12,
  output        _EVAL_13,
  input  [2:0]  _EVAL_14,
  output        _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  output [3:0]  _EVAL_18,
  output [3:0]  _EVAL_19,
  input         _EVAL_20,
  input         _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  output        _EVAL_24,
  output [31:0] _EVAL_25,
  input         _EVAL_26,
  output        _EVAL_27,
  output        _EVAL_28,
  output        _EVAL_29,
  input         _EVAL_30,
  output        _EVAL_31,
  input         _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_34,
  output        _EVAL_35,
  input  [31:0] _EVAL_36,
  output        _EVAL_37,
  input         _EVAL_38,
  output        _EVAL_39,
  input         _EVAL_40,
  output        _EVAL_41,
  output [2:0]  _EVAL_42,
  output        _EVAL_43,
  output        _EVAL_44,
  output [31:0] _EVAL_45,
  output [2:0]  _EVAL_46,
  input  [31:0] _EVAL_47,
  input  [2:0]  _EVAL_48,
  input         _EVAL_49,
  input  [31:0] _EVAL_50,
  input         _EVAL_51,
  output [31:0] _EVAL_52,
  output        _EVAL_53,
  output        _EVAL_54,
  output [31:0] _EVAL_55,
  input  [3:0]  _EVAL_56,
  input  [2:0]  _EVAL_57,
  input  [2:0]  _EVAL_58,
  output [3:0]  _EVAL_59,
  output        _EVAL_60,
  output [3:0]  _EVAL_61,
  input         _EVAL_62,
  output [1:0]  _EVAL_63,
  output [3:0]  _EVAL_64,
  output [3:0]  _EVAL_65,
  input         _EVAL_66,
  output [31:0] _EVAL_67,
  input         _EVAL_68,
  input         _EVAL_69,
  input         _EVAL_70,
  input         _EVAL_71,
  input         _EVAL_72,
  output        _EVAL_73,
  input         _EVAL_74,
  input         _EVAL_75,
  input         _EVAL_76,
  output        _EVAL_77,
  output        _EVAL_78,
  output        _EVAL_79,
  output [31:0] _EVAL_80,
  output        _EVAL_81,
  output        _EVAL_82,
  output        _EVAL_83,
  output [2:0]  _EVAL_84,
  output        _EVAL_85,
  input  [3:0]  _EVAL_86,
  input  [3:0]  _EVAL_87,
  output        _EVAL_88,
  output        _EVAL_89,
  input         _EVAL_90,
  output        _EVAL_91,
  output        _EVAL_92,
  output        _EVAL_93,
  input  [3:0]  _EVAL_94,
  output        _EVAL_95,
  input         _EVAL_96,
  input  [3:0]  _EVAL_97,
  input         _EVAL_98,
  input  [31:0] _EVAL_99,
  input  [2:0]  _EVAL_100,
  input  [31:0] _EVAL_101,
  output        _EVAL_102,
  input         _EVAL_103,
  input  [2:0]  _EVAL_104,
  input  [31:0] _EVAL_105,
  input         _EVAL_106,
  output [1:0]  _EVAL_107,
  input         _EVAL_108
);
  wire [5:0] _EVAL_111;
  wire [32:0] _EVAL_112;
  wire [7:0] _EVAL_114;
  wire [32:0] _EVAL_116;
  wire [32:0] _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_124;
  wire [22:0] _EVAL_126;
  wire  _EVAL_127;
  wire [32:0] _EVAL_128;
  wire  _EVAL_130;
  wire  _EVAL_135;
  wire  _EVAL_137;
  wire [32:0] _EVAL_143;
  wire [32:0] _EVAL_144;
  wire [1:0] _EVAL_149;
  wire [32:0] _EVAL_150;
  wire  _EVAL_151;
  wire [1:0] _EVAL_155;
  wire  _EVAL_157;
  wire [5:0] _EVAL_160;
  wire [32:0] _EVAL_164;
  wire  _EVAL_165;
  wire [5:0] _EVAL_166;
  wire [7:0] _EVAL_173;
  wire [22:0] _EVAL_174;
  wire [6:0] _EVAL_176;
  wire [31:0] _EVAL_177;
  wire [6:0] _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_184;
  wire  _EVAL_187;
  wire  _EVAL_188;
  reg  _EVAL_191;
  reg [31:0] _RAND_0;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_200;
  wire  _EVAL_203;
  wire [31:0] _EVAL_207;
  reg  _EVAL_208;
  reg [31:0] _RAND_1;
  wire [32:0] _EVAL_209;
  reg [1:0] _EVAL_212;
  reg [31:0] _RAND_2;
  wire [1:0] _EVAL_216;
  wire  _EVAL_218;
  wire  _EVAL_220;
  reg [5:0] _EVAL_224;
  reg [31:0] _RAND_3;
  wire  _EVAL_225;
  wire [7:0] _EVAL_227;
  wire  _EVAL_228;
  wire [5:0] _EVAL_236;
  wire  _EVAL_241;
  wire  _EVAL_245;
  reg [5:0] _EVAL_246;
  reg [31:0] _RAND_4;
  wire  _EVAL_247;
  wire [7:0] _EVAL_249;
  assign _EVAL_13 = _EVAL_76;
  assign _EVAL_53 = _EVAL_9;
  assign _EVAL_165 = ~_EVAL_187;
  assign _EVAL_59 = _EVAL_86;
  assign _EVAL_15 = _EVAL_66;
  assign _EVAL_84 = _EVAL_100;
  assign _EVAL_35 = _EVAL_108;
  assign _EVAL_102 = _EVAL_96;
  assign _EVAL_19 = _EVAL_12;
  assign _EVAL_184 = $signed(_EVAL_164) == 33'sh0;
  assign _EVAL_31 = _EVAL_51;
  assign _EVAL_236 = _EVAL_227[7:2];
  assign _EVAL_112 = {1'b0,$signed(_EVAL_207)};
  assign _EVAL_126 = 23'hff << _EVAL_97;
  assign _EVAL_4 = _EVAL_17;
  assign _EVAL_93 = _EVAL_34;
  assign _EVAL_194 = _EVAL_191 | _EVAL_208;
  assign _EVAL_89 = _EVAL_70;
  assign _EVAL_2 = _EVAL_14;
  assign _EVAL_46 = _EVAL_57;
  assign _EVAL_55 = _EVAL_50;
  assign _EVAL_166 = _EVAL_180[5:0];
  assign _EVAL_54 = _EVAL_3;
  assign _EVAL_67 = _EVAL_101;
  assign _EVAL_228 = $signed(_EVAL_150) == 33'sh0;
  assign _EVAL_77 = _EVAL_74;
  assign _EVAL_91 = _EVAL_69;
  assign _EVAL_95 = _EVAL_16;
  assign _EVAL_151 = _EVAL_49 & _EVAL_195;
  assign _EVAL_195 = _EVAL_228 | _EVAL_165;
  assign _EVAL_207 = _EVAL_50 ^ 32'h80000000;
  assign _EVAL_116 = {1'b0,$signed(_EVAL_50)};
  assign _EVAL_160 = _EVAL_176[5:0];
  assign _EVAL_81 = _EVAL_6;
  assign _EVAL_188 = _EVAL_220 & _EVAL_245;
  assign _EVAL_43 = _EVAL_75;
  assign _EVAL_176 = _EVAL_246 - 6'h1;
  assign _EVAL_181 = _EVAL_246 == 6'h0;
  assign _EVAL_45 = _EVAL_36;
  assign _EVAL_73 = _EVAL_49 & _EVAL_195;
  assign _EVAL_28 = _EVAL_21;
  assign _EVAL_245 = _EVAL_30 & _EVAL_62;
  assign _EVAL_157 = ~_EVAL_121;
  assign _EVAL_11 = _EVAL_48;
  assign _EVAL_39 = _EVAL_38;
  assign _EVAL_218 = _EVAL_124 & _EVAL_247;
  assign _EVAL_79 = _EVAL_33;
  assign _EVAL_227 = ~_EVAL_114;
  assign _EVAL_209 = $signed(_EVAL_112) & 33'sh80000000;
  assign _EVAL_196 = _EVAL_104 != 3'h6;
  assign _EVAL_174 = 23'hff << _EVAL_12;
  assign _EVAL_249 = ~_EVAL_173;
  assign _EVAL_52 = _EVAL_105;
  assign _EVAL_27 = _EVAL_72;
  assign _EVAL_144 = _EVAL_128;
  assign _EVAL_130 = _EVAL_203 | _EVAL_200;
  assign _EVAL_177 = _EVAL_50 ^ 32'h40000000;
  assign _EVAL = _EVAL_58;
  assign _EVAL_150 = _EVAL_209;
  assign _EVAL_149 = _EVAL_216 | _EVAL_155;
  assign _EVAL_225 = $signed(_EVAL_144) == 33'sh0;
  assign _EVAL_216 = {{1'd0}, _EVAL_225};
  assign _EVAL_128 = $signed(_EVAL_143) & 33'sh40000000;
  assign _EVAL_124 = _EVAL_151 & _EVAL_103;
  assign _EVAL_173 = _EVAL_126[7:0];
  assign _EVAL_203 = _EVAL_149 == 2'h0;
  assign _EVAL_164 = _EVAL_120;
  assign _EVAL_187 = _EVAL_241 & _EVAL_130;
  assign _EVAL_92 = _EVAL_22;
  assign _EVAL_137 = _EVAL_104[0];
  assign _EVAL_64 = _EVAL_97;
  assign _EVAL_220 = _EVAL_135 & _EVAL_196;
  assign _EVAL_111 = _EVAL_249[7:2];
  assign _EVAL_200 = _EVAL_212 != _EVAL_149;
  assign _EVAL_155 = _EVAL_184 ? 2'h2 : 2'h0;
  assign _EVAL_44 = _EVAL_10;
  assign _EVAL_121 = _EVAL_57[2];
  assign _EVAL_82 = _EVAL_71;
  assign _EVAL_180 = _EVAL_224 - 6'h1;
  assign _EVAL_25 = _EVAL_47;
  assign _EVAL_127 = _EVAL_181 & _EVAL_124;
  assign _EVAL_247 = ~_EVAL_228;
  assign _EVAL_80 = _EVAL_99;
  assign _EVAL_241 = _EVAL_181 & _EVAL_194;
  assign _EVAL_85 = _EVAL_40;
  assign _EVAL_65 = _EVAL_56;
  assign _EVAL_42 = _EVAL_104;
  assign _EVAL_8 = _EVAL_103 & _EVAL_195;
  assign _EVAL_88 = _EVAL_98;
  assign _EVAL_24 = _EVAL_90;
  assign _EVAL_135 = _EVAL_224 == 6'h0;
  assign _EVAL_41 = _EVAL_26;
  assign _EVAL_120 = $signed(_EVAL_116) & 33'sh40000000;
  assign _EVAL_61 = _EVAL_94;
  assign _EVAL_29 = _EVAL_106;
  assign _EVAL_18 = _EVAL_87;
  assign _EVAL_37 = _EVAL_23;
  assign _EVAL_83 = _EVAL_32;
  assign _EVAL_114 = _EVAL_174[7:0];
  assign _EVAL_143 = {1'b0,$signed(_EVAL_177)};
  assign _EVAL_60 = _EVAL_62;
  assign _EVAL_5 = _EVAL_20;
  assign _EVAL_63 = _EVAL_0;
  assign _EVAL_78 = _EVAL_30;
  assign _EVAL_107 = _EVAL_7;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_191 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_208 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_212 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_224 = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_246 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_68) begin
    if (_EVAL_1) begin
      _EVAL_191 <= 1'h0;
    end else if (_EVAL_188) begin
      if (~_EVAL_66) begin
        _EVAL_191 <= 1'h0;
      end else if (_EVAL_127) begin
        if (~_EVAL_16) begin
          _EVAL_191 <= _EVAL_247;
        end
      end
    end else if (_EVAL_127) begin
      if (~_EVAL_16) begin
        _EVAL_191 <= _EVAL_247;
      end
    end
    if (_EVAL_1) begin
      _EVAL_208 <= 1'h0;
    end else if (_EVAL_188) begin
      if (_EVAL_66) begin
        _EVAL_208 <= 1'h0;
      end else if (_EVAL_127) begin
        if (_EVAL_16) begin
          _EVAL_208 <= _EVAL_247;
        end
      end
    end else if (_EVAL_127) begin
      if (_EVAL_16) begin
        _EVAL_208 <= _EVAL_247;
      end
    end
    if (_EVAL_218) begin
      _EVAL_212 <= _EVAL_149;
    end
    if (_EVAL_1) begin
      _EVAL_224 <= 6'h0;
    end else if (_EVAL_245) begin
      if (_EVAL_135) begin
        if (_EVAL_137) begin
          _EVAL_224 <= _EVAL_111;
        end else begin
          _EVAL_224 <= 6'h0;
        end
      end else begin
        _EVAL_224 <= _EVAL_166;
      end
    end
    if (_EVAL_1) begin
      _EVAL_246 <= 6'h0;
    end else if (_EVAL_124) begin
      if (_EVAL_181) begin
        if (_EVAL_157) begin
          _EVAL_246 <= _EVAL_236;
        end else begin
          _EVAL_246 <= 6'h0;
        end
      end else begin
        _EVAL_246 <= _EVAL_160;
      end
    end
  end
endmodule
