//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_64_assert(
  input  [2:0]  _EVAL,
  input  [2:0]  _EVAL_0,
  input  [3:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [3:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [1:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [2:0]  _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input  [2:0]  _EVAL_16,
  input  [29:0] _EVAL_17,
  input  [3:0]  _EVAL_18
);
  wire  _EVAL_19;
  wire [22:0] _EVAL_20;
  wire  _EVAL_21;
  wire [6:0] _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire [3:0] _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire [4:0] _EVAL_29;
  wire [29:0] _EVAL_30;
  wire [5:0] _EVAL_31;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire [30:0] _EVAL_46;
  wire  _EVAL_47;
  wire [31:0] plusarg_reader_out;
  wire [29:0] _EVAL_49;
  wire [22:0] _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire [6:0] _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire [29:0] _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire [7:0] _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire [30:0] _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire [4:0] _EVAL_78;
  wire [7:0] _EVAL_79;
  wire  _EVAL_80;
  wire [30:0] _EVAL_81;
  wire  _EVAL_82;
  reg [3:0] _EVAL_83;
  reg [31:0] _RAND_0;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire [6:0] _EVAL_87;
  wire [4:0] _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire [30:0] _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire [1:0] _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire [1:0] _EVAL_98;
  reg [3:0] _EVAL_99;
  reg [31:0] _RAND_1;
  wire [32:0] _EVAL_100;
  wire  _EVAL_101;
  reg [5:0] _EVAL_102;
  reg [31:0] _RAND_2;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  reg [2:0] _EVAL_106;
  reg [31:0] _RAND_3;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire [3:0] _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  reg [5:0] _EVAL_121;
  reg [31:0] _RAND_4;
  wire  _EVAL_122;
  wire [5:0] _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  reg [4:0] _EVAL_127;
  reg [31:0] _RAND_5;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_143;
  wire [6:0] _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire [30:0] _EVAL_152;
  wire [7:0] _EVAL_153;
  wire  _EVAL_154;
  reg [31:0] _EVAL_155;
  reg [31:0] _RAND_6;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire [1:0] _EVAL_170;
  wire  _EVAL_171;
  wire [30:0] _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire [29:0] _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire [4:0] _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire [4:0] _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire [7:0] _EVAL_202;
  reg [2:0] _EVAL_203;
  reg [31:0] _RAND_7;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire [4:0] _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  reg [5:0] _EVAL_213;
  reg [31:0] _RAND_8;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire [30:0] _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire [5:0] _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_239;
  wire [5:0] _EVAL_240;
  wire  _EVAL_241;
  wire [4:0] _EVAL_242;
  wire [29:0] _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire [30:0] _EVAL_250;
  wire  _EVAL_251;
  wire [30:0] _EVAL_252;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire [1:0] _EVAL_256;
  wire  _EVAL_257;
  reg [5:0] _EVAL_258;
  reg [31:0] _RAND_9;
  wire [7:0] _EVAL_259;
  wire  _EVAL_260;
  wire [7:0] _EVAL_261;
  wire [7:0] _EVAL_262;
  wire [7:0] _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire [3:0] _EVAL_266;
  wire  _EVAL_267;
  wire [31:0] _EVAL_268;
  wire  _EVAL_269;
  reg [2:0] _EVAL_270;
  reg [31:0] _RAND_10;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire [5:0] _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  reg [2:0] _EVAL_281;
  reg [31:0] _RAND_11;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  reg [2:0] _EVAL_285;
  reg [31:0] _RAND_12;
  reg [1:0] _EVAL_286;
  reg [31:0] _RAND_13;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire [5:0] _EVAL_289;
  wire  _EVAL_290;
  wire [4:0] _EVAL_291;
  wire [30:0] _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  reg  _EVAL_301;
  reg [31:0] _RAND_14;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire [30:0] _EVAL_308;
  reg  _EVAL_309;
  reg [31:0] _RAND_15;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire [3:0] _EVAL_312;
  reg [29:0] _EVAL_313;
  reg [31:0] _RAND_16;
  wire  _EVAL_314;
  wire [30:0] _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire  _EVAL_321;
  wire  _EVAL_323;
  wire  _EVAL_324;
  wire  _EVAL_325;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_308 = {1'b0,$signed(_EVAL_59)};
  assign _EVAL_36 = _EVAL_11 & _EVAL_149;
  assign _EVAL_277 = _EVAL_214 | _EVAL_15;
  assign _EVAL_19 = ~_EVAL_269;
  assign _EVAL_67 = _EVAL_169 | _EVAL_15;
  assign _EVAL_239 = ~_EVAL_41;
  assign _EVAL_119 = _EVAL_188 | _EVAL_15;
  assign _EVAL_30 = _EVAL_17 ^ 30'h2000000;
  assign _EVAL_266 = {_EVAL_321,_EVAL_201,_EVAL_249,_EVAL_186};
  assign _EVAL_124 = ~_EVAL_217;
  assign _EVAL_54 = _EVAL_260 | _EVAL_15;
  assign _EVAL_134 = _EVAL_11 & _EVAL_133;
  assign _EVAL_171 = ~_EVAL_60;
  assign _EVAL_245 = $signed(_EVAL_91) == 31'sh0;
  assign _EVAL_90 = ~_EVAL_193;
  assign _EVAL_82 = _EVAL_241 & _EVAL_131;
  assign _EVAL_85 = _EVAL_257 | _EVAL_15;
  assign _EVAL_193 = _EVAL_77 | _EVAL_15;
  assign _EVAL_175 = _EVAL_11 & _EVAL_57;
  assign _EVAL_125 = _EVAL_310 | _EVAL_15;
  assign _EVAL_79 = ~_EVAL_66;
  assign _EVAL_173 = ~_EVAL_86;
  assign _EVAL_25 = _EVAL_3 & _EVAL_118;
  assign _EVAL_72 = _EVAL_248 | _EVAL_23;
  assign _EVAL_20 = 23'hff << _EVAL_18;
  assign _EVAL_182 = ~_EVAL_73;
  assign _EVAL_236 = _EVAL_79[7:2];
  assign _EVAL_144 = _EVAL_121 - 6'h1;
  assign _EVAL_27 = _EVAL_18 >= 4'h2;
  assign _EVAL_292 = $signed(_EVAL_252) & -31'sh5000;
  assign _EVAL_55 = $signed(_EVAL_250) == 31'sh0;
  assign _EVAL_88 = _EVAL_153[4:0];
  assign _EVAL_40 = _EVAL_1 >= 4'h2;
  assign _EVAL_101 = ~_EVAL_158;
  assign _EVAL_28 = ~_EVAL_112;
  assign _EVAL_154 = ~_EVAL_139;
  assign _EVAL_242 = ~_EVAL_199;
  assign _EVAL_259 = _EVAL_111 ? _EVAL_261 : 8'h0;
  assign _EVAL_138 = _EVAL_0 == 3'h1;
  assign _EVAL_299 = _EVAL_165 | _EVAL_15;
  assign _EVAL_269 = _EVAL_221 | _EVAL_15;
  assign _EVAL_255 = _EVAL_5 & _EVAL_180;
  assign _EVAL_307 = _EVAL_258 == 6'h0;
  assign _EVAL_311 = _EVAL_6 == _EVAL_286;
  assign _EVAL_303 = _EVAL_11 & _EVAL_265;
  assign _EVAL_198 = ~_EVAL_85;
  assign _EVAL_157 = _EVAL <= 3'h3;
  assign _EVAL_316 = _EVAL_318 | _EVAL_15;
  assign _EVAL_149 = _EVAL_16 == 3'h6;
  assign _EVAL_306 = _EVAL_17[0];
  assign _EVAL_34 = _EVAL_98 == 2'h1;
  assign _EVAL_211 = _EVAL_70 & _EVAL_84;
  assign _EVAL_261 = 8'h1 << _EVAL_13;
  assign _EVAL_64 = _EVAL_1 <= 4'h8;
  assign _EVAL_248 = _EVAL_204 | _EVAL_245;
  assign _EVAL_179 = _EVAL_192 | _EVAL_15;
  assign _EVAL_52 = _EVAL_16[2];
  assign _EVAL_271 = ~_EVAL_277;
  assign _EVAL_282 = _EVAL_53 | _EVAL_143;
  assign _EVAL_293 = _EVAL_16 == 3'h1;
  assign _EVAL_89 = _EVAL_40 | _EVAL_95;
  assign _EVAL_216 = _EVAL_233 & _EVAL_306;
  assign _EVAL_228 = ~_EVAL_272;
  assign _EVAL_165 = _EVAL_145 | _EVAL_229;
  assign _EVAL_191 = ~_EVAL_247;
  assign _EVAL_272 = _EVAL_24 | _EVAL_15;
  assign _EVAL_279 = _EVAL_0 == 3'h6;
  assign _EVAL_222 = _EVAL_273 | _EVAL_15;
  assign _EVAL_200 = _EVAL_246 | _EVAL_15;
  assign _EVAL_69 = _EVAL_152;
  assign _EVAL_120 = _EVAL_256[0];
  assign _EVAL_204 = $signed(_EVAL_224) == 31'sh0;
  assign _EVAL_109 = _EVAL_11 & _EVAL_323;
  assign _EVAL_315 = $signed(_EVAL_308) & -31'sh1000;
  assign _EVAL_201 = _EVAL_187 | _EVAL_167;
  assign _EVAL_217 = _EVAL_110 | _EVAL_15;
  assign _EVAL_22 = _EVAL_258 - 6'h1;
  assign _EVAL_156 = ~_EVAL_314;
  assign _EVAL_91 = _EVAL_292;
  assign _EVAL_166 = plusarg_reader_out == 32'h0;
  assign _EVAL_188 = _EVAL_312 == 4'h0;
  assign _EVAL_197 = _EVAL_88 != _EVAL_199;
  assign _EVAL_133 = _EVAL_16 == 3'h2;
  assign _EVAL_45 = _EVAL_96 | _EVAL_15;
  assign _EVAL_92 = ~_EVAL_63;
  assign _EVAL_190 = _EVAL_16 == _EVAL_270;
  assign _EVAL_76 = _EVAL_297 | _EVAL_15;
  assign _EVAL_122 = ~_EVAL_254;
  assign _EVAL_128 = _EVAL_16 == 3'h7;
  assign _EVAL_310 = _EVAL_295 | _EVAL_234;
  assign _EVAL_302 = _EVAL_0 == 3'h0;
  assign _EVAL_146 = _EVAL_97 | _EVAL_15;
  assign _EVAL_221 = _EVAL_25 == 4'h0;
  assign _EVAL_70 = _EVAL_7 & _EVAL_11;
  assign _EVAL_94 = 2'h1 << _EVAL_235;
  assign _EVAL_71 = _EVAL_5 & _EVAL_280;
  assign _EVAL_161 = _EVAL_88 != 5'h0;
  assign _EVAL_323 = ~_EVAL_84;
  assign _EVAL_135 = _EVAL_190 | _EVAL_15;
  assign _EVAL_163 = _EVAL_120 & _EVAL_216;
  assign _EVAL_187 = _EVAL_40 | _EVAL_162;
  assign _EVAL_312 = ~_EVAL_3;
  assign _EVAL_162 = _EVAL_195 & _EVAL_233;
  assign _EVAL_80 = ~_EVAL_125;
  assign _EVAL_153 = _EVAL_237 ? _EVAL_202 : 8'h0;
  assign _EVAL_50 = 23'hff << _EVAL_1;
  assign _EVAL_189 = _EVAL_136 & _EVAL_55;
  assign _EVAL_274 = ~_EVAL_126;
  assign _EVAL_51 = _EVAL_282 | _EVAL_15;
  assign _EVAL_260 = _EVAL <= 3'h1;
  assign _EVAL_86 = _EVAL_215 | _EVAL_15;
  assign _EVAL_62 = _EVAL_207 | _EVAL_15;
  assign _EVAL_212 = ~_EVAL_26;
  assign _EVAL_53 = _EVAL_43 | _EVAL_141;
  assign _EVAL_249 = _EVAL_89 | _EVAL_39;
  assign _EVAL_250 = _EVAL_315;
  assign _EVAL_321 = _EVAL_187 | _EVAL_163;
  assign _EVAL_319 = ~_EVAL_146;
  assign _EVAL_178 = _EVAL_0 == 3'h5;
  assign _EVAL_23 = $signed(_EVAL_69) == 31'sh0;
  assign _EVAL_140 = _EVAL_120 & _EVAL_82;
  assign _EVAL_263 = ~_EVAL_262;
  assign _EVAL_247 = _EVAL_181 | _EVAL_15;
  assign _EVAL_174 = _EVAL_16 == 3'h4;
  assign _EVAL_252 = {1'b0,$signed(_EVAL_17)};
  assign _EVAL_233 = _EVAL_17[1];
  assign _EVAL_224 = _EVAL_172;
  assign _EVAL_65 = ~_EVAL_12;
  assign _EVAL_254 = _EVAL_78[0];
  assign _EVAL_192 = _EVAL_6 == 2'h0;
  assign _EVAL_78 = _EVAL_127 >> _EVAL_2;
  assign _EVAL_232 = _EVAL <= 3'h4;
  assign _EVAL_136 = _EVAL_1 <= 4'h2;
  assign _EVAL_251 = ~_EVAL_288;
  assign _EVAL_287 = ~_EVAL_76;
  assign _EVAL_103 = _EVAL_98 == 2'h0;
  assign _EVAL_57 = _EVAL_16 == 3'h0;
  assign _EVAL_275 = _EVAL_87[5:0];
  assign _EVAL_265 = _EVAL_16 == 3'h3;
  assign _EVAL_325 = ~_EVAL_58;
  assign _EVAL_113 = ~_EVAL_15;
  assign _EVAL_63 = _EVAL_189 | _EVAL_15;
  assign _EVAL_320 = _EVAL_0 == 3'h2;
  assign _EVAL_96 = _EVAL == _EVAL_106;
  assign _EVAL_229 = _EVAL_2 == 3'h4;
  assign _EVAL_244 = _EVAL_17 & _EVAL_185;
  assign _EVAL_60 = _EVAL_37 | _EVAL_15;
  assign _EVAL_278 = ~_EVAL_54;
  assign _EVAL_206 = ~_EVAL_179;
  assign _EVAL_264 = _EVAL_14 & _EVAL_5;
  assign _EVAL_118 = ~_EVAL_266;
  assign _EVAL_164 = _EVAL_10 == _EVAL_309;
  assign _EVAL_304 = ~_EVAL_21;
  assign _EVAL_46 = {1'b0,$signed(_EVAL_49)};
  assign _EVAL_87 = _EVAL_213 - 6'h1;
  assign _EVAL_231 = _EVAL_5 & _EVAL_279;
  assign _EVAL_215 = _EVAL_0 <= 3'h6;
  assign _EVAL_273 = ~_EVAL_4;
  assign _EVAL_220 = _EVAL_210 | _EVAL_284;
  assign _EVAL_129 = ~_EVAL_116;
  assign _EVAL_68 = ~_EVAL_51;
  assign _EVAL_305 = _EVAL_244 == 30'h0;
  assign _EVAL_172 = $signed(_EVAL_81) & -31'sh1000000;
  assign _EVAL_283 = ~_EVAL_105;
  assign _EVAL_317 = _EVAL_44 | _EVAL_15;
  assign _EVAL_74 = ~_EVAL_316;
  assign _EVAL_288 = _EVAL_127 != 5'h0;
  assign _EVAL_226 = ~_EVAL_119;
  assign _EVAL_110 = _EVAL_2 == _EVAL_281;
  assign _EVAL_160 = ~_EVAL_299;
  assign _EVAL_181 = _EVAL_13 == _EVAL_203;
  assign _EVAL_170 = _EVAL_13[2:1];
  assign _EVAL_43 = _EVAL_170 == 2'h1;
  assign _EVAL_318 = _EVAL_17 == _EVAL_313;
  assign _EVAL_41 = _EVAL_35 | _EVAL_15;
  assign _EVAL_73 = _EVAL_122 | _EVAL_15;
  assign _EVAL_246 = _EVAL_210 | _EVAL_132;
  assign _EVAL_145 = _EVAL_34 | _EVAL_103;
  assign _EVAL_105 = _EVAL_305 | _EVAL_15;
  assign _EVAL_97 = _EVAL <= 3'h2;
  assign _EVAL_262 = _EVAL_50[7:0];
  assign _EVAL_93 = _EVAL_5 & _EVAL_138;
  assign _EVAL_267 = _EVAL_11 & _EVAL_176;
  assign _EVAL_290 = _EVAL_311 | _EVAL_15;
  assign _EVAL_44 = ~_EVAL_9;
  assign _EVAL_31 = _EVAL_144[5:0];
  assign _EVAL_209 = _EVAL_5 & _EVAL_302;
  assign _EVAL_241 = ~_EVAL_233;
  assign _EVAL_81 = {1'b0,$signed(_EVAL_30)};
  assign _EVAL_168 = _EVAL_65 | _EVAL_15;
  assign _EVAL_21 = _EVAL_232 | _EVAL_15;
  assign _EVAL_284 = _EVAL_136 & _EVAL_23;
  assign _EVAL_123 = _EVAL_56[5:0];
  assign _EVAL_294 = ~_EVAL_135;
  assign _EVAL_47 = _EVAL != 3'h0;
  assign _EVAL_234 = _EVAL_155 < plusarg_reader_out;
  assign _EVAL_111 = _EVAL_115 & _EVAL_38;
  assign _EVAL_291 = _EVAL_127 | _EVAL_88;
  assign _EVAL_108 = _EVAL_11 & _EVAL_128;
  assign _EVAL_176 = _EVAL_16 == 3'h5;
  assign _EVAL_77 = _EVAL_197 | _EVAL_104;
  assign _EVAL_115 = _EVAL_264 & _EVAL_75;
  assign _EVAL_240 = _EVAL_263[7:2];
  assign _EVAL_184 = ~_EVAL_290;
  assign _EVAL_167 = _EVAL_120 & _EVAL_227;
  assign _EVAL_225 = ~_EVAL_218;
  assign _EVAL_289 = _EVAL_22[5:0];
  assign _EVAL_56 = _EVAL_102 - 6'h1;
  assign _EVAL_112 = _EVAL_47 | _EVAL_15;
  assign _EVAL_237 = _EVAL_70 & _EVAL_307;
  assign _EVAL_59 = _EVAL_17 ^ 30'h3000;
  assign _EVAL_158 = _EVAL_27 | _EVAL_15;
  assign _EVAL_295 = _EVAL_251 | _EVAL_166;
  assign _EVAL_131 = ~_EVAL_306;
  assign _EVAL_152 = $signed(_EVAL_46) & -31'sh2000;
  assign _EVAL_207 = _EVAL_6 != 2'h2;
  assign _EVAL_42 = _EVAL_11 & _EVAL_293;
  assign _EVAL_100 = _EVAL_155 + 32'h1;
  assign _EVAL_186 = _EVAL_89 | _EVAL_140;
  assign _EVAL_177 = ~_EVAL_52;
  assign _EVAL_257 = _EVAL == 3'h0;
  assign _EVAL_107 = _EVAL_241 & _EVAL_306;
  assign _EVAL_196 = ~_EVAL_45;
  assign _EVAL_300 = _EVAL_11 & _EVAL_174;
  assign _EVAL_210 = _EVAL_64 & _EVAL_55;
  assign _EVAL_24 = _EVAL_1 == _EVAL_83;
  assign _EVAL_223 = ~_EVAL_222;
  assign _EVAL_148 = ~_EVAL_62;
  assign _EVAL_150 = _EVAL_6 <= 2'h2;
  assign _EVAL_195 = _EVAL_256[1];
  assign _EVAL_276 = _EVAL_121 == 6'h0;
  assign _EVAL_39 = _EVAL_120 & _EVAL_107;
  assign _EVAL_95 = _EVAL_195 & _EVAL_241;
  assign _EVAL_185 = {{22'd0}, _EVAL_263};
  assign _EVAL_268 = _EVAL_100[31:0];
  assign _EVAL_117 = _EVAL_18 == _EVAL_99;
  assign _EVAL_26 = _EVAL_117 | _EVAL_15;
  assign _EVAL_208 = _EVAL_194 >> _EVAL_13;
  assign _EVAL_84 = _EVAL_213 == 6'h0;
  assign _EVAL_143 = _EVAL_13 == 3'h4;
  assign _EVAL_183 = _EVAL_4 == _EVAL_301;
  assign _EVAL_141 = _EVAL_170 == 2'h0;
  assign _EVAL_180 = _EVAL_0 == 3'h4;
  assign _EVAL_147 = ~_EVAL_317;
  assign _EVAL_159 = _EVAL_264 & _EVAL_276;
  assign _EVAL_61 = _EVAL_70 | _EVAL_264;
  assign _EVAL_58 = _EVAL_164 | _EVAL_15;
  assign _EVAL_194 = _EVAL_88 | _EVAL_127;
  assign _EVAL_126 = _EVAL_220 | _EVAL_15;
  assign _EVAL_235 = _EVAL_1[0];
  assign _EVAL_314 = _EVAL_150 | _EVAL_15;
  assign _EVAL_214 = _EVAL_210 | _EVAL_151;
  assign _EVAL_132 = _EVAL_136 & _EVAL_72;
  assign _EVAL_98 = _EVAL_2[2:1];
  assign _EVAL_297 = _EVAL_208[0];
  assign _EVAL_139 = _EVAL_157 | _EVAL_15;
  assign _EVAL_35 = _EVAL_3 == _EVAL_266;
  assign _EVAL_280 = ~_EVAL_276;
  assign _EVAL_202 = 8'h1 << _EVAL_2;
  assign _EVAL_256 = _EVAL_94 | 2'h1;
  assign _EVAL_66 = _EVAL_20[7:0];
  assign _EVAL_75 = _EVAL_102 == 6'h0;
  assign _EVAL_104 = ~_EVAL_161;
  assign _EVAL_49 = _EVAL_17 ^ 30'h20000000;
  assign _EVAL_324 = ~_EVAL_200;
  assign _EVAL_29 = _EVAL_291 & _EVAL_242;
  assign _EVAL_199 = _EVAL_259[4:0];
  assign _EVAL_219 = ~_EVAL_168;
  assign _EVAL_298 = _EVAL_5 & _EVAL_178;
  assign _EVAL_38 = ~_EVAL_279;
  assign _EVAL_116 = _EVAL_183 | _EVAL_15;
  assign _EVAL_114 = _EVAL_0[0];
  assign _EVAL_227 = _EVAL_233 & _EVAL_131;
  assign _EVAL_230 = ~_EVAL_67;
  assign _EVAL_151 = _EVAL_136 & _EVAL_248;
  assign _EVAL_37 = _EVAL_0 == _EVAL_285;
  assign _EVAL_169 = _EVAL_273 | _EVAL_12;
  assign _EVAL_218 = _EVAL_40 | _EVAL_15;
  assign _EVAL_205 = _EVAL_5 & _EVAL_320;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_83 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_99 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_102 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_106 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_121 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_127 = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_155 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_203 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_213 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_258 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_270 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_281 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_285 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_286 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_301 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_309 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_313 = _RAND_16[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_8) begin
    if (_EVAL_211) begin
      _EVAL_83 <= _EVAL_1;
    end
    if (_EVAL_159) begin
      _EVAL_99 <= _EVAL_18;
    end
    if (_EVAL_15) begin
      _EVAL_102 <= 6'h0;
    end else if (_EVAL_264) begin
      if (_EVAL_75) begin
        if (_EVAL_114) begin
          _EVAL_102 <= _EVAL_236;
        end else begin
          _EVAL_102 <= 6'h0;
        end
      end else begin
        _EVAL_102 <= _EVAL_123;
      end
    end
    if (_EVAL_211) begin
      _EVAL_106 <= _EVAL;
    end
    if (_EVAL_15) begin
      _EVAL_121 <= 6'h0;
    end else if (_EVAL_264) begin
      if (_EVAL_276) begin
        if (_EVAL_114) begin
          _EVAL_121 <= _EVAL_236;
        end else begin
          _EVAL_121 <= 6'h0;
        end
      end else begin
        _EVAL_121 <= _EVAL_31;
      end
    end
    if (_EVAL_15) begin
      _EVAL_127 <= 5'h0;
    end else begin
      _EVAL_127 <= _EVAL_29;
    end
    if (_EVAL_15) begin
      _EVAL_155 <= 32'h0;
    end else if (_EVAL_61) begin
      _EVAL_155 <= 32'h0;
    end else begin
      _EVAL_155 <= _EVAL_268;
    end
    if (_EVAL_159) begin
      _EVAL_203 <= _EVAL_13;
    end
    if (_EVAL_15) begin
      _EVAL_213 <= 6'h0;
    end else if (_EVAL_70) begin
      if (_EVAL_84) begin
        if (_EVAL_177) begin
          _EVAL_213 <= _EVAL_240;
        end else begin
          _EVAL_213 <= 6'h0;
        end
      end else begin
        _EVAL_213 <= _EVAL_275;
      end
    end
    if (_EVAL_15) begin
      _EVAL_258 <= 6'h0;
    end else if (_EVAL_70) begin
      if (_EVAL_307) begin
        if (_EVAL_177) begin
          _EVAL_258 <= _EVAL_240;
        end else begin
          _EVAL_258 <= 6'h0;
        end
      end else begin
        _EVAL_258 <= _EVAL_289;
      end
    end
    if (_EVAL_211) begin
      _EVAL_270 <= _EVAL_16;
    end
    if (_EVAL_211) begin
      _EVAL_281 <= _EVAL_2;
    end
    if (_EVAL_159) begin
      _EVAL_285 <= _EVAL_0;
    end
    if (_EVAL_159) begin
      _EVAL_286 <= _EVAL_6;
    end
    if (_EVAL_159) begin
      _EVAL_301 <= _EVAL_4;
    end
    if (_EVAL_159) begin
      _EVAL_309 <= _EVAL_10;
    end
    if (_EVAL_211) begin
      _EVAL_313 <= _EVAL_17;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8428faf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d77b65ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90aae722)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(611d3b8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f478a69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(384b59e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_287) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36a4e27e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_319) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d034e8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d59053d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a89e372)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76d81914)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b3e90c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c579f6aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40ba1e8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_325) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c644570b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e93167ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d8a163a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39eddded)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19123089)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(524fb139)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4aef044)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5125e001)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd0e2ce4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db36575c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43da67f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89d9f565)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_319) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42b3ac1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68f5f053)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe4e764d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52ec8279)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_319) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c0e8c9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91493d0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(505eb8ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56b92340)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(893d4a91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fddc9f07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3314386d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d95fad5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_324) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(887056c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_324) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c67cbd9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc7c6af4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9479a1f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_304) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ffcc44c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a0ceb91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a3cf0d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b3af82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(610ceab8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a25b9d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_287) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_324) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf38762a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56383e95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_274) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4932cb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dca44891)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_294) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a735a469)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62f9fccd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d96cacd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5008eb29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_324) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ff626ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1da6d26c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f026b06e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84d75274)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6894f228)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1feea408)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a39b514)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f4c3b3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5eee380)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81bf773c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e55a53e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_294) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebb24a2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a0a2600)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45ea674d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb1e6dc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bb7d36a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2372ad37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0dce96a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23bbc7fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a427ffef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eee05a44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c981dfb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_319) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac6a588d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_325) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8acda915)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e10768cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87e38e13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8226cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be789897)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a00f49b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ed9fcf1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5182ba3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82f84f90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6b98ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(999c6a46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbb4149e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
