//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_128_assert(
  input        _EVAL,
  input  [8:0] _EVAL_0,
  input        _EVAL_1,
  input  [1:0] _EVAL_2,
  input        _EVAL_3,
  input  [2:0] _EVAL_4,
  input        _EVAL_5,
  input        _EVAL_6,
  input  [1:0] _EVAL_7,
  input        _EVAL_8,
  input  [2:0] _EVAL_9,
  input        _EVAL_10,
  input  [3:0] _EVAL_11,
  input        _EVAL_12,
  input        _EVAL_13,
  input        _EVAL_14
);
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  reg [1:0] _EVAL_19;
  reg [31:0] _RAND_0;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  reg [31:0] _EVAL_35;
  reg [31:0] _RAND_1;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire [1:0] _EVAL_44;
  reg [1:0] _EVAL_45;
  reg [31:0] _RAND_2;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  reg  _EVAL_56;
  reg [31:0] _RAND_3;
  wire  _EVAL_57;
  reg  _EVAL_58;
  reg [31:0] _RAND_4;
  wire [8:0] _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  reg  _EVAL_63;
  reg [31:0] _RAND_5;
  wire  _EVAL_64;
  wire  _EVAL_65;
  reg [2:0] _EVAL_66;
  reg [31:0] _RAND_6;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire [9:0] _EVAL_75;
  reg [8:0] _EVAL_76;
  reg [31:0] _RAND_7;
  wire  _EVAL_77;
  wire [8:0] _EVAL_78;
  wire [9:0] _EVAL_79;
  wire  _EVAL_80;
  wire [9:0] _EVAL_81;
  wire [9:0] _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire [1:0] _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire [9:0] _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  reg  _EVAL_97;
  reg [31:0] _RAND_8;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire [9:0] _EVAL_102;
  wire [8:0] _EVAL_103;
  wire  _EVAL_104;
  wire [9:0] _EVAL_105;
  wire  _EVAL_106;
  wire [9:0] _EVAL_107;
  wire  _EVAL_108;
  reg  _EVAL_109;
  reg [31:0] _RAND_9;
  wire [9:0] _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire [9:0] _EVAL_113;
  wire [9:0] _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire [9:0] _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire [9:0] _EVAL_136;
  wire  _EVAL_137;
  reg  _EVAL_138;
  reg [31:0] _RAND_10;
  wire [9:0] _EVAL_139;
  wire [9:0] _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire [1:0] _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_147;
  wire [3:0] _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire [31:0] _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire [8:0] _EVAL_158;
  wire  _EVAL_159;
  wire [9:0] _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  reg  _EVAL_166;
  reg [31:0] _RAND_11;
  wire [1:0] _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire [8:0] _EVAL_172;
  wire  _EVAL_173;
  reg  _EVAL_174;
  reg [31:0] _RAND_12;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire [1:0] _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire [1:0] _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire [32:0] _EVAL_186;
  wire [8:0] _EVAL_187;
  wire  _EVAL_189;
  wire [9:0] _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire [9:0] _EVAL_193;
  reg [2:0] _EVAL_194;
  reg [31:0] _RAND_13;
  wire  _EVAL_195;
  wire [1:0] _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_107 = $signed(_EVAL_113) & -10'sh80;
  assign _EVAL_98 = ~_EVAL_77;
  assign _EVAL_75 = {1'b0,$signed(_EVAL_187)};
  assign _EVAL_122 = ~_EVAL_138;
  assign _EVAL_158 = _EVAL_0 ^ 9'h100;
  assign _EVAL_34 = _EVAL_9 <= 3'h6;
  assign _EVAL_100 = ~_EVAL_153;
  assign _EVAL_39 = _EVAL_34 | _EVAL_115;
  assign _EVAL_130 = _EVAL_170 & _EVAL_94;
  assign _EVAL_126 = ~_EVAL_28;
  assign _EVAL_61 = _EVAL_163 | _EVAL_115;
  assign _EVAL_74 = ~_EVAL_177;
  assign _EVAL_105 = $signed(_EVAL_160) & -10'sh18;
  assign _EVAL_135 = ~_EVAL_56;
  assign _EVAL_26 = ~_EVAL_135;
  assign _EVAL_70 = plusarg_reader_out == 32'h0;
  assign _EVAL_207 = ~_EVAL_25;
  assign _EVAL_192 = ~_EVAL_181;
  assign _EVAL_153 = _EVAL_65 | _EVAL_115;
  assign _EVAL_131 = _EVAL_4 == 3'h7;
  assign _EVAL_211 = _EVAL_6 & _EVAL_26;
  assign _EVAL_145 = ~_EVAL_161;
  assign _EVAL_41 = _EVAL_196[0];
  assign _EVAL_106 = _EVAL_2 == 2'h0;
  assign _EVAL_203 = _EVAL_9 == 3'h0;
  assign _EVAL_60 = _EVAL_210 | _EVAL_115;
  assign _EVAL_91 = $signed(_EVAL_110) == 10'sh0;
  assign _EVAL_175 = $signed(_EVAL_140) == 10'sh0;
  assign _EVAL_29 = _EVAL_197 | _EVAL_70;
  assign _EVAL_182 = _EVAL_4 == 3'h4;
  assign _EVAL_42 = _EVAL_6 & _EVAL_111;
  assign _EVAL_54 = _EVAL_197 | _EVAL_115;
  assign _EVAL_129 = _EVAL_109 | _EVAL_46;
  assign _EVAL_50 = _EVAL_157 | _EVAL_115;
  assign _EVAL_142 = _EVAL_7 == _EVAL_45;
  assign _EVAL_208 = _EVAL_2 == _EVAL_19;
  assign _EVAL_123 = _EVAL_149 | _EVAL_115;
  assign _EVAL_191 = _EVAL_208 | _EVAL_115;
  assign _EVAL_128 = _EVAL_48 | _EVAL_30;
  assign _EVAL_48 = _EVAL_175 | _EVAL_22;
  assign _EVAL_171 = _EVAL_65 | _EVAL_10;
  assign _EVAL_116 = _EVAL_12 & _EVAL_6;
  assign _EVAL_68 = _EVAL_14 & _EVAL_182;
  assign _EVAL_127 = {1'b0,$signed(_EVAL_0)};
  assign _EVAL_28 = _EVAL_195 | _EVAL_115;
  assign _EVAL_181 = _EVAL_179 | _EVAL_115;
  assign _EVAL_84 = _EVAL_106 | _EVAL_115;
  assign _EVAL_201 = _EVAL_128 | _EVAL_91;
  assign _EVAL_20 = ~_EVAL_156;
  assign _EVAL_55 = _EVAL_0 == _EVAL_76;
  assign _EVAL_18 = _EVAL_51 | _EVAL_115;
  assign _EVAL_114 = $signed(_EVAL_75) & -10'sh4;
  assign _EVAL_95 = ~_EVAL_50;
  assign _EVAL_80 = _EVAL_108 | _EVAL_115;
  assign _EVAL_94 = ~_EVAL_63;
  assign _EVAL_205 = _EVAL_125 | _EVAL_115;
  assign _EVAL_176 = ~_EVAL_52;
  assign _EVAL_165 = _EVAL_21 | _EVAL_115;
  assign _EVAL_52 = _EVAL_209 | _EVAL_115;
  assign _EVAL_81 = $signed(_EVAL_82) & -10'sh100;
  assign _EVAL_199 = _EVAL_183[0];
  assign _EVAL_44 = _EVAL_38 ? _EVAL_89 : 2'h0;
  assign _EVAL_15 = _EVAL_14 & _EVAL_131;
  assign _EVAL_148 = ~_EVAL_11;
  assign _EVAL_187 = _EVAL_0 ^ 9'h44;
  assign _EVAL_137 = _EVAL_144[0];
  assign _EVAL_161 = _EVAL_168 | _EVAL_115;
  assign _EVAL_27 = ~_EVAL_32;
  assign _EVAL_49 = ~_EVAL_205;
  assign _EVAL_112 = _EVAL_9 == 3'h1;
  assign _EVAL_59 = _EVAL_0 ^ 9'h80;
  assign _EVAL_88 = _EVAL_55 | _EVAL_115;
  assign _EVAL_82 = {1'b0,$signed(_EVAL_158)};
  assign _EVAL_140 = _EVAL_190;
  assign _EVAL_120 = ~_EVAL_165;
  assign _EVAL_43 = _EVAL_167[0];
  assign _EVAL_36 = _EVAL_14 & _EVAL_162;
  assign _EVAL_177 = _EVAL_96 | _EVAL_115;
  assign _EVAL_150 = _EVAL_14 & _EVAL_87;
  assign _EVAL_93 = _EVAL_105;
  assign _EVAL_21 = _EVAL_13 == _EVAL_97;
  assign _EVAL_155 = _EVAL_4 == 3'h3;
  assign _EVAL_108 = _EVAL_92 | _EVAL_69;
  assign _EVAL_125 = _EVAL_4 == _EVAL_66;
  assign _EVAL_212 = _EVAL_46 | _EVAL_109;
  assign _EVAL_46 = _EVAL_178[0];
  assign _EVAL_141 = ~_EVAL_54;
  assign _EVAL_64 = _EVAL_6 & _EVAL_104;
  assign _EVAL_160 = {1'b0,$signed(_EVAL_78)};
  assign _EVAL_134 = ~_EVAL_191;
  assign _EVAL_154 = _EVAL_171 | _EVAL_115;
  assign _EVAL_197 = ~_EVAL_109;
  assign _EVAL_102 = {1'b0,$signed(_EVAL_172)};
  assign _EVAL_157 = _EVAL_11 == 4'hf;
  assign _EVAL_156 = _EVAL_37 | _EVAL_115;
  assign _EVAL_30 = $signed(_EVAL_93) == 10'sh0;
  assign _EVAL_167 = _EVAL_174 - 1'h1;
  assign _EVAL_117 = _EVAL_142 | _EVAL_115;
  assign _EVAL_136 = _EVAL_107;
  assign _EVAL_209 = _EVAL_2 != 2'h2;
  assign _EVAL_184 = _EVAL_4 == 3'h5;
  assign _EVAL_186 = _EVAL_35 + 32'h1;
  assign _EVAL_111 = _EVAL_9 == 3'h4;
  assign _EVAL_163 = _EVAL_148 == 4'h0;
  assign _EVAL_190 = $signed(_EVAL_127) & -10'sh40;
  assign _EVAL_24 = _EVAL_170 | _EVAL_116;
  assign _EVAL_17 = ~_EVAL_200;
  assign _EVAL_77 = _EVAL_85 | _EVAL_115;
  assign _EVAL_210 = ~_EVAL_13;
  assign _EVAL_113 = {1'b0,$signed(_EVAL_59)};
  assign _EVAL_101 = _EVAL_14 & _EVAL_121;
  assign _EVAL_206 = ~_EVAL_61;
  assign _EVAL_92 = _EVAL_201 | _EVAL_124;
  assign _EVAL_185 = _EVAL_14 & _EVAL_202;
  assign _EVAL_202 = ~_EVAL_159;
  assign _EVAL_47 = _EVAL_119 | _EVAL_115;
  assign _EVAL_71 = ~_EVAL_117;
  assign _EVAL_32 = _EVAL_44[0];
  assign _EVAL_90 = ~_EVAL_84;
  assign _EVAL_151 = _EVAL_186[31:0];
  assign _EVAL_67 = _EVAL_6 & _EVAL_203;
  assign _EVAL_96 = _EVAL_3 == _EVAL_58;
  assign _EVAL_23 = _EVAL_6 & _EVAL_86;
  assign _EVAL_85 = _EVAL_212 >> _EVAL_13;
  assign _EVAL_40 = _EVAL_6 & _EVAL_112;
  assign _EVAL_143 = _EVAL_170 & _EVAL_159;
  assign _EVAL_121 = _EVAL_4 == 3'h6;
  assign _EVAL_73 = ~_EVAL_46;
  assign _EVAL_51 = _EVAL_103 == 9'h0;
  assign _EVAL_25 = _EVAL_9 == 3'h6;
  assign _EVAL_79 = _EVAL_81;
  assign _EVAL_37 = ~_EVAL_10;
  assign _EVAL_139 = _EVAL_114;
  assign _EVAL_172 = _EVAL_0 ^ 9'h60;
  assign _EVAL_38 = _EVAL_16 & _EVAL_207;
  assign _EVAL_179 = _EVAL_8 == _EVAL_166;
  assign _EVAL_196 = _EVAL_56 - 1'h1;
  assign _EVAL_53 = _EVAL_116 & _EVAL_135;
  assign _EVAL_159 = ~_EVAL_174;
  assign _EVAL_173 = ~_EVAL_80;
  assign _EVAL_124 = $signed(_EVAL_136) == 10'sh0;
  assign _EVAL_144 = _EVAL_138 - 1'h1;
  assign _EVAL_78 = _EVAL_0 ^ 9'h48;
  assign _EVAL_89 = 2'h1 << _EVAL_13;
  assign _EVAL_162 = _EVAL_4 == 3'h2;
  assign _EVAL_69 = $signed(_EVAL_79) == 10'sh0;
  assign _EVAL_86 = _EVAL_9 == 3'h2;
  assign _EVAL_198 = ~_EVAL_154;
  assign _EVAL_147 = ~_EVAL_88;
  assign _EVAL_33 = ~_EVAL_123;
  assign _EVAL_115 = _EVAL_5;
  assign _EVAL_103 = _EVAL_0 & 9'h3;
  assign _EVAL_178 = _EVAL_130 ? 2'h1 : 2'h0;
  assign _EVAL_132 = _EVAL_14 & _EVAL_184;
  assign _EVAL_200 = _EVAL_57 | _EVAL_115;
  assign _EVAL_65 = ~_EVAL_8;
  assign _EVAL_57 = _EVAL_2 <= 2'h2;
  assign _EVAL_133 = _EVAL_14 & _EVAL_31;
  assign _EVAL_62 = _EVAL_6 & _EVAL_25;
  assign _EVAL_169 = ~_EVAL_47;
  assign _EVAL_204 = ~_EVAL_115;
  assign _EVAL_164 = _EVAL_46 != _EVAL_32;
  assign _EVAL_193 = $signed(_EVAL_102) & -10'sh20;
  assign _EVAL_183 = _EVAL_63 - 1'h1;
  assign _EVAL_168 = _EVAL_29 | _EVAL_152;
  assign _EVAL_119 = _EVAL_164 | _EVAL_73;
  assign _EVAL_195 = _EVAL_7 >= 2'h2;
  assign _EVAL_16 = _EVAL_116 & _EVAL_122;
  assign _EVAL_83 = ~_EVAL_60;
  assign _EVAL_149 = _EVAL_9 == _EVAL_194;
  assign _EVAL_99 = _EVAL_14 & _EVAL_155;
  assign _EVAL_104 = _EVAL_9 == 3'h5;
  assign _EVAL_22 = $signed(_EVAL_139) == 10'sh0;
  assign _EVAL_152 = _EVAL_35 < plusarg_reader_out;
  assign _EVAL_87 = _EVAL_4 == 3'h0;
  assign _EVAL_118 = ~_EVAL_18;
  assign _EVAL_110 = _EVAL_193;
  assign _EVAL_189 = ~_EVAL_39;
  assign _EVAL_31 = _EVAL_4 == 3'h1;
  assign _EVAL_170 = _EVAL_1 & _EVAL_14;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_19 = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_35 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_45 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_56 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_58 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_63 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_66 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_76 = _RAND_7[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_97 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_109 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_138 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_166 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_174 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_194 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  if (_EVAL_5) begin
    _EVAL_35 = 32'h0;
  end
  if (_EVAL_5) begin
    _EVAL_56 = 1'h0;
  end
  if (_EVAL_5) begin
    _EVAL_63 = 1'h0;
  end
  if (_EVAL_5) begin
    _EVAL_109 = 1'h0;
  end
  if (_EVAL_5) begin
    _EVAL_138 = 1'h0;
  end
  if (_EVAL_5) begin
    _EVAL_174 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL) begin
    if (_EVAL_53) begin
      _EVAL_19 <= _EVAL_2;
    end
    if (_EVAL_53) begin
      _EVAL_45 <= _EVAL_7;
    end
    if (_EVAL_53) begin
      _EVAL_58 <= _EVAL_3;
    end
    if (_EVAL_143) begin
      _EVAL_66 <= _EVAL_4;
    end
    if (_EVAL_143) begin
      _EVAL_76 <= _EVAL_0;
    end
    if (_EVAL_53) begin
      _EVAL_97 <= _EVAL_13;
    end
    if (_EVAL_53) begin
      _EVAL_166 <= _EVAL_8;
    end
    if (_EVAL_53) begin
      _EVAL_194 <= _EVAL_9;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37492696)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81707802)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(957bd015)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(236403ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57e22c91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8ba45bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdd7b19d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(844086e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc0cff4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a98b4a1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fa1f5e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40e3b2d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c854aa44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71e57c02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23d4a95f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2111838)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7881ad44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1331bbc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c844693)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bba917c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1f04661)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f23f1c66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92fd31cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe822b00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a4040ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c338041)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(626b6d34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(931cf324)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3fdb3f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a24ebfdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(110eb0d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f025ce70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67634f02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(956c0ed9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b52bed78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e95488ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92a43d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f70ef477)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(576bf4b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d201084c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11daf33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfb9aa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fae4995)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65b19d39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c18e991a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5dc59ee5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(659374c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5684ae8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee69534c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a997895)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec4ac0a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e52482e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ffb2ad8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(772cd13a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f33001f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3aa279e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd49a342)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72cde62c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96c6def9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbb34d5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5df39e07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ed9bbe5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5834b5bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99a24102)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0a1efb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5b50bd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(998f99af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6fb575e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5351dabb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd10bc28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge _EVAL or posedge _EVAL_5) begin
    if (_EVAL_5) begin
      _EVAL_35 <= 32'h0;
    end else if (_EVAL_24) begin
      _EVAL_35 <= 32'h0;
    end else begin
      _EVAL_35 <= _EVAL_151;
    end
  end
  always @(posedge _EVAL or posedge _EVAL_5) begin
    if (_EVAL_5) begin
      _EVAL_56 <= 1'h0;
    end else if (_EVAL_116) begin
      if (_EVAL_135) begin
        _EVAL_56 <= 1'h0;
      end else begin
        _EVAL_56 <= _EVAL_41;
      end
    end
  end
  always @(posedge _EVAL or posedge _EVAL_5) begin
    if (_EVAL_5) begin
      _EVAL_63 <= 1'h0;
    end else if (_EVAL_170) begin
      if (_EVAL_94) begin
        _EVAL_63 <= 1'h0;
      end else begin
        _EVAL_63 <= _EVAL_199;
      end
    end
  end
  always @(posedge _EVAL or posedge _EVAL_5) begin
    if (_EVAL_5) begin
      _EVAL_109 <= 1'h0;
    end else begin
      _EVAL_109 <= _EVAL_129 & _EVAL_27;
    end
  end
  always @(posedge _EVAL or posedge _EVAL_5) begin
    if (_EVAL_5) begin
      _EVAL_138 <= 1'h0;
    end else if (_EVAL_116) begin
      if (_EVAL_122) begin
        _EVAL_138 <= 1'h0;
      end else begin
        _EVAL_138 <= _EVAL_137;
      end
    end
  end
  always @(posedge _EVAL or posedge _EVAL_5) begin
    if (_EVAL_5) begin
      _EVAL_174 <= 1'h0;
    end else if (_EVAL_170) begin
      if (_EVAL_159) begin
        _EVAL_174 <= 1'h0;
      end else begin
        _EVAL_174 <= _EVAL_43;
      end
    end
  end

endmodule
