//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_159_assert(
  input  [3:0]  _EVAL,
  input         _EVAL_0,
  input  [3:0]  _EVAL_1,
  input  [31:0] _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input  [1:0]  _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [2:0]  _EVAL_17,
  input  [3:0]  _EVAL_18
);
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire [22:0] _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire [32:0] _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire [5:0] _EVAL_37;
  wire [6:0] _EVAL_38;
  wire  _EVAL_39;
  wire [31:0] _EVAL_40;
  wire [31:0] _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire [31:0] plusarg_reader_out;
  wire [7:0] _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire [1:0] _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire [32:0] _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_62;
  wire [3:0] _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire [32:0] _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire [32:0] _EVAL_70;
  wire  _EVAL_71;
  reg [2:0] _EVAL_72;
  reg [31:0] _RAND_0;
  wire [32:0] _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire [1:0] _EVAL_77;
  reg [31:0] _EVAL_78;
  reg [31:0] _RAND_1;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire [32:0] _EVAL_82;
  wire [31:0] _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire [1:0] _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire [32:0] _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  reg [31:0] _EVAL_98;
  reg [31:0] _RAND_2;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire [1:0] _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire [5:0] _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire [32:0] _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire [7:0] _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire [1:0] _EVAL_120;
  wire  _EVAL_121;
  wire [31:0] _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire [32:0] _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_133;
  wire [32:0] _EVAL_134;
  wire [32:0] _EVAL_135;
  wire  _EVAL_136;
  wire [6:0] _EVAL_137;
  reg [1:0] _EVAL_138;
  reg [31:0] _RAND_3;
  wire [31:0] _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire [22:0] _EVAL_142;
  wire  _EVAL_143;
  wire [31:0] _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  reg  _EVAL_150;
  reg [31:0] _RAND_4;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  reg [3:0] _EVAL_158;
  reg [31:0] _RAND_5;
  wire [1:0] _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  reg [5:0] _EVAL_172;
  reg [31:0] _RAND_6;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  reg [1:0] _EVAL_177;
  reg [31:0] _RAND_7;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  reg [2:0] _EVAL_184;
  reg [31:0] _RAND_8;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire [5:0] _EVAL_190;
  wire  _EVAL_191;
  reg  _EVAL_192;
  reg [31:0] _RAND_9;
  wire  _EVAL_194;
  wire [32:0] _EVAL_195;
  wire [32:0] _EVAL_196;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire [5:0] _EVAL_202;
  wire [1:0] _EVAL_203;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire [32:0] _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire [32:0] _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire [6:0] _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire [32:0] _EVAL_229;
  wire  _EVAL_230;
  wire [1:0] _EVAL_231;
  wire  _EVAL_232;
  reg [5:0] _EVAL_234;
  reg [31:0] _RAND_10;
  reg [3:0] _EVAL_235;
  reg [31:0] _RAND_11;
  wire [32:0] _EVAL_236;
  wire [32:0] _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  reg  _EVAL_240;
  reg [31:0] _RAND_12;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire [31:0] _EVAL_246;
  wire  _EVAL_248;
  wire [1:0] _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire [5:0] _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire [31:0] _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  reg [5:0] _EVAL_259;
  reg [31:0] _RAND_13;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire [6:0] _EVAL_263;
  wire [1:0] _EVAL_264;
  reg [5:0] _EVAL_265;
  reg [31:0] _RAND_14;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire [3:0] _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_274;
  wire  _EVAL_275;
  reg  _EVAL_276;
  reg [31:0] _RAND_15;
  wire  _EVAL_277;
  wire [3:0] _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire [3:0] _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire [1:0] _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire [1:0] _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire [5:0] _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  reg [2:0] _EVAL_311;
  reg [31:0] _RAND_16;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire [7:0] _EVAL_318;
  wire [7:0] _EVAL_319;
  wire  _EVAL_320;
  wire  _EVAL_321;
  wire  _EVAL_322;
  wire [32:0] _EVAL_323;
  wire  _EVAL_324;
  wire  _EVAL_325;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_219 = _EVAL_99 & _EVAL_29;
  assign _EVAL_136 = _EVAL_1[0];
  assign _EVAL_250 = ~_EVAL_13;
  assign _EVAL_280 = ~_EVAL_166;
  assign _EVAL_324 = ~_EVAL_320;
  assign _EVAL_129 = ~_EVAL_69;
  assign _EVAL_294 = _EVAL_5 == 3'h6;
  assign _EVAL_123 = _EVAL_14 & _EVAL_106;
  assign _EVAL_95 = _EVAL_134;
  assign _EVAL_37 = _EVAL_226[5:0];
  assign _EVAL_160 = plusarg_reader_out == 32'h0;
  assign _EVAL_320 = _EVAL_255 | _EVAL_6;
  assign _EVAL_142 = 23'hff << _EVAL_1;
  assign _EVAL_157 = _EVAL_99 & _EVAL_287;
  assign _EVAL_56 = ~_EVAL_297;
  assign _EVAL_176 = ~_EVAL_261;
  assign _EVAL_87 = _EVAL_283 | _EVAL_6;
  assign _EVAL_22 = 23'hff << _EVAL_18;
  assign _EVAL_52 = _EVAL_321 | _EVAL_6;
  assign _EVAL_261 = _EVAL_25 | _EVAL_6;
  assign _EVAL_57 = _EVAL_127 | _EVAL_6;
  assign _EVAL_322 = ~_EVAL_218;
  assign _EVAL_77 = _EVAL_177 | _EVAL_249;
  assign _EVAL_120 = _EVAL_165 ? _EVAL_301 : 2'h0;
  assign _EVAL_256 = _EVAL_26[31:0];
  assign _EVAL_147 = _EVAL_4 & _EVAL_14;
  assign _EVAL_186 = _EVAL_227 | _EVAL_64;
  assign _EVAL_71 = _EVAL_105 | _EVAL_188;
  assign _EVAL_216 = _EVAL_42 | _EVAL_6;
  assign _EVAL_321 = ~_EVAL_0;
  assign _EVAL_303 = _EVAL == _EVAL_269;
  assign _EVAL_58 = _EVAL_236;
  assign _EVAL_302 = _EVAL_12 & _EVAL_294;
  assign _EVAL_49 = _EVAL_131 | _EVAL_6;
  assign _EVAL_208 = _EVAL_283 | _EVAL_80;
  assign _EVAL_159 = _EVAL_177 >> _EVAL_15;
  assign _EVAL_105 = _EVAL_274 & _EVAL_181;
  assign _EVAL_191 = _EVAL_59 | _EVAL_6;
  assign _EVAL_251 = _EVAL_2[1];
  assign _EVAL_196 = _EVAL_73;
  assign _EVAL_152 = _EVAL_7 == 2'h0;
  assign _EVAL_30 = _EVAL_296 | _EVAL_6;
  assign _EVAL_284 = _EVAL_133 & _EVAL_251;
  assign _EVAL_66 = _EVAL_323;
  assign _EVAL_65 = ~_EVAL_84;
  assign _EVAL_270 = _EVAL_177 != 2'h0;
  assign _EVAL_281 = _EVAL_17[0];
  assign _EVAL_325 = _EVAL_210 | _EVAL_6;
  assign _EVAL_133 = _EVAL_107[1];
  assign _EVAL_69 = _EVAL_93 | _EVAL_6;
  assign _EVAL_180 = _EVAL_175 | _EVAL_315;
  assign _EVAL_243 = _EVAL_155 & _EVAL_157;
  assign _EVAL_169 = _EVAL_14 & _EVAL_271;
  assign _EVAL_317 = $signed(_EVAL_196) == 33'sh0;
  assign _EVAL_185 = _EVAL_12 & _EVAL_300;
  assign _EVAL_174 = _EVAL_5 == 3'h4;
  assign _EVAL_189 = _EVAL_17 == 3'h4;
  assign _EVAL_210 = _EVAL_241 | _EVAL_188;
  assign _EVAL_171 = _EVAL_5 == 3'h2;
  assign _EVAL_108 = _EVAL_152 | _EVAL_6;
  assign _EVAL_111 = _EVAL_25 | _EVAL_13;
  assign _EVAL_26 = _EVAL_98 + 32'h1;
  assign _EVAL_76 = _EVAL_111 | _EVAL_6;
  assign _EVAL_127 = ~_EVAL_35;
  assign _EVAL_190 = _EVAL_137[5:0];
  assign _EVAL_198 = _EVAL_23 | _EVAL_6;
  assign _EVAL_124 = _EVAL_17 <= 3'h6;
  assign _EVAL_33 = _EVAL_12 & _EVAL_262;
  assign _EVAL_173 = _EVAL_231[0];
  assign _EVAL_308 = ~_EVAL_143;
  assign _EVAL_293 = _EVAL_172 == 6'h0;
  assign _EVAL_262 = _EVAL_5 == 3'h5;
  assign _EVAL_154 = _EVAL_9 <= 3'h4;
  assign _EVAL_102 = _EVAL_147 & _EVAL_312;
  assign _EVAL_148 = _EVAL_180 | _EVAL_88;
  assign _EVAL_54 = _EVAL_250 | _EVAL_6;
  assign _EVAL_223 = _EVAL_251 & _EVAL_29;
  assign _EVAL_131 = _EVAL_71 | _EVAL_314;
  assign _EVAL_230 = _EVAL_154 | _EVAL_6;
  assign _EVAL_306 = _EVAL_263[5:0];
  assign _EVAL_178 = _EVAL_258 | _EVAL_6;
  assign _EVAL_92 = ~_EVAL_244;
  assign _EVAL_93 = _EVAL_9 != 3'h0;
  assign _EVAL_291 = ~_EVAL_325;
  assign _EVAL_114 = _EVAL_10 == _EVAL_192;
  assign _EVAL_70 = $signed(_EVAL_113) & -33'sh1000;
  assign _EVAL_44 = _EVAL_22[7:0];
  assign _EVAL_86 = _EVAL_7 != 2'h2;
  assign _EVAL_146 = _EVAL_7 <= 2'h2;
  assign _EVAL_229 = {1'b0,$signed(_EVAL_40)};
  assign _EVAL_255 = _EVAL_47 & _EVAL_148;
  assign _EVAL_232 = ~_EVAL_245;
  assign _EVAL_200 = _EVAL_155 & _EVAL_85;
  assign _EVAL_166 = _EVAL_205 | _EVAL_6;
  assign _EVAL_257 = _EVAL_9 == 3'h0;
  assign _EVAL_246 = _EVAL_2 ^ 32'h80000000;
  assign _EVAL_202 = _EVAL_117[7:2];
  assign _EVAL_80 = _EVAL_133 & _EVAL_99;
  assign _EVAL_279 = ~_EVAL_125;
  assign _EVAL_297 = _EVAL_249 != 2'h0;
  assign _EVAL_286 = _EVAL_147 & _EVAL_242;
  assign _EVAL_211 = _EVAL_237;
  assign _EVAL_239 = _EVAL_5[2];
  assign _EVAL_101 = _EVAL_282 | _EVAL_6;
  assign _EVAL_167 = _EVAL_12 & _EVAL_141;
  assign _EVAL_236 = $signed(_EVAL_195) & -33'sh2000;
  assign _EVAL_110 = _EVAL_38[5:0];
  assign _EVAL_312 = _EVAL_234 == 6'h0;
  assign _EVAL_201 = ~_EVAL_198;
  assign _EVAL_310 = _EVAL_5 == 3'h0;
  assign _EVAL_258 = _EVAL_32 | _EVAL_56;
  assign _EVAL_274 = _EVAL_1 <= 4'h6;
  assign _EVAL_161 = _EVAL_155 & _EVAL_219;
  assign _EVAL_85 = _EVAL_251 & _EVAL_287;
  assign _EVAL_181 = $signed(_EVAL_58) == 33'sh0;
  assign _EVAL_179 = _EVAL_5 == 3'h1;
  assign _EVAL_134 = $signed(_EVAL_214) & -33'shc000;
  assign _EVAL_268 = _EVAL_14 & _EVAL_260;
  assign _EVAL_113 = {1'b0,$signed(_EVAL_122)};
  assign _EVAL_20 = ~_EVAL_39;
  assign _EVAL_115 = ~_EVAL_76;
  assign _EVAL_100 = ~_EVAL_109;
  assign _EVAL_63 = ~_EVAL_269;
  assign _EVAL_316 = _EVAL_303 | _EVAL_6;
  assign _EVAL_96 = _EVAL_12 & _EVAL_179;
  assign _EVAL_218 = _EVAL_151 | _EVAL_6;
  assign _EVAL_313 = _EVAL_145 | _EVAL_6;
  assign _EVAL_83 = _EVAL_2 & _EVAL_144;
  assign _EVAL_209 = _EVAL_187 | _EVAL_6;
  assign _EVAL_307 = _EVAL_18 >= 4'h2;
  assign _EVAL_213 = ~_EVAL_36;
  assign _EVAL_73 = $signed(_EVAL_229) & -33'sh1000000;
  assign _EVAL_315 = $signed(_EVAL_66) == 33'sh0;
  assign _EVAL_41 = _EVAL_2 ^ 32'h20000000;
  assign _EVAL_309 = ~_EVAL_270;
  assign _EVAL_289 = _EVAL_12 & _EVAL_168;
  assign _EVAL_31 = _EVAL_9 <= 3'h3;
  assign _EVAL_143 = _EVAL_146 | _EVAL_6;
  assign _EVAL_225 = _EVAL_12 & _EVAL_174;
  assign _EVAL_267 = _EVAL_31 | _EVAL_6;
  assign _EVAL_241 = _EVAL_47 & _EVAL_19;
  assign _EVAL_46 = _EVAL_2 == _EVAL_78;
  assign _EVAL_224 = ~_EVAL_87;
  assign _EVAL_194 = _EVAL_14 & _EVAL_140;
  assign _EVAL_305 = _EVAL_307 | _EVAL_6;
  assign _EVAL_59 = _EVAL_9 <= 3'h1;
  assign _EVAL_298 = ~_EVAL_120;
  assign _EVAL_34 = $signed(_EVAL_126) == 33'sh0;
  assign _EVAL_269 = {_EVAL_164,_EVAL_186,_EVAL_119,_EVAL_206};
  assign _EVAL_222 = _EVAL_17 == 3'h2;
  assign _EVAL_145 = _EVAL_292 == 4'h0;
  assign _EVAL_43 = _EVAL_5 == _EVAL_72;
  assign _EVAL_238 = _EVAL_254 & _EVAL_75;
  assign _EVAL_227 = _EVAL_283 | _EVAL_284;
  assign _EVAL_212 = ~_EVAL_272;
  assign _EVAL_89 = _EVAL_77 & _EVAL_298;
  assign _EVAL_25 = ~_EVAL_10;
  assign _EVAL_104 = ~_EVAL_316;
  assign _EVAL_287 = _EVAL_2[0];
  assign _EVAL_283 = _EVAL_1 >= 4'h2;
  assign _EVAL_107 = _EVAL_264 | 2'h1;
  assign _EVAL_144 = {{24'd0}, _EVAL_318};
  assign _EVAL_126 = _EVAL_70;
  assign _EVAL_296 = _EVAL_7 == _EVAL_138;
  assign _EVAL_99 = ~_EVAL_251;
  assign _EVAL_38 = _EVAL_172 - 6'h1;
  assign _EVAL_90 = ~_EVAL_178;
  assign _EVAL_271 = ~_EVAL_242;
  assign _EVAL_228 = _EVAL_27 | _EVAL_183;
  assign _EVAL_125 = _EVAL_128 | _EVAL_6;
  assign _EVAL_199 = _EVAL_83 == 32'h0;
  assign _EVAL_141 = _EVAL_5 == 3'h7;
  assign _EVAL_40 = _EVAL_2 ^ 32'h2000000;
  assign _EVAL_263 = _EVAL_234 - 6'h1;
  assign _EVAL_121 = _EVAL_124 | _EVAL_6;
  assign _EVAL_155 = _EVAL_107[0];
  assign _EVAL_203 = _EVAL_249 | _EVAL_177;
  assign _EVAL_50 = ~_EVAL_130;
  assign _EVAL_139 = _EVAL_2 ^ 32'h40000000;
  assign _EVAL_252 = ~_EVAL_30;
  assign _EVAL_135 = {1'b0,$signed(_EVAL_2)};
  assign _EVAL_39 = _EVAL_43 | _EVAL_6;
  assign _EVAL_64 = _EVAL_155 & _EVAL_223;
  assign _EVAL_217 = _EVAL_15 == _EVAL_240;
  assign _EVAL_60 = _EVAL_14 & _EVAL_189;
  assign _EVAL_122 = _EVAL_2 ^ 32'h3000;
  assign _EVAL_153 = _EVAL_14 & _EVAL_116;
  assign _EVAL_248 = _EVAL_74 | _EVAL_6;
  assign _EVAL_195 = {1'b0,$signed(_EVAL_139)};
  assign _EVAL_82 = {1'b0,$signed(_EVAL_41)};
  assign _EVAL_103 = ~_EVAL_108;
  assign _EVAL_67 = ~_EVAL_191;
  assign _EVAL_314 = _EVAL_47 & _EVAL_88;
  assign _EVAL_35 = _EVAL_159[0];
  assign _EVAL_323 = $signed(_EVAL_135) & -33'sh5000;
  assign _EVAL_36 = _EVAL_228 | _EVAL_6;
  assign _EVAL_168 = ~_EVAL_293;
  assign _EVAL_97 = _EVAL_1 <= 4'h8;
  assign _EVAL_237 = $signed(_EVAL_82) & -33'sh2000;
  assign _EVAL_260 = _EVAL_17 == 3'h6;
  assign _EVAL_226 = _EVAL_259 - 6'h1;
  assign _EVAL_156 = ~_EVAL_230;
  assign _EVAL_68 = ~_EVAL_121;
  assign _EVAL_23 = _EVAL_8 == _EVAL_150;
  assign _EVAL_118 = ~_EVAL_49;
  assign _EVAL_116 = _EVAL_17 == 3'h0;
  assign _EVAL_244 = _EVAL_114 | _EVAL_6;
  assign _EVAL_245 = _EVAL_46 | _EVAL_6;
  assign _EVAL_301 = 2'h1 << _EVAL_8;
  assign _EVAL_162 = _EVAL_254 | _EVAL_147;
  assign _EVAL_137 = _EVAL_265 - 6'h1;
  assign _EVAL_292 = _EVAL & _EVAL_63;
  assign _EVAL_140 = _EVAL_17 == 3'h1;
  assign _EVAL_84 = _EVAL_86 | _EVAL_6;
  assign _EVAL_128 = _EVAL_304 | _EVAL_188;
  assign _EVAL_62 = $signed(_EVAL_95) == 33'sh0;
  assign _EVAL_24 = ~_EVAL_221;
  assign _EVAL_242 = _EVAL_259 == 6'h0;
  assign _EVAL_32 = _EVAL_249 != _EVAL_120;
  assign _EVAL_117 = ~_EVAL_44;
  assign _EVAL_277 = ~_EVAL_52;
  assign _EVAL_205 = _EVAL_9 <= 3'h2;
  assign _EVAL_55 = _EVAL_12 & _EVAL_171;
  assign _EVAL_163 = ~_EVAL_267;
  assign _EVAL_27 = _EVAL_309 | _EVAL_160;
  assign _EVAL_231 = _EVAL_203 >> _EVAL_8;
  assign _EVAL_106 = _EVAL_17 == 3'h5;
  assign _EVAL_88 = $signed(_EVAL_211) == 33'sh0;
  assign _EVAL_221 = _EVAL_217 | _EVAL_6;
  assign _EVAL_48 = ~_EVAL_305;
  assign _EVAL_272 = _EVAL_53 | _EVAL_6;
  assign _EVAL_164 = _EVAL_227 | _EVAL_200;
  assign _EVAL_170 = _EVAL_19 | _EVAL_88;
  assign _EVAL_288 = ~_EVAL_290;
  assign _EVAL_79 = _EVAL_12 & _EVAL_310;
  assign _EVAL_220 = ~_EVAL_239;
  assign _EVAL_206 = _EVAL_208 | _EVAL_161;
  assign _EVAL_275 = ~_EVAL_101;
  assign _EVAL_94 = ~_EVAL_6;
  assign _EVAL_149 = ~_EVAL_209;
  assign _EVAL_21 = ~_EVAL_248;
  assign _EVAL_207 = _EVAL_47 & _EVAL_170;
  assign _EVAL_119 = _EVAL_208 | _EVAL_243;
  assign _EVAL_29 = ~_EVAL_287;
  assign _EVAL_282 = _EVAL_18 == _EVAL_235;
  assign _EVAL_182 = _EVAL_62 | _EVAL_317;
  assign _EVAL_51 = 2'h1 << _EVAL_15;
  assign _EVAL_215 = ~_EVAL_313;
  assign _EVAL_112 = ~_EVAL_54;
  assign _EVAL_319 = _EVAL_142[7:0];
  assign _EVAL_19 = _EVAL_182 | _EVAL_315;
  assign _EVAL_304 = _EVAL_207 | _EVAL_105;
  assign _EVAL_75 = _EVAL_265 == 6'h0;
  assign _EVAL_253 = _EVAL_318[7:2];
  assign _EVAL_74 = _EVAL_1 == _EVAL_158;
  assign _EVAL_130 = _EVAL_257 | _EVAL_6;
  assign _EVAL_81 = ~_EVAL_57;
  assign _EVAL_266 = ~_EVAL_260;
  assign _EVAL_249 = _EVAL_238 ? _EVAL_51 : 2'h0;
  assign _EVAL_300 = _EVAL_5 == 3'h3;
  assign _EVAL_254 = _EVAL_3 & _EVAL_12;
  assign _EVAL_214 = {1'b0,$signed(_EVAL_246)};
  assign _EVAL_42 = _EVAL_278 == 4'h0;
  assign _EVAL_290 = _EVAL_173 | _EVAL_6;
  assign _EVAL_53 = _EVAL_9 == _EVAL_184;
  assign _EVAL_264 = 2'h1 << _EVAL_136;
  assign _EVAL_278 = ~_EVAL;
  assign _EVAL_183 = _EVAL_98 < plusarg_reader_out;
  assign _EVAL_47 = _EVAL_1 <= 4'h2;
  assign _EVAL_165 = _EVAL_102 & _EVAL_266;
  assign _EVAL_151 = _EVAL_11 == _EVAL_276;
  assign _EVAL_188 = _EVAL_97 & _EVAL_34;
  assign _EVAL_295 = _EVAL_14 & _EVAL_222;
  assign _EVAL_109 = _EVAL_199 | _EVAL_6;
  assign _EVAL_45 = _EVAL_254 & _EVAL_293;
  assign _EVAL_187 = _EVAL_17 == _EVAL_311;
  assign _EVAL_318 = ~_EVAL_319;
  assign _EVAL_175 = _EVAL_34 | _EVAL_317;
  assign _EVAL_299 = ~_EVAL_216;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_72 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_78 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_98 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_138 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_150 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_158 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_172 = _RAND_6[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_177 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_184 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_192 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_234 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_235 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_240 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_259 = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_265 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_276 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_311 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_16) begin
    if (_EVAL_45) begin
      _EVAL_72 <= _EVAL_5;
    end
    if (_EVAL_45) begin
      _EVAL_78 <= _EVAL_2;
    end
    if (_EVAL_6) begin
      _EVAL_98 <= 32'h0;
    end else if (_EVAL_162) begin
      _EVAL_98 <= 32'h0;
    end else begin
      _EVAL_98 <= _EVAL_256;
    end
    if (_EVAL_286) begin
      _EVAL_138 <= _EVAL_7;
    end
    if (_EVAL_286) begin
      _EVAL_150 <= _EVAL_8;
    end
    if (_EVAL_45) begin
      _EVAL_158 <= _EVAL_1;
    end
    if (_EVAL_6) begin
      _EVAL_172 <= 6'h0;
    end else if (_EVAL_254) begin
      if (_EVAL_293) begin
        if (_EVAL_220) begin
          _EVAL_172 <= _EVAL_253;
        end else begin
          _EVAL_172 <= 6'h0;
        end
      end else begin
        _EVAL_172 <= _EVAL_110;
      end
    end
    if (_EVAL_6) begin
      _EVAL_177 <= 2'h0;
    end else begin
      _EVAL_177 <= _EVAL_89;
    end
    if (_EVAL_45) begin
      _EVAL_184 <= _EVAL_9;
    end
    if (_EVAL_286) begin
      _EVAL_192 <= _EVAL_10;
    end
    if (_EVAL_6) begin
      _EVAL_234 <= 6'h0;
    end else if (_EVAL_147) begin
      if (_EVAL_312) begin
        if (_EVAL_281) begin
          _EVAL_234 <= _EVAL_202;
        end else begin
          _EVAL_234 <= 6'h0;
        end
      end else begin
        _EVAL_234 <= _EVAL_306;
      end
    end
    if (_EVAL_286) begin
      _EVAL_235 <= _EVAL_18;
    end
    if (_EVAL_45) begin
      _EVAL_240 <= _EVAL_15;
    end
    if (_EVAL_6) begin
      _EVAL_259 <= 6'h0;
    end else if (_EVAL_147) begin
      if (_EVAL_242) begin
        if (_EVAL_281) begin
          _EVAL_259 <= _EVAL_202;
        end else begin
          _EVAL_259 <= 6'h0;
        end
      end else begin
        _EVAL_259 <= _EVAL_37;
      end
    end
    if (_EVAL_6) begin
      _EVAL_265 <= 6'h0;
    end else if (_EVAL_254) begin
      if (_EVAL_75) begin
        if (_EVAL_220) begin
          _EVAL_265 <= _EVAL_253;
        end else begin
          _EVAL_265 <= 6'h0;
        end
      end else begin
        _EVAL_265 <= _EVAL_190;
      end
    end
    if (_EVAL_286) begin
      _EVAL_276 <= _EVAL_11;
    end
    if (_EVAL_286) begin
      _EVAL_311 <= _EVAL_17;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cf83e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_324) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f192b70b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7dc03179)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a2d2b60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_308) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c95356ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_299) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f5e3eec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d31a7aac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86db0dfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bb6bb30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ef594a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7171687)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdc57f02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41701d9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64bb9d58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a668857)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_275) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da52d4a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3edf12e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_308) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(965523e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7f86806)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_308) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2cfcb90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d21b4c75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_324) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(595728b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1ad69e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5609bc4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d31a10f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8481d6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71116efb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_308) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f842a1a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af08ba9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f78791f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e687a695)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5983c0a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa04fbdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_288) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4beb552e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa6faffc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fa2fb1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4f6495f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_324) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b307929)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(501813f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c1dd985)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(342e968)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2f8acb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_324) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66ce2347)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(220938fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6680e4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c14a362)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(432a2b02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eeaaaa73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2515227b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_299) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59bdcbdb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd2f2626)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(977e546b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_299) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4aa871e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f05b4b2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_275) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7c64d30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_322) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd801533)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b2ec15f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e16a5762)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f4d13fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_299) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(960d12d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f5628cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b8550a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ee2b2c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b51a699)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76ff606c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6c4e5b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db311713)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f969b1b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_288) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bc75703)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f67516e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_322) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bebbcc9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77ebe19c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a4e0c32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f220088)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ed212cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86fd1323)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34b6ef46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
