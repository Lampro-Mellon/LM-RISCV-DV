//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_48_assert(
  input         _EVAL,
  input  [31:0] _EVAL_0,
  input         _EVAL_1,
  input  [3:0]  _EVAL_2,
  input  [3:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input  [1:0]  _EVAL_12,
  input         _EVAL_13,
  input  [3:0]  _EVAL_14,
  input         _EVAL_15
);
  wire  _EVAL_16;
  wire  _EVAL_17;
  reg [31:0] _EVAL_18;
  reg [31:0] _RAND_0;
  wire  _EVAL_19;
  reg [1:0] _EVAL_20;
  reg [31:0] _RAND_1;
  wire  _EVAL_21;
  wire [1:0] _EVAL_22;
  reg [3:0] _EVAL_23;
  reg [31:0] _RAND_2;
  wire [32:0] _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  reg [2:0] _EVAL_28;
  reg [31:0] _RAND_3;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire [7:0] _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  reg [5:0] _EVAL_48;
  reg [31:0] _RAND_4;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire [5:0] _EVAL_51;
  wire [1:0] _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire [6:0] _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire [32:0] _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire [32:0] _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire [32:0] _EVAL_94;
  wire [3:0] _EVAL_96;
  wire  _EVAL_97;
  wire [3:0] _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire [31:0] _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire [6:0] _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire [31:0] _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire [1:0] _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  reg [2:0] _EVAL_119;
  reg [31:0] _RAND_5;
  wire  _EVAL_120;
  reg [5:0] _EVAL_121;
  reg [31:0] _RAND_6;
  wire [31:0] _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  reg [31:0] _EVAL_125;
  reg [31:0] _RAND_7;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire [5:0] _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire [3:0] _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire [7:0] _EVAL_142;
  wire  _EVAL_143;
  wire [32:0] _EVAL_144;
  wire [31:0] _EVAL_145;
  wire  _EVAL_146;
  wire [31:0] _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  reg  _EVAL_153;
  reg [31:0] _RAND_8;
  wire [32:0] _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire [6:0] _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire [5:0] _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire [32:0] _EVAL_168;
  wire  _EVAL_169;
  wire [22:0] _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  reg [5:0] _EVAL_173;
  reg [31:0] _RAND_9;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  reg  _EVAL_188;
  reg [31:0] _RAND_10;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire [32:0] _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire [7:0] _EVAL_197;
  wire [3:0] _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire [22:0] _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  reg  _EVAL_209;
  reg [31:0] _RAND_11;
  wire [31:0] plusarg_reader_out;
  wire [5:0] _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire [32:0] _EVAL_213;
  wire  _EVAL_214;
  wire [32:0] _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire [32:0] _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire [31:0] _EVAL_227;
  wire [5:0] _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire [1:0] _EVAL_234;
  wire [32:0] _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire [32:0] _EVAL_239;
  wire [32:0] _EVAL_240;
  wire  _EVAL_241;
  wire [32:0] _EVAL_242;
  wire  _EVAL_243;
  reg [3:0] _EVAL_244;
  reg [31:0] _RAND_12;
  wire [6:0] _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire [5:0] _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire [31:0] _EVAL_254;
  wire [32:0] _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_260;
  wire [32:0] _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire [32:0] _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire [7:0] _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  reg [5:0] _EVAL_277;
  reg [31:0] _RAND_13;
  wire  _EVAL_278;
  wire [31:0] _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire [1:0] _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire [32:0] _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  reg  _EVAL_290;
  reg [31:0] _RAND_14;
  wire  _EVAL_291;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_147 = _EVAL_0 ^ 32'h40000000;
  assign _EVAL_97 = _EVAL_7[0];
  assign _EVAL_251 = _EVAL_36 | _EVAL_6;
  assign _EVAL_85 = _EVAL_53 | _EVAL_6;
  assign _EVAL_24 = {1'b0,$signed(_EVAL_0)};
  assign _EVAL_118 = _EVAL_12 != 2'h2;
  assign _EVAL_51 = _EVAL_245[5:0];
  assign _EVAL_114 = _EVAL_136 | _EVAL_6;
  assign _EVAL_57 = _EVAL_181 | _EVAL_195;
  assign _EVAL_49 = _EVAL_14 <= 4'h2;
  assign _EVAL_229 = _EVAL_10 == 3'h1;
  assign _EVAL_112 = _EVAL_173 == 6'h0;
  assign _EVAL_102 = _EVAL_7 <= 3'h6;
  assign _EVAL_45 = _EVAL_14[0];
  assign _EVAL_177 = _EVAL_134 == 4'h0;
  assign _EVAL_101 = _EVAL_0 ^ 32'h80000000;
  assign _EVAL_134 = _EVAL_2 & _EVAL_98;
  assign _EVAL_216 = _EVAL_137 & _EVAL_149;
  assign _EVAL_246 = ~_EVAL_131;
  assign _EVAL_89 = _EVAL_128 | _EVAL_190;
  assign _EVAL_215 = $signed(_EVAL_144) & -33'sh2000;
  assign _EVAL_136 = _EVAL == _EVAL_290;
  assign _EVAL_38 = ~_EVAL_107;
  assign _EVAL_226 = _EVAL_138 & _EVAL_224;
  assign _EVAL_162 = _EVAL_173 - 6'h1;
  assign _EVAL_35 = _EVAL_283 | _EVAL_6;
  assign _EVAL_267 = _EVAL_49 & _EVAL_217;
  assign _EVAL_124 = ~_EVAL_149;
  assign _EVAL_74 = _EVAL_18 < plusarg_reader_out;
  assign _EVAL_62 = ~_EVAL_85;
  assign _EVAL_183 = _EVAL_12 <= 2'h2;
  assign _EVAL_80 = _EVAL_10 == 3'h3;
  assign _EVAL_59 = _EVAL_48 == 6'h0;
  assign _EVAL_143 = ~_EVAL_260;
  assign _EVAL_240 = {1'b0,$signed(_EVAL_122)};
  assign _EVAL_144 = {1'b0,$signed(_EVAL_145)};
  assign _EVAL_65 = _EVAL_121 == 6'h0;
  assign _EVAL_108 = ~_EVAL_47;
  assign _EVAL_63 = _EVAL_127 | _EVAL_6;
  assign _EVAL_43 = _EVAL_87 | _EVAL_6;
  assign _EVAL_60 = _EVAL_25 >> _EVAL_5;
  assign _EVAL_148 = _EVAL_17 | _EVAL_6;
  assign _EVAL_99 = _EVAL_7 == 3'h4;
  assign _EVAL_189 = ~_EVAL_15;
  assign _EVAL_73 = _EVAL_242;
  assign _EVAL_105 = $signed(_EVAL_255) == 33'sh0;
  assign _EVAL_92 = _EVAL_183 | _EVAL_6;
  assign _EVAL_137 = _EVAL_1 & _EVAL_13;
  assign _EVAL_67 = _EVAL_121 - 6'h1;
  assign _EVAL_207 = _EVAL_7 == 3'h1;
  assign _EVAL_150 = _EVAL_141 & _EVAL_250;
  assign _EVAL_174 = _EVAL_123 | _EVAL_226;
  assign _EVAL_122 = _EVAL_0 ^ 32'h3000;
  assign _EVAL_90 = _EVAL_60 | _EVAL_6;
  assign _EVAL_131 = _EVAL_238 | _EVAL_6;
  assign _EVAL_171 = ~_EVAL_75;
  assign _EVAL_53 = _EVAL_15 == _EVAL_209;
  assign _EVAL_227 = _EVAL_79[31:0];
  assign _EVAL_224 = _EVAL_175 & _EVAL_275;
  assign _EVAL_31 = _EVAL_137 & _EVAL_65;
  assign _EVAL_287 = _EVAL_50 | _EVAL_74;
  assign _EVAL_279 = _EVAL_0 & _EVAL_254;
  assign _EVAL_116 = _EVAL_89 | _EVAL_100;
  assign _EVAL_130 = ~_EVAL_249;
  assign _EVAL_120 = ~_EVAL_140;
  assign _EVAL_86 = ~_EVAL_188;
  assign _EVAL_286 = $signed(_EVAL_24) & -33'sh5000;
  assign _EVAL_40 = _EVAL_30 | _EVAL_190;
  assign _EVAL_206 = ~_EVAL_271;
  assign _EVAL_26 = _EVAL_9 & _EVAL_237;
  assign _EVAL_280 = _EVAL_82 | _EVAL_6;
  assign _EVAL_164 = ~_EVAL_288;
  assign _EVAL_235 = _EVAL_261;
  assign _EVAL_157 = _EVAL_7 == 3'h5;
  assign _EVAL_257 = _EVAL_14 <= 4'h8;
  assign _EVAL_167 = _EVAL_7 == 3'h6;
  assign _EVAL_140 = _EVAL_113 | _EVAL_6;
  assign _EVAL_236 = _EVAL_123 | _EVAL_172;
  assign _EVAL_203 = 23'hff << _EVAL_3;
  assign _EVAL_273 = ~_EVAL_220;
  assign _EVAL_250 = ~_EVAL_175;
  assign _EVAL_276 = _EVAL_250 & _EVAL_275;
  assign _EVAL_195 = _EVAL_49 & _EVAL_100;
  assign _EVAL_255 = _EVAL_94;
  assign _EVAL_109 = _EVAL_0 ^ 32'h2000000;
  assign _EVAL_193 = _EVAL_10 == 3'h0;
  assign _EVAL_222 = _EVAL_154;
  assign _EVAL_249 = _EVAL_70 | _EVAL_6;
  assign _EVAL_248 = _EVAL_67[5:0];
  assign _EVAL_243 = _EVAL_14 >= 4'h2;
  assign _EVAL_239 = {1'b0,$signed(_EVAL_109)};
  assign _EVAL_104 = _EVAL_277 - 6'h1;
  assign _EVAL_234 = 2'h1 << _EVAL_5;
  assign _EVAL_230 = _EVAL_13 & _EVAL_229;
  assign _EVAL_37 = _EVAL_49 & _EVAL_40;
  assign _EVAL_154 = $signed(_EVAL_240) & -33'sh1000;
  assign _EVAL_245 = _EVAL_48 - 6'h1;
  assign _EVAL_79 = _EVAL_18 + 32'h1;
  assign _EVAL_289 = _EVAL_188 | _EVAL_166;
  assign _EVAL_211 = _EVAL_10 == 3'h7;
  assign _EVAL_187 = _EVAL_257 & _EVAL_111;
  assign _EVAL_94 = $signed(_EVAL_213) & -33'sh2000;
  assign _EVAL_68 = ~_EVAL_35;
  assign _EVAL_254 = {{24'd0}, _EVAL_272};
  assign _EVAL_16 = _EVAL_10 == _EVAL_119;
  assign _EVAL_100 = $signed(_EVAL_168) == 33'sh0;
  assign _EVAL_242 = $signed(_EVAL_191) & -33'shc000;
  assign _EVAL_128 = _EVAL_111 | _EVAL_265;
  assign _EVAL_194 = ~_EVAL_5;
  assign _EVAL_221 = ~_EVAL_205;
  assign _EVAL_264 = _EVAL_8 & _EVAL_9;
  assign _EVAL_271 = _EVAL_256 | _EVAL_6;
  assign _EVAL_50 = _EVAL_86 | _EVAL_155;
  assign _EVAL_252 = ~_EVAL_114;
  assign _EVAL_30 = _EVAL_93 | _EVAL_265;
  assign _EVAL_285 = _EVAL_138 & _EVAL_103;
  assign _EVAL_237 = ~_EVAL_59;
  assign _EVAL_232 = _EVAL_9 & _EVAL_207;
  assign _EVAL_253 = ~_EVAL_92;
  assign _EVAL_161 = _EVAL_141 & _EVAL_175;
  assign _EVAL_179 = _EVAL_58 & _EVAL_105;
  assign _EVAL_212 = ~_EVAL_90;
  assign _EVAL_225 = _EVAL_284 & _EVAL_231;
  assign _EVAL_214 = _EVAL_86 | _EVAL_6;
  assign _EVAL_54 = _EVAL_267 | _EVAL_179;
  assign _EVAL_159 = _EVAL_189 | _EVAL_11;
  assign _EVAL_247 = _EVAL_12 == 2'h0;
  assign _EVAL_58 = _EVAL_14 <= 4'h6;
  assign _EVAL_272 = ~_EVAL_142;
  assign _EVAL_82 = _EVAL_279 == 32'h0;
  assign _EVAL_127 = _EVAL_12 == _EVAL_20;
  assign _EVAL_233 = _EVAL_243 | _EVAL_150;
  assign _EVAL_208 = _EVAL_9 & _EVAL_99;
  assign _EVAL_284 = _EVAL_264 & _EVAL_112;
  assign _EVAL_69 = _EVAL_13 & _EVAL_124;
  assign _EVAL_160 = ~_EVAL_6;
  assign _EVAL_138 = _EVAL_22[0];
  assign _EVAL_64 = _EVAL_189 | _EVAL_6;
  assign _EVAL_77 = _EVAL_13 & _EVAL_193;
  assign _EVAL_172 = _EVAL_138 & _EVAL_56;
  assign _EVAL_17 = _EVAL_3 == _EVAL_244;
  assign _EVAL_32 = ~_EVAL_197;
  assign _EVAL_149 = _EVAL_277 == 6'h0;
  assign _EVAL_141 = _EVAL_22[1];
  assign _EVAL_241 = _EVAL_13 & _EVAL_270;
  assign _EVAL_204 = _EVAL_0 == _EVAL_125;
  assign _EVAL_182 = _EVAL_13 & _EVAL_211;
  assign _EVAL_123 = _EVAL_243 | _EVAL_161;
  assign _EVAL_70 = _EVAL_5 == _EVAL_153;
  assign _EVAL_181 = _EVAL_179 | _EVAL_187;
  assign _EVAL_76 = ~_EVAL_43;
  assign _EVAL_168 = _EVAL_215;
  assign _EVAL_110 = _EVAL_37 | _EVAL_187;
  assign _EVAL_185 = _EVAL_166 != _EVAL_169;
  assign _EVAL_258 = ~_EVAL_63;
  assign _EVAL_42 = _EVAL_118 | _EVAL_6;
  assign _EVAL_200 = _EVAL_9 & _EVAL_126;
  assign _EVAL_135 = _EVAL_243 | _EVAL_6;
  assign _EVAL_288 = _EVAL_16 | _EVAL_6;
  assign _EVAL_111 = $signed(_EVAL_222) == 33'sh0;
  assign _EVAL_145 = _EVAL_0 ^ 32'h20000000;
  assign _EVAL_165 = _EVAL_162[5:0];
  assign _EVAL_33 = _EVAL_233 | _EVAL_285;
  assign _EVAL_202 = _EVAL_264 & _EVAL_59;
  assign _EVAL_274 = _EVAL_10[2];
  assign _EVAL_199 = _EVAL_13 & _EVAL_21;
  assign _EVAL_55 = _EVAL_233 | _EVAL_176;
  assign _EVAL_146 = ~_EVAL_291;
  assign _EVAL_220 = _EVAL_177 | _EVAL_6;
  assign _EVAL_81 = _EVAL_10 == 3'h6;
  assign _EVAL_166 = _EVAL_52[0];
  assign _EVAL_282 = _EVAL_225 ? _EVAL_234 : 2'h0;
  assign _EVAL_197 = _EVAL_203[7:0];
  assign _EVAL_269 = _EVAL_286;
  assign _EVAL_44 = _EVAL_156 | _EVAL_6;
  assign _EVAL_129 = _EVAL_32[7:2];
  assign _EVAL_186 = _EVAL_13 & _EVAL_80;
  assign _EVAL_83 = ~_EVAL_280;
  assign _EVAL_231 = ~_EVAL_167;
  assign _EVAL_34 = ~_EVAL_275;
  assign _EVAL_163 = ~_EVAL_214;
  assign _EVAL_126 = _EVAL_7 == 3'h0;
  assign _EVAL_184 = ~_EVAL_42;
  assign _EVAL_238 = ~_EVAL_11;
  assign _EVAL_87 = _EVAL_2 == _EVAL_96;
  assign _EVAL_19 = ~_EVAL_135;
  assign _EVAL_278 = _EVAL_247 | _EVAL_6;
  assign _EVAL_142 = _EVAL_170[7:0];
  assign _EVAL_263 = ~_EVAL_251;
  assign _EVAL_291 = _EVAL_204 | _EVAL_6;
  assign _EVAL_210 = _EVAL_104[5:0];
  assign _EVAL_93 = $signed(_EVAL_73) == 33'sh0;
  assign _EVAL_132 = _EVAL_7 == 3'h2;
  assign _EVAL_223 = ~_EVAL_169;
  assign _EVAL_228 = _EVAL_272[7:2];
  assign _EVAL_133 = ~_EVAL_274;
  assign _EVAL_201 = _EVAL_72 | _EVAL_6;
  assign _EVAL_117 = ~_EVAL_166;
  assign _EVAL_115 = 2'h1 << _EVAL_45;
  assign _EVAL_61 = _EVAL_39 | _EVAL_6;
  assign _EVAL_213 = {1'b0,$signed(_EVAL_147)};
  assign _EVAL_261 = $signed(_EVAL_239) & -33'sh1000000;
  assign _EVAL_262 = _EVAL_137 | _EVAL_264;
  assign _EVAL_56 = _EVAL_175 & _EVAL_34;
  assign _EVAL_283 = _EVAL_14 == _EVAL_23;
  assign _EVAL_98 = ~_EVAL_96;
  assign _EVAL_107 = _EVAL_110 | _EVAL_6;
  assign _EVAL_191 = {1'b0,$signed(_EVAL_101)};
  assign _EVAL_218 = ~_EVAL_278;
  assign _EVAL_205 = _EVAL_102 | _EVAL_6;
  assign _EVAL_21 = _EVAL_10 == 3'h5;
  assign _EVAL_270 = _EVAL_10 == 3'h2;
  assign _EVAL_281 = ~_EVAL_61;
  assign _EVAL_36 = _EVAL_49 & _EVAL_116;
  assign _EVAL_139 = _EVAL_9 & _EVAL_132;
  assign _EVAL_66 = _EVAL_13 & _EVAL_84;
  assign _EVAL_219 = _EVAL_57 | _EVAL_6;
  assign _EVAL_52 = _EVAL_31 ? 2'h1 : 2'h0;
  assign _EVAL_198 = ~_EVAL_2;
  assign _EVAL_25 = _EVAL_166 | _EVAL_188;
  assign _EVAL_96 = {_EVAL_174,_EVAL_236,_EVAL_55,_EVAL_33};
  assign _EVAL_217 = _EVAL_40 | _EVAL_100;
  assign _EVAL_39 = _EVAL_7 == _EVAL_28;
  assign _EVAL_22 = _EVAL_115 | 2'h1;
  assign _EVAL_260 = _EVAL_194 | _EVAL_6;
  assign _EVAL_84 = _EVAL_10 == 3'h4;
  assign _EVAL_41 = ~_EVAL_219;
  assign _EVAL_178 = ~_EVAL_148;
  assign _EVAL_156 = _EVAL_185 | _EVAL_117;
  assign _EVAL_192 = ~_EVAL_201;
  assign _EVAL_275 = _EVAL_0[0];
  assign _EVAL_180 = _EVAL_9 & _EVAL_157;
  assign _EVAL_46 = _EVAL_9 & _EVAL_167;
  assign _EVAL_196 = _EVAL_289 & _EVAL_223;
  assign _EVAL_75 = _EVAL_287 | _EVAL_6;
  assign _EVAL_155 = plusarg_reader_out == 32'h0;
  assign _EVAL_175 = _EVAL_0[1];
  assign _EVAL_176 = _EVAL_138 & _EVAL_276;
  assign _EVAL_113 = _EVAL_198 == 4'h0;
  assign _EVAL_47 = _EVAL_159 | _EVAL_6;
  assign _EVAL_103 = _EVAL_250 & _EVAL_34;
  assign _EVAL_266 = ~_EVAL_64;
  assign _EVAL_170 = 23'hff << _EVAL_14;
  assign _EVAL_71 = ~_EVAL_44;
  assign _EVAL_169 = _EVAL_282[0];
  assign _EVAL_190 = $signed(_EVAL_269) == 33'sh0;
  assign _EVAL_72 = _EVAL_54 | _EVAL_187;
  assign _EVAL_256 = _EVAL_3 >= 4'h2;
  assign _EVAL_91 = _EVAL_13 & _EVAL_81;
  assign _EVAL_265 = $signed(_EVAL_235) == 33'sh0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_18 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_20 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_23 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_28 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_48 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_119 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_121 = _RAND_6[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_125 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_153 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_173 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_188 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_209 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_244 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_277 = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_290 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_4) begin
    if (_EVAL_6) begin
      _EVAL_18 <= 32'h0;
    end else if (_EVAL_262) begin
      _EVAL_18 <= 32'h0;
    end else begin
      _EVAL_18 <= _EVAL_227;
    end
    if (_EVAL_202) begin
      _EVAL_20 <= _EVAL_12;
    end
    if (_EVAL_216) begin
      _EVAL_23 <= _EVAL_14;
    end
    if (_EVAL_202) begin
      _EVAL_28 <= _EVAL_7;
    end
    if (_EVAL_6) begin
      _EVAL_48 <= 6'h0;
    end else if (_EVAL_264) begin
      if (_EVAL_59) begin
        if (_EVAL_97) begin
          _EVAL_48 <= _EVAL_129;
        end else begin
          _EVAL_48 <= 6'h0;
        end
      end else begin
        _EVAL_48 <= _EVAL_51;
      end
    end
    if (_EVAL_216) begin
      _EVAL_119 <= _EVAL_10;
    end
    if (_EVAL_6) begin
      _EVAL_121 <= 6'h0;
    end else if (_EVAL_137) begin
      if (_EVAL_65) begin
        if (_EVAL_133) begin
          _EVAL_121 <= _EVAL_228;
        end else begin
          _EVAL_121 <= 6'h0;
        end
      end else begin
        _EVAL_121 <= _EVAL_248;
      end
    end
    if (_EVAL_216) begin
      _EVAL_125 <= _EVAL_0;
    end
    if (_EVAL_202) begin
      _EVAL_153 <= _EVAL_5;
    end
    if (_EVAL_6) begin
      _EVAL_173 <= 6'h0;
    end else if (_EVAL_264) begin
      if (_EVAL_112) begin
        if (_EVAL_97) begin
          _EVAL_173 <= _EVAL_129;
        end else begin
          _EVAL_173 <= 6'h0;
        end
      end else begin
        _EVAL_173 <= _EVAL_165;
      end
    end
    if (_EVAL_6) begin
      _EVAL_188 <= 1'h0;
    end else begin
      _EVAL_188 <= _EVAL_196;
    end
    if (_EVAL_202) begin
      _EVAL_209 <= _EVAL_15;
    end
    if (_EVAL_202) begin
      _EVAL_244 <= _EVAL_3;
    end
    if (_EVAL_6) begin
      _EVAL_277 <= 6'h0;
    end else if (_EVAL_137) begin
      if (_EVAL_149) begin
        if (_EVAL_133) begin
          _EVAL_277 <= _EVAL_228;
        end else begin
          _EVAL_277 <= 6'h0;
        end
      end else begin
        _EVAL_277 <= _EVAL_210;
      end
    end
    if (_EVAL_202) begin
      _EVAL_290 <= _EVAL;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(476aaeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fbcc887)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cccf737a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89fb1a31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c651f444)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff8c6e60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4343d68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e2076cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31c54afe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c48e4b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9707cfce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1b282ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d9a9bab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd88a06b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a092a7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a8f04d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbe82c8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f472a9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17ded2ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78eed859)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d80e5b60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c54d4dff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c453dae9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de664525)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9467647)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61de9819)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4822e930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc49096f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6e083b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2745ea79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bd7ca9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f18c15d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bba0d9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5da3a832)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6403b68a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38c2f2ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7dd908d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(513aedb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42da7f7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bec3b726)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98523ede)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7e73e6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa236aba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf63551c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d261ecc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d6e8fd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24d0773d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fa14966)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b579320e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4531ea97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2175f1cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad9fd30c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(811987fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b755fd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c220aaf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e31a331)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bbd1c78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53df6ac1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be6846aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19fa1ad6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(692d37e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef44954)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a854b0ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33d27c11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1edcd4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78134d0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8c06efa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5e6264d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(476d920b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
