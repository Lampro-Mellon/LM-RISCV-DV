//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_136(
  output        _EVAL,
  output [8:0]  _EVAL_0,
  input  [6:0]  _EVAL_1,
  input  [31:0] _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  output [2:0]  _EVAL_5,
  output        _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  output        _EVAL_12,
  input  [31:0] _EVAL_13,
  output        _EVAL_14,
  output        _EVAL_15,
  output        _EVAL_16,
  input  [1:0]  _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19,
  output        _EVAL_20,
  output [3:0]  _EVAL_21,
  output        _EVAL_22,
  output        _EVAL_23,
  input         _EVAL_24,
  output [1:0]  _EVAL_25,
  output        _EVAL_26,
  input         _EVAL_27,
  output [31:0] _EVAL_28,
  input  [1:0]  _EVAL_29,
  output [31:0] _EVAL_30,
  input         _EVAL_31
);
  wire  _EVAL_32;
  wire [2:0] asource__EVAL;
  wire [8:0] asource__EVAL_0;
  wire [31:0] asource__EVAL_1;
  wire  asource__EVAL_2;
  wire  asource__EVAL_3;
  wire [8:0] asource__EVAL_4;
  wire [31:0] asource__EVAL_5;
  wire  asource__EVAL_6;
  wire  asource__EVAL_7;
  wire  asource__EVAL_8;
  wire  asource__EVAL_9;
  wire [1:0] asource__EVAL_10;
  wire [2:0] asource__EVAL_11;
  wire  asource__EVAL_12;
  wire  asource__EVAL_13;
  wire  asource__EVAL_14;
  wire [3:0] asource__EVAL_15;
  wire  asource__EVAL_16;
  wire [31:0] asource__EVAL_17;
  wire  asource__EVAL_18;
  wire [31:0] asource__EVAL_19;
  wire [1:0] asource__EVAL_20;
  wire [3:0] asource__EVAL_21;
  wire [2:0] asource__EVAL_22;
  wire [1:0] asource__EVAL_23;
  wire  asource__EVAL_24;
  wire [2:0] asource__EVAL_25;
  wire  asource__EVAL_26;
  wire  asource__EVAL_27;
  wire  asource__EVAL_28;
  wire  AsyncQueueSource__EVAL;
  wire  AsyncQueueSource__EVAL_0;
  wire  AsyncQueueSource__EVAL_1;
  wire  AsyncQueueSource__EVAL_2;
  wire  AsyncQueueSource__EVAL_3;
  wire  AsyncQueueSource__EVAL_4;
  wire  AsyncQueueSource__EVAL_5;
  wire  AsyncQueueSource__EVAL_6;
  wire  AsyncQueueSource__EVAL_7;
  wire  AsyncQueueSource__EVAL_8;
  wire  AsyncQueueSource__EVAL_9;
  wire  AsyncQueueSource__EVAL_10;
  wire [2:0] dmiXbar__EVAL;
  wire [31:0] dmiXbar__EVAL_0;
  wire  dmiXbar__EVAL_1;
  wire [3:0] dmiXbar__EVAL_2;
  wire  dmiXbar__EVAL_3;
  wire [31:0] dmiXbar__EVAL_4;
  wire [31:0] dmiXbar__EVAL_5;
  wire [2:0] dmiXbar__EVAL_6;
  wire [3:0] dmiXbar__EVAL_7;
  wire  dmiXbar__EVAL_8;
  wire  dmiXbar__EVAL_9;
  wire [2:0] dmiXbar__EVAL_10;
  wire  dmiXbar__EVAL_11;
  wire [8:0] dmiXbar__EVAL_12;
  wire  dmiXbar__EVAL_13;
  wire  dmiXbar__EVAL_14;
  wire  dmiXbar__EVAL_15;
  wire  dmiXbar__EVAL_16;
  wire [1:0] dmiXbar__EVAL_17;
  wire [31:0] dmiXbar__EVAL_18;
  wire [1:0] dmiXbar__EVAL_19;
  wire  dmiXbar__EVAL_20;
  wire  dmiXbar__EVAL_21;
  wire [8:0] dmiXbar__EVAL_22;
  wire [31:0] dmiXbar__EVAL_23;
  wire [3:0] dmiXbar__EVAL_24;
  wire  dmiXbar__EVAL_25;
  wire  dmiXbar__EVAL_26;
  wire [2:0] dmiXbar__EVAL_27;
  wire  dmiXbar__EVAL_28;
  wire  dmiXbar__EVAL_29;
  wire [2:0] dmiXbar__EVAL_30;
  wire  dmiXbar__EVAL_31;
  wire  dmiXbar__EVAL_32;
  wire  dmiXbar__EVAL_33;
  wire  dmiXbar__EVAL_34;
  wire [31:0] dmiXbar__EVAL_35;
  wire [6:0] dmiXbar__EVAL_36;
  wire  dmiXbar__EVAL_37;
  wire  dmactiveAckSync__EVAL;
  wire  dmactiveAckSync__EVAL_0;
  wire  dmactiveAckSync__EVAL_1;
  wire  dmactiveAckSync__EVAL_2;
  wire [31:0] dmOuter__EVAL;
  wire [31:0] dmOuter__EVAL_0;
  wire [6:0] dmOuter__EVAL_1;
  wire  dmOuter__EVAL_2;
  wire  dmOuter__EVAL_3;
  wire  dmOuter__EVAL_4;
  wire  dmOuter__EVAL_5;
  wire  dmOuter__EVAL_6;
  wire  dmOuter__EVAL_7;
  wire  dmOuter__EVAL_8;
  wire  dmOuter__EVAL_9;
  wire  dmOuter__EVAL_10;
  wire [2:0] dmOuter__EVAL_11;
  wire  dmOuter__EVAL_12;
  wire  dmOuter__EVAL_13;
  wire  dmOuter__EVAL_14;
  wire  dmOuter__EVAL_15;
  wire [2:0] dmOuter__EVAL_16;
  wire  dmOuter__EVAL_17;
  wire  dmOuter__EVAL_18;
  wire  dmOuter__EVAL_19;
  wire [3:0] dmOuter__EVAL_20;
  wire [9:0] dmOuter__EVAL_21;
  wire  intsource__EVAL;
  wire  intsource__EVAL_0;
  wire  _EVAL_33;
  wire  dmi2tl__EVAL;
  wire [6:0] dmi2tl__EVAL_0;
  wire  dmi2tl__EVAL_1;
  wire  dmi2tl__EVAL_2;
  wire [31:0] dmi2tl__EVAL_3;
  wire  dmi2tl__EVAL_4;
  wire [1:0] dmi2tl__EVAL_5;
  wire [2:0] dmi2tl__EVAL_6;
  wire [31:0] dmi2tl__EVAL_7;
  wire  dmi2tl__EVAL_8;
  wire  dmi2tl__EVAL_9;
  wire [31:0] dmi2tl__EVAL_10;
  wire  dmi2tl__EVAL_11;
  wire  dmi2tl__EVAL_12;
  wire [31:0] dmi2tl__EVAL_13;
  wire [3:0] dmi2tl__EVAL_14;
  wire  dmi2tl__EVAL_15;
  wire  dmi2tl__EVAL_16;
  wire [8:0] dmi2tl__EVAL_17;
  wire [1:0] dmi2tl__EVAL_18;
  wire  _EVAL_34;
  wire  dmiBypass__EVAL;
  wire [3:0] dmiBypass__EVAL_0;
  wire [2:0] dmiBypass__EVAL_1;
  wire [2:0] dmiBypass__EVAL_2;
  wire [1:0] dmiBypass__EVAL_3;
  wire  dmiBypass__EVAL_4;
  wire [1:0] dmiBypass__EVAL_5;
  wire  dmiBypass__EVAL_6;
  wire  dmiBypass__EVAL_7;
  wire  dmiBypass__EVAL_8;
  wire  dmiBypass__EVAL_9;
  wire  dmiBypass__EVAL_10;
  wire [1:0] dmiBypass__EVAL_11;
  wire [31:0] dmiBypass__EVAL_12;
  wire [31:0] dmiBypass__EVAL_13;
  wire [2:0] dmiBypass__EVAL_14;
  wire  dmiBypass__EVAL_15;
  wire [2:0] dmiBypass__EVAL_16;
  wire [31:0] dmiBypass__EVAL_17;
  wire [8:0] dmiBypass__EVAL_18;
  wire [31:0] dmiBypass__EVAL_19;
  wire  dmiBypass__EVAL_20;
  wire  dmiBypass__EVAL_21;
  wire  dmiBypass__EVAL_22;
  wire  dmiBypass__EVAL_23;
  wire  dmiBypass__EVAL_24;
  wire  dmiBypass__EVAL_25;
  wire  dmiBypass__EVAL_26;
  wire [1:0] dmiBypass__EVAL_27;
  wire  dmiBypass__EVAL_28;
  wire  dmiBypass__EVAL_29;
  wire [3:0] dmiBypass__EVAL_30;
  wire [8:0] dmiBypass__EVAL_31;
  wire  dmiBypass__EVAL_32;
  wire  dmiBypass__EVAL_33;
  _EVAL_134 asource (
    ._EVAL(asource__EVAL),
    ._EVAL_0(asource__EVAL_0),
    ._EVAL_1(asource__EVAL_1),
    ._EVAL_2(asource__EVAL_2),
    ._EVAL_3(asource__EVAL_3),
    ._EVAL_4(asource__EVAL_4),
    ._EVAL_5(asource__EVAL_5),
    ._EVAL_6(asource__EVAL_6),
    ._EVAL_7(asource__EVAL_7),
    ._EVAL_8(asource__EVAL_8),
    ._EVAL_9(asource__EVAL_9),
    ._EVAL_10(asource__EVAL_10),
    ._EVAL_11(asource__EVAL_11),
    ._EVAL_12(asource__EVAL_12),
    ._EVAL_13(asource__EVAL_13),
    ._EVAL_14(asource__EVAL_14),
    ._EVAL_15(asource__EVAL_15),
    ._EVAL_16(asource__EVAL_16),
    ._EVAL_17(asource__EVAL_17),
    ._EVAL_18(asource__EVAL_18),
    ._EVAL_19(asource__EVAL_19),
    ._EVAL_20(asource__EVAL_20),
    ._EVAL_21(asource__EVAL_21),
    ._EVAL_22(asource__EVAL_22),
    ._EVAL_23(asource__EVAL_23),
    ._EVAL_24(asource__EVAL_24),
    ._EVAL_25(asource__EVAL_25),
    ._EVAL_26(asource__EVAL_26),
    ._EVAL_27(asource__EVAL_27),
    ._EVAL_28(asource__EVAL_28)
  );
  _EVAL_135 AsyncQueueSource (
    ._EVAL(AsyncQueueSource__EVAL),
    ._EVAL_0(AsyncQueueSource__EVAL_0),
    ._EVAL_1(AsyncQueueSource__EVAL_1),
    ._EVAL_2(AsyncQueueSource__EVAL_2),
    ._EVAL_3(AsyncQueueSource__EVAL_3),
    ._EVAL_4(AsyncQueueSource__EVAL_4),
    ._EVAL_5(AsyncQueueSource__EVAL_5),
    ._EVAL_6(AsyncQueueSource__EVAL_6),
    ._EVAL_7(AsyncQueueSource__EVAL_7),
    ._EVAL_8(AsyncQueueSource__EVAL_8),
    ._EVAL_9(AsyncQueueSource__EVAL_9),
    ._EVAL_10(AsyncQueueSource__EVAL_10)
  );
  _EVAL_118 dmiXbar (
    ._EVAL(dmiXbar__EVAL),
    ._EVAL_0(dmiXbar__EVAL_0),
    ._EVAL_1(dmiXbar__EVAL_1),
    ._EVAL_2(dmiXbar__EVAL_2),
    ._EVAL_3(dmiXbar__EVAL_3),
    ._EVAL_4(dmiXbar__EVAL_4),
    ._EVAL_5(dmiXbar__EVAL_5),
    ._EVAL_6(dmiXbar__EVAL_6),
    ._EVAL_7(dmiXbar__EVAL_7),
    ._EVAL_8(dmiXbar__EVAL_8),
    ._EVAL_9(dmiXbar__EVAL_9),
    ._EVAL_10(dmiXbar__EVAL_10),
    ._EVAL_11(dmiXbar__EVAL_11),
    ._EVAL_12(dmiXbar__EVAL_12),
    ._EVAL_13(dmiXbar__EVAL_13),
    ._EVAL_14(dmiXbar__EVAL_14),
    ._EVAL_15(dmiXbar__EVAL_15),
    ._EVAL_16(dmiXbar__EVAL_16),
    ._EVAL_17(dmiXbar__EVAL_17),
    ._EVAL_18(dmiXbar__EVAL_18),
    ._EVAL_19(dmiXbar__EVAL_19),
    ._EVAL_20(dmiXbar__EVAL_20),
    ._EVAL_21(dmiXbar__EVAL_21),
    ._EVAL_22(dmiXbar__EVAL_22),
    ._EVAL_23(dmiXbar__EVAL_23),
    ._EVAL_24(dmiXbar__EVAL_24),
    ._EVAL_25(dmiXbar__EVAL_25),
    ._EVAL_26(dmiXbar__EVAL_26),
    ._EVAL_27(dmiXbar__EVAL_27),
    ._EVAL_28(dmiXbar__EVAL_28),
    ._EVAL_29(dmiXbar__EVAL_29),
    ._EVAL_30(dmiXbar__EVAL_30),
    ._EVAL_31(dmiXbar__EVAL_31),
    ._EVAL_32(dmiXbar__EVAL_32),
    ._EVAL_33(dmiXbar__EVAL_33),
    ._EVAL_34(dmiXbar__EVAL_34),
    ._EVAL_35(dmiXbar__EVAL_35),
    ._EVAL_36(dmiXbar__EVAL_36),
    ._EVAL_37(dmiXbar__EVAL_37)
  );
  _EVAL_130 dmactiveAckSync (
    ._EVAL(dmactiveAckSync__EVAL),
    ._EVAL_0(dmactiveAckSync__EVAL_0),
    ._EVAL_1(dmactiveAckSync__EVAL_1),
    ._EVAL_2(dmactiveAckSync__EVAL_2)
  );
  _EVAL_121 dmOuter (
    ._EVAL(dmOuter__EVAL),
    ._EVAL_0(dmOuter__EVAL_0),
    ._EVAL_1(dmOuter__EVAL_1),
    ._EVAL_2(dmOuter__EVAL_2),
    ._EVAL_3(dmOuter__EVAL_3),
    ._EVAL_4(dmOuter__EVAL_4),
    ._EVAL_5(dmOuter__EVAL_5),
    ._EVAL_6(dmOuter__EVAL_6),
    ._EVAL_7(dmOuter__EVAL_7),
    ._EVAL_8(dmOuter__EVAL_8),
    ._EVAL_9(dmOuter__EVAL_9),
    ._EVAL_10(dmOuter__EVAL_10),
    ._EVAL_11(dmOuter__EVAL_11),
    ._EVAL_12(dmOuter__EVAL_12),
    ._EVAL_13(dmOuter__EVAL_13),
    ._EVAL_14(dmOuter__EVAL_14),
    ._EVAL_15(dmOuter__EVAL_15),
    ._EVAL_16(dmOuter__EVAL_16),
    ._EVAL_17(dmOuter__EVAL_17),
    ._EVAL_18(dmOuter__EVAL_18),
    ._EVAL_19(dmOuter__EVAL_19),
    ._EVAL_20(dmOuter__EVAL_20),
    ._EVAL_21(dmOuter__EVAL_21)
  );
  _EVAL_122 intsource (
    ._EVAL(intsource__EVAL),
    ._EVAL_0(intsource__EVAL_0)
  );
  _EVAL_119 dmi2tl (
    ._EVAL(dmi2tl__EVAL),
    ._EVAL_0(dmi2tl__EVAL_0),
    ._EVAL_1(dmi2tl__EVAL_1),
    ._EVAL_2(dmi2tl__EVAL_2),
    ._EVAL_3(dmi2tl__EVAL_3),
    ._EVAL_4(dmi2tl__EVAL_4),
    ._EVAL_5(dmi2tl__EVAL_5),
    ._EVAL_6(dmi2tl__EVAL_6),
    ._EVAL_7(dmi2tl__EVAL_7),
    ._EVAL_8(dmi2tl__EVAL_8),
    ._EVAL_9(dmi2tl__EVAL_9),
    ._EVAL_10(dmi2tl__EVAL_10),
    ._EVAL_11(dmi2tl__EVAL_11),
    ._EVAL_12(dmi2tl__EVAL_12),
    ._EVAL_13(dmi2tl__EVAL_13),
    ._EVAL_14(dmi2tl__EVAL_14),
    ._EVAL_15(dmi2tl__EVAL_15),
    ._EVAL_16(dmi2tl__EVAL_16),
    ._EVAL_17(dmi2tl__EVAL_17),
    ._EVAL_18(dmi2tl__EVAL_18)
  );
  _EVAL_127 dmiBypass (
    ._EVAL(dmiBypass__EVAL),
    ._EVAL_0(dmiBypass__EVAL_0),
    ._EVAL_1(dmiBypass__EVAL_1),
    ._EVAL_2(dmiBypass__EVAL_2),
    ._EVAL_3(dmiBypass__EVAL_3),
    ._EVAL_4(dmiBypass__EVAL_4),
    ._EVAL_5(dmiBypass__EVAL_5),
    ._EVAL_6(dmiBypass__EVAL_6),
    ._EVAL_7(dmiBypass__EVAL_7),
    ._EVAL_8(dmiBypass__EVAL_8),
    ._EVAL_9(dmiBypass__EVAL_9),
    ._EVAL_10(dmiBypass__EVAL_10),
    ._EVAL_11(dmiBypass__EVAL_11),
    ._EVAL_12(dmiBypass__EVAL_12),
    ._EVAL_13(dmiBypass__EVAL_13),
    ._EVAL_14(dmiBypass__EVAL_14),
    ._EVAL_15(dmiBypass__EVAL_15),
    ._EVAL_16(dmiBypass__EVAL_16),
    ._EVAL_17(dmiBypass__EVAL_17),
    ._EVAL_18(dmiBypass__EVAL_18),
    ._EVAL_19(dmiBypass__EVAL_19),
    ._EVAL_20(dmiBypass__EVAL_20),
    ._EVAL_21(dmiBypass__EVAL_21),
    ._EVAL_22(dmiBypass__EVAL_22),
    ._EVAL_23(dmiBypass__EVAL_23),
    ._EVAL_24(dmiBypass__EVAL_24),
    ._EVAL_25(dmiBypass__EVAL_25),
    ._EVAL_26(dmiBypass__EVAL_26),
    ._EVAL_27(dmiBypass__EVAL_27),
    ._EVAL_28(dmiBypass__EVAL_28),
    ._EVAL_29(dmiBypass__EVAL_29),
    ._EVAL_30(dmiBypass__EVAL_30),
    ._EVAL_31(dmiBypass__EVAL_31),
    ._EVAL_32(dmiBypass__EVAL_32),
    ._EVAL_33(dmiBypass__EVAL_33)
  );
  assign dmi2tl__EVAL_18 = _EVAL_29;
  assign dmOuter__EVAL_20 = dmiXbar__EVAL_7;
  assign dmiBypass__EVAL = _EVAL_8;
  assign dmiBypass__EVAL_32 = asource__EVAL_24;
  assign dmOuter__EVAL_10 = _EVAL_8;
  assign dmi2tl__EVAL_1 = dmiXbar__EVAL_14;
  assign dmOuter__EVAL_16 = dmiXbar__EVAL_27;
  assign _EVAL_20 = AsyncQueueSource__EVAL_6;
  assign dmi2tl__EVAL_10 = dmiXbar__EVAL_35;
  assign dmiXbar__EVAL_24 = dmi2tl__EVAL_14;
  assign dmiBypass__EVAL_29 = asource__EVAL_26;
  assign dmOuter__EVAL = dmiXbar__EVAL_18;
  assign _EVAL_22 = AsyncQueueSource__EVAL_10;
  assign dmi2tl__EVAL_3 = _EVAL_2;
  assign dmiXbar__EVAL_16 = dmiBypass__EVAL_20;
  assign asource__EVAL_7 = _EVAL_8;
  assign dmiXbar__EVAL_23 = dmOuter__EVAL_0;
  assign AsyncQueueSource__EVAL_3 = dmOuter__EVAL_7;
  assign dmiXbar__EVAL_29 = dmiBypass__EVAL_28;
  assign _EVAL_14 = dmOuter__EVAL_6;
  assign asource__EVAL_1 = _EVAL_13;
  assign intsource__EVAL_0 = dmOuter__EVAL_12;
  assign dmiBypass__EVAL_14 = dmiXbar__EVAL_30;
  assign _EVAL_0 = asource__EVAL_4;
  assign AsyncQueueSource__EVAL_9 = _EVAL_8;
  assign dmOuter__EVAL_5 = dmiXbar__EVAL_33;
  assign AsyncQueueSource__EVAL_1 = _EVAL_31;
  assign asource__EVAL_14 = _EVAL_19;
  assign dmOuter__EVAL_4 = AsyncQueueSource__EVAL;
  assign dmi2tl__EVAL_12 = _EVAL_24;
  assign dmiXbar__EVAL_6 = dmOuter__EVAL_11;
  assign asource__EVAL_16 = _EVAL_3;
  assign dmi2tl__EVAL_4 = _EVAL_4;
  assign dmiXbar__EVAL_28 = dmOuter__EVAL_8;
  assign dmactiveAckSync__EVAL_0 = _EVAL_8;
  assign dmiXbar__EVAL_10 = dmiBypass__EVAL_1;
  assign _EVAL_6 = AsyncQueueSource__EVAL_0;
  assign dmiXbar__EVAL_5 = dmiBypass__EVAL_13;
  assign dmiXbar__EVAL_3 = dmi2tl__EVAL_16;
  assign AsyncQueueSource__EVAL_2 = dmOuter__EVAL_18;
  assign _EVAL_15 = dmi2tl__EVAL_11;
  assign _EVAL_23 = AsyncQueueSource__EVAL_7;
  assign dmactiveAckSync__EVAL = _EVAL_27;
  assign dmiXbar__EVAL_11 = dmiBypass__EVAL_6;
  assign asource__EVAL_11 = dmiBypass__EVAL_2;
  assign asource__EVAL_25 = _EVAL_11;
  assign dmi2tl__EVAL_0 = _EVAL_1;
  assign dmiXbar__EVAL_37 = dmOuter__EVAL_19;
  assign dmiXbar__EVAL_12 = dmi2tl__EVAL_17;
  assign _EVAL_26 = intsource__EVAL;
  assign dmiBypass__EVAL_17 = dmiXbar__EVAL_4;
  assign AsyncQueueSource__EVAL_4 = dmOuter__EVAL_14;
  assign dmiBypass__EVAL_7 = asource__EVAL_13;
  assign dmiXbar__EVAL = dmi2tl__EVAL_6;
  assign dmi2tl__EVAL_15 = dmiXbar__EVAL_25;
  assign dmiXbar__EVAL_26 = dmiBypass__EVAL_21;
  assign _EVAL_16 = asource__EVAL_2;
  assign dmiBypass__EVAL_25 = _EVAL_32 | _EVAL_33;
  assign dmiXbar__EVAL_34 = dmiBypass__EVAL_4;
  assign _EVAL_32 = ~_EVAL;
  assign asource__EVAL_17 = dmiBypass__EVAL_12;
  assign dmOuter__EVAL_1 = dmiXbar__EVAL_36;
  assign _EVAL_28 = asource__EVAL_5;
  assign _EVAL_12 = dmi2tl__EVAL_2;
  assign _EVAL_21 = asource__EVAL_21;
  assign _EVAL_18 = asource__EVAL_3;
  assign AsyncQueueSource__EVAL_5 = dmOuter__EVAL_9;
  assign asource__EVAL_6 = dmiBypass__EVAL_15;
  assign dmOuter__EVAL_15 = dmiXbar__EVAL_9;
  assign _EVAL_34 = dmactiveAckSync__EVAL_1;
  assign asource__EVAL_28 = _EVAL_7;
  assign dmiBypass__EVAL_30 = dmiXbar__EVAL_2;
  assign _EVAL_30 = dmi2tl__EVAL_7;
  assign dmiXbar__EVAL_32 = dmiBypass__EVAL_33;
  assign _EVAL = dmOuter__EVAL_13;
  assign AsyncQueueSource__EVAL_8 = _EVAL_3;
  assign _EVAL_25 = dmi2tl__EVAL_5;
  assign dmiXbar__EVAL_19 = dmiBypass__EVAL_27;
  assign dmiXbar__EVAL_31 = dmi2tl__EVAL_8;
  assign dmiBypass__EVAL_24 = dmiXbar__EVAL_1;
  assign dmiXbar__EVAL_0 = dmi2tl__EVAL_13;
  assign dmactiveAckSync__EVAL_2 = _EVAL_3;
  assign asource__EVAL_20 = _EVAL_17;
  assign dmi2tl__EVAL = dmiXbar__EVAL_15;
  assign dmiBypass__EVAL_3 = asource__EVAL_10;
  assign dmiBypass__EVAL_26 = asource__EVAL_8;
  assign dmiBypass__EVAL_18 = dmiXbar__EVAL_22;
  assign dmiBypass__EVAL_9 = asource__EVAL_27;
  assign dmiXbar__EVAL_13 = _EVAL_3;
  assign _EVAL_5 = asource__EVAL_22;
  assign _EVAL_33 = ~_EVAL_34;
  assign dmiBypass__EVAL_16 = asource__EVAL;
  assign dmOuter__EVAL_17 = dmactiveAckSync__EVAL_1;
  assign dmOuter__EVAL_2 = _EVAL_9;
  assign asource__EVAL_9 = _EVAL_10;
  assign dmiBypass__EVAL_5 = asource__EVAL_23;
  assign asource__EVAL_12 = dmiBypass__EVAL_10;
  assign dmiBypass__EVAL_23 = asource__EVAL_18;
  assign dmiXbar__EVAL_21 = _EVAL_8;
  assign dmiBypass__EVAL_8 = dmiXbar__EVAL_20;
  assign dmiBypass__EVAL_19 = asource__EVAL_19;
  assign asource__EVAL_15 = dmiBypass__EVAL_0;
  assign dmiBypass__EVAL_22 = _EVAL_3;
  assign dmiXbar__EVAL_17 = dmiBypass__EVAL_11;
  assign dmOuter__EVAL_3 = _EVAL_3;
  assign dmi2tl__EVAL_9 = dmiXbar__EVAL_8;
  assign asource__EVAL_0 = dmiBypass__EVAL_31;
endmodule
