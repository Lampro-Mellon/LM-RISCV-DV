//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_75(
  input         _EVAL,
  input  [3:0]  _EVAL_0,
  output        _EVAL_1,
  input         _EVAL_2,
  output        _EVAL_3,
  output [2:0]  _EVAL_4,
  output [2:0]  _EVAL_5,
  output [2:0]  _EVAL_6,
  output [3:0]  _EVAL_7,
  output        _EVAL_8,
  input  [2:0]  _EVAL_9,
  output [31:0] _EVAL_10,
  input         _EVAL_11,
  output [3:0]  _EVAL_12,
  output        _EVAL_13,
  input  [3:0]  _EVAL_14,
  output        _EVAL_15,
  input  [2:0]  _EVAL_16,
  output        _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  output [1:0]  _EVAL_20,
  output [2:0]  _EVAL_21,
  output [3:0]  _EVAL_22,
  input  [2:0]  _EVAL_23,
  output        _EVAL_24,
  input         _EVAL_25,
  input  [2:0]  _EVAL_26,
  input         _EVAL_27,
  input  [13:0] _EVAL_28,
  input         _EVAL_29,
  input  [3:0]  _EVAL_30,
  input  [2:0]  _EVAL_31,
  output [13:0] _EVAL_32,
  output [2:0]  _EVAL_33,
  output        _EVAL_34
);
  wire [2:0] Queue__EVAL;
  wire [2:0] Queue__EVAL_0;
  wire  Queue__EVAL_1;
  wire  Queue__EVAL_2;
  wire  Queue__EVAL_3;
  wire [2:0] Queue__EVAL_4;
  wire [13:0] Queue__EVAL_5;
  wire [2:0] Queue__EVAL_6;
  wire [3:0] Queue__EVAL_7;
  wire  Queue__EVAL_8;
  wire [3:0] Queue__EVAL_9;
  wire [2:0] Queue__EVAL_10;
  wire [2:0] Queue__EVAL_11;
  wire [3:0] Queue__EVAL_12;
  wire  Queue__EVAL_13;
  wire  Queue__EVAL_14;
  wire  Queue__EVAL_15;
  wire  Queue__EVAL_16;
  wire [3:0] Queue__EVAL_17;
  wire [13:0] Queue__EVAL_18;
  wire  Queue_1__EVAL;
  wire [2:0] Queue_1__EVAL_0;
  wire  Queue_1__EVAL_1;
  wire  Queue_1__EVAL_2;
  wire  Queue_1__EVAL_3;
  wire  Queue_1__EVAL_4;
  wire  Queue_1__EVAL_5;
  wire [3:0] Queue_1__EVAL_6;
  wire  Queue_1__EVAL_7;
  wire [1:0] Queue_1__EVAL_8;
  wire [31:0] Queue_1__EVAL_9;
  wire [1:0] Queue_1__EVAL_10;
  wire [31:0] Queue_1__EVAL_11;
  wire [2:0] Queue_1__EVAL_12;
  wire [3:0] Queue_1__EVAL_13;
  wire  Queue_1__EVAL_14;
  wire  Queue_1__EVAL_15;
  wire [2:0] Queue_1__EVAL_16;
  wire  Queue_1__EVAL_17;
  wire  Queue_1__EVAL_18;
  wire  Queue_1__EVAL_19;
  wire [2:0] Queue_1__EVAL_20;
  _EVAL_74 Queue (
    ._EVAL(Queue__EVAL),
    ._EVAL_0(Queue__EVAL_0),
    ._EVAL_1(Queue__EVAL_1),
    ._EVAL_2(Queue__EVAL_2),
    ._EVAL_3(Queue__EVAL_3),
    ._EVAL_4(Queue__EVAL_4),
    ._EVAL_5(Queue__EVAL_5),
    ._EVAL_6(Queue__EVAL_6),
    ._EVAL_7(Queue__EVAL_7),
    ._EVAL_8(Queue__EVAL_8),
    ._EVAL_9(Queue__EVAL_9),
    ._EVAL_10(Queue__EVAL_10),
    ._EVAL_11(Queue__EVAL_11),
    ._EVAL_12(Queue__EVAL_12),
    ._EVAL_13(Queue__EVAL_13),
    ._EVAL_14(Queue__EVAL_14),
    ._EVAL_15(Queue__EVAL_15),
    ._EVAL_16(Queue__EVAL_16),
    ._EVAL_17(Queue__EVAL_17),
    ._EVAL_18(Queue__EVAL_18)
  );
  _EVAL_66 Queue_1 (
    ._EVAL(Queue_1__EVAL),
    ._EVAL_0(Queue_1__EVAL_0),
    ._EVAL_1(Queue_1__EVAL_1),
    ._EVAL_2(Queue_1__EVAL_2),
    ._EVAL_3(Queue_1__EVAL_3),
    ._EVAL_4(Queue_1__EVAL_4),
    ._EVAL_5(Queue_1__EVAL_5),
    ._EVAL_6(Queue_1__EVAL_6),
    ._EVAL_7(Queue_1__EVAL_7),
    ._EVAL_8(Queue_1__EVAL_8),
    ._EVAL_9(Queue_1__EVAL_9),
    ._EVAL_10(Queue_1__EVAL_10),
    ._EVAL_11(Queue_1__EVAL_11),
    ._EVAL_12(Queue_1__EVAL_12),
    ._EVAL_13(Queue_1__EVAL_13),
    ._EVAL_14(Queue_1__EVAL_14),
    ._EVAL_15(Queue_1__EVAL_15),
    ._EVAL_16(Queue_1__EVAL_16),
    ._EVAL_17(Queue_1__EVAL_17),
    ._EVAL_18(Queue_1__EVAL_18),
    ._EVAL_19(Queue_1__EVAL_19),
    ._EVAL_20(Queue_1__EVAL_20)
  );
  assign Queue__EVAL_16 = _EVAL_18;
  assign _EVAL_21 = Queue_1__EVAL_12;
  assign Queue_1__EVAL_1 = _EVAL_25;
  assign _EVAL_3 = Queue_1__EVAL_17;
  assign Queue__EVAL_6 = _EVAL_31;
  assign _EVAL_15 = Queue__EVAL_2;
  assign Queue_1__EVAL_2 = 1'h0;
  assign _EVAL_5 = Queue_1__EVAL_16;
  assign _EVAL_20 = Queue_1__EVAL_8;
  assign _EVAL_1 = Queue_1__EVAL_15;
  assign _EVAL_6 = Queue__EVAL_0;
  assign Queue_1__EVAL_13 = _EVAL_14;
  assign Queue__EVAL_10 = _EVAL_23;
  assign _EVAL_22 = Queue_1__EVAL_6;
  assign Queue__EVAL_15 = _EVAL;
  assign Queue_1__EVAL_20 = _EVAL_9;
  assign _EVAL_24 = Queue_1__EVAL_4;
  assign _EVAL_13 = Queue_1__EVAL;
  assign Queue_1__EVAL_7 = 1'h1;
  assign _EVAL_8 = Queue__EVAL_8;
  assign _EVAL_17 = Queue_1__EVAL_14;
  assign _EVAL_7 = Queue__EVAL_9;
  assign _EVAL_33 = Queue__EVAL_4;
  assign Queue__EVAL_12 = _EVAL_30;
  assign _EVAL_12 = Queue__EVAL_17;
  assign _EVAL_34 = Queue__EVAL_1;
  assign Queue_1__EVAL_5 = _EVAL_11;
  assign Queue__EVAL_3 = _EVAL_19;
  assign Queue__EVAL_14 = _EVAL_29;
  assign Queue__EVAL_18 = _EVAL_28;
  assign Queue_1__EVAL_0 = _EVAL_16;
  assign Queue_1__EVAL_18 = _EVAL_19;
  assign Queue_1__EVAL_9 = 32'h0;
  assign Queue__EVAL_7 = _EVAL_0;
  assign Queue__EVAL_13 = _EVAL_27;
  assign Queue_1__EVAL_10 = 2'h0;
  assign Queue_1__EVAL_19 = _EVAL_2;
  assign Queue__EVAL = _EVAL_26;
  assign _EVAL_10 = Queue_1__EVAL_11;
  assign _EVAL_4 = Queue__EVAL_11;
  assign Queue_1__EVAL_3 = _EVAL_27;
  assign _EVAL_32 = Queue__EVAL_5;
endmodule
