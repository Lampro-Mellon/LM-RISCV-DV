//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_151(
  output        _EVAL,
  input  [31:0] _EVAL_0,
  output        _EVAL_1,
  output [4:0]  _EVAL_2,
  output [4:0]  _EVAL_3,
  output        _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  output [4:0]  _EVAL_7,
  output        _EVAL_8,
  output        _EVAL_9,
  input         _EVAL_10,
  output [31:0] _EVAL_11,
  input         _EVAL_12,
  input  [31:0] _EVAL_13,
  input         _EVAL_14,
  output [31:0] _EVAL_15,
  input         _EVAL_16,
  output [4:0]  _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  output        _EVAL_20,
  input  [31:0] _EVAL_21,
  output        _EVAL_22,
  input         _EVAL_23
);
  reg [15:0] _EVAL_25;
  reg [31:0] _RAND_0;
  wire [2:0] _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  reg [15:0] _EVAL_38;
  reg [31:0] _RAND_1;
  wire [2:0] _EVAL_40;
  wire  _EVAL_42;
  reg  _EVAL_43;
  reg [31:0] _RAND_2;
  wire  _EVAL_44;
  wire [2:0] _EVAL_46;
  wire  _EVAL_47;
  wire [3:0] _EVAL_48;
  wire [2:0] _EVAL_49;
  wire  _EVAL_52;
  wire [15:0] _EVAL_54;
  reg  _EVAL_55;
  reg [31:0] _RAND_3;
  wire  _EVAL_58;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_65;
  reg [15:0] _EVAL_66;
  reg [31:0] _RAND_4;
  wire  _EVAL_67;
  wire  _EVAL_72;
  wire  _EVAL_74;
  reg [2:0] _EVAL_75;
  reg [31:0] _RAND_5;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire [2:0] _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_85;
  wire  _EVAL_86;
  reg [2:0] _EVAL_87;
  reg [31:0] _RAND_6;
  wire [1:0] _EVAL_89;
  wire  _EVAL_90;
  wire [3:0] _EVAL_91;
  reg  _EVAL_92;
  reg [31:0] _RAND_7;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire [2:0] _EVAL_98;
  wire [3:0] _EVAL_100;
  reg [15:0] _EVAL_101;
  reg [31:0] _RAND_8;
  wire  _EVAL_103;
  wire  _EVAL_105;
  wire [2:0] _EVAL_106;
  wire  _EVAL_107;
  wire [2:0] _EVAL_108;
  wire [3:0] _EVAL_114;
  reg [15:0] _EVAL_115;
  reg [31:0] _RAND_9;
  wire  _EVAL_116;
  reg  _EVAL_118;
  reg [31:0] _RAND_10;
  wire  _EVAL_119;
  wire  _EVAL_120;
  reg  _EVAL_122;
  reg [31:0] _RAND_11;
  wire [2:0] _EVAL_123;
  wire  _EVAL_124;
  reg [31:0] _EVAL_128;
  reg [31:0] _RAND_12;
  wire  _EVAL_132;
  wire [2:0] _EVAL_133;
  wire  _EVAL_138;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_144;
  wire [2:0] _EVAL_145;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire [2:0] _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire [15:0] _EVAL_155;
  wire [3:0] _EVAL_156;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire [2:0] _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_175;
  wire [3:0] _EVAL_181;
  wire  _EVAL_184;
  reg  _EVAL_185;
  reg [31:0] _RAND_13;
  wire  _EVAL_186;
  reg  _EVAL_188;
  reg [31:0] _RAND_14;
  reg [2:0] _EVAL_190;
  reg [31:0] _RAND_15;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire [4:0] expander__EVAL;
  wire [4:0] expander__EVAL_0;
  wire  expander__EVAL_1;
  wire [31:0] expander__EVAL_2;
  wire [4:0] expander__EVAL_3;
  wire [31:0] expander__EVAL_4;
  reg  _EVAL_196;
  reg [31:0] _RAND_16;
  wire  _EVAL_199;
  reg  _EVAL_201;
  reg [31:0] _RAND_17;
  wire [2:0] _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_206;
  wire [15:0] _EVAL_207;
  reg [15:0] _EVAL_209;
  reg [31:0] _RAND_18;
  reg  _EVAL_210;
  reg [31:0] _RAND_19;
  reg [15:0] _EVAL_211;
  reg [31:0] _RAND_20;
  reg  _EVAL_212;
  reg [31:0] _RAND_21;
  reg  _EVAL_213;
  reg [31:0] _RAND_22;
  wire [3:0] _EVAL_215;
  wire  _EVAL_216;
  wire [2:0] _EVAL_217;
  reg  _EVAL_218;
  reg [31:0] _RAND_23;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire [3:0] _EVAL_221;
  wire [15:0] _EVAL_225;
  wire  _EVAL_230;
  wire [2:0] _EVAL_233;
  reg  _EVAL_238;
  reg [31:0] _RAND_24;
  wire  _EVAL_240;
  wire [2:0] _EVAL_242;
  wire [15:0] _EVAL_244;
  wire [15:0] _EVAL_245;
  wire [1:0] _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  _EVAL_150 expander (
    ._EVAL(expander__EVAL),
    ._EVAL_0(expander__EVAL_0),
    ._EVAL_1(expander__EVAL_1),
    ._EVAL_2(expander__EVAL_2),
    ._EVAL_3(expander__EVAL_3),
    ._EVAL_4(expander__EVAL_4)
  );
  assign _EVAL_216 = ~_EVAL_55;
  assign _EVAL_9 = _EVAL_122 | _EVAL_201;
  assign _EVAL_144 = _EVAL_108 == 3'h1;
  assign _EVAL_147 = _EVAL_87 > 3'h3;
  assign _EVAL_203 = _EVAL_220 ? 1'h0 : _EVAL_118;
  assign _EVAL_62 = _EVAL_233 == 3'h1;
  assign _EVAL_17 = {_EVAL_181, 1'h0};
  assign _EVAL_58 = _EVAL_18 != _EVAL_55;
  assign _EVAL_48 = _EVAL_87 - _EVAL_80;
  assign _EVAL_78 = _EVAL_33 & _EVAL_184;
  assign _EVAL_46 = _EVAL_201 ? _EVAL_26 : 3'h0;
  assign _EVAL_162 = _EVAL_55 ? _EVAL_201 : _EVAL_122;
  assign _EVAL_202 = {{2'd0}, _EVAL_138};
  assign _EVAL_168 = _EVAL_103 & _EVAL_163;
  assign _EVAL_54 = _EVAL_220 ? _EVAL_225 : _EVAL_244;
  assign _EVAL_89 = _EVAL_52 ? _EVAL_246 : 2'h0;
  assign _EVAL_199 = _EVAL_87 >= 3'h1;
  assign _EVAL_233 = _EVAL_48[2:0];
  assign _EVAL_225 = _EVAL_128[31:16];
  assign _EVAL_206 = _EVAL_216 | _EVAL_166;
  assign _EVAL_163 = _EVAL_246 >= 2'h1;
  assign _EVAL_107 = _EVAL_87 > 3'h6;
  assign _EVAL_40 = _EVAL_100[2:0];
  assign _EVAL_221 = 3'h7 - _EVAL_151;
  assign _EVAL_217 = _EVAL_221[2:0];
  assign _EVAL_242 = _EVAL_248 ? _EVAL_49 : 3'h0;
  assign _EVAL_100 = 3'h2 - _EVAL_190;
  assign _EVAL_1 = _EVAL_81 & _EVAL_210;
  assign _EVAL_204 = _EVAL_175 | _EVAL_203;
  assign _EVAL_33 = _EVAL_87 > 3'h5;
  assign _EVAL_32 = _EVAL_124 ? _EVAL_206 : _EVAL_166;
  assign _EVAL_181 = _EVAL_242 + _EVAL_87;
  assign _EVAL_133 = _EVAL_215[2:0];
  assign _EVAL_207 = _EVAL_220 ? _EVAL_155 : _EVAL_245;
  assign _EVAL_7 = expander__EVAL;
  assign _EVAL_186 = _EVAL_147 & _EVAL_184;
  assign _EVAL_22 = _EVAL_42 & _EVAL_116;
  assign _EVAL_11 = expander__EVAL_4;
  assign _EVAL_165 = _EVAL_140 & _EVAL_162;
  assign _EVAL_140 = _EVAL_14 & _EVAL_58;
  assign _EVAL_27 = _EVAL_233 == 3'h0;
  assign _EVAL_120 = ~_EVAL_94;
  assign _EVAL_142 = _EVAL_216 | _EVAL_32;
  assign _EVAL_167 = {{1'd0}, _EVAL_246};
  assign _EVAL_219 = _EVAL_87 > 3'h2;
  assign _EVAL_116 = ~_EVAL_162;
  assign _EVAL_108 = _EVAL_47 ? _EVAL_75 : _EVAL_190;
  assign _EVAL_152 = _EVAL_67 | _EVAL_220;
  assign _EVAL_240 = _EVAL_22 & _EVAL_6;
  assign _EVAL_141 = _EVAL_55 | _EVAL_30;
  assign _EVAL_94 = _EVAL_169 & _EVAL_42;
  assign _EVAL_215 = 3'h2 - _EVAL_108;
  assign _EVAL_106 = _EVAL_122 ? _EVAL_40 : 3'h0;
  assign _EVAL_65 = ~_EVAL_248;
  assign _EVAL_138 = _EVAL_21[1];
  assign _EVAL_15 = expander__EVAL_2;
  assign _EVAL_80 = {{1'd0}, _EVAL_89};
  assign _EVAL_86 = _EVAL_18 ? 1'h0 : _EVAL_201;
  assign _EVAL_30 = _EVAL_14 ? _EVAL_86 : _EVAL_201;
  assign _EVAL_103 = _EVAL_87 > 3'h4;
  assign _EVAL_67 = _EVAL_14 & _EVAL_120;
  assign _EVAL_3 = expander__EVAL_3;
  assign _EVAL_4 = _EVAL_238;
  assign _EVAL_114 = 3'h2 - _EVAL_75;
  assign _EVAL_8 = expander__EVAL_1;
  assign _EVAL_98 = _EVAL_91[2:0];
  assign _EVAL_148 = _EVAL_103 & _EVAL_184;
  assign _EVAL_132 = _EVAL_220 ? _EVAL_212 : _EVAL_5;
  assign _EVAL_124 = _EVAL_16 & _EVAL_1;
  assign expander__EVAL_4 = {_EVAL_38,_EVAL_66};
  assign _EVAL = _EVAL_153 | _EVAL_230;
  assign _EVAL_47 = _EVAL_220 ? _EVAL_185 : _EVAL_18;
  assign _EVAL_151 = 3'h2 << _EVAL_248;
  assign _EVAL_184 = _EVAL_246 >= 2'h2;
  assign _EVAL_246 = 2'h2 >> expander__EVAL_1;
  assign _EVAL_91 = _EVAL_233 + _EVAL_145;
  assign _EVAL_123 = {{2'd0}, _EVAL_90};
  assign _EVAL_72 = _EVAL_124 ? _EVAL_141 : _EVAL_30;
  assign _EVAL_79 = _EVAL_233 == 3'h4;
  assign _EVAL_247 = _EVAL_33 & _EVAL_163;
  assign _EVAL_61 = _EVAL_42 & _EVAL_116;
  assign _EVAL_194 = _EVAL_233 == 3'h3;
  assign _EVAL_164 = _EVAL_55 | _EVAL_72;
  assign _EVAL_26 = _EVAL_114[2:0];
  assign _EVAL_156 = _EVAL_106 + _EVAL_46;
  assign _EVAL_31 = _EVAL_219 & _EVAL_163;
  assign _EVAL_248 = _EVAL_122 | _EVAL_201;
  assign _EVAL_145 = _EVAL_152 ? _EVAL_133 : 3'h0;
  assign _EVAL_153 = _EVAL_87 >= _EVAL_167;
  assign _EVAL_105 = _EVAL_233 == 3'h5;
  assign _EVAL_245 = _EVAL_0[15:0];
  assign _EVAL_155 = _EVAL_128[15:0];
  assign _EVAL_52 = _EVAL_10 & _EVAL;
  assign _EVAL_93 = _EVAL_233 == 3'h2;
  assign _EVAL_220 = _EVAL_118 & _EVAL_65;
  assign _EVAL_230 = _EVAL_199 & _EVAL_238;
  assign _EVAL_119 = _EVAL_107 & _EVAL_163;
  assign _EVAL_193 = ~_EVAL_18 ? 1'h0 : _EVAL_122;
  assign _EVAL_49 = _EVAL_156[2:0];
  assign _EVAL_175 = _EVAL_165 & _EVAL_42;
  assign _EVAL_81 = _EVAL_61 & _EVAL_44;
  assign _EVAL_85 = _EVAL_107 & _EVAL_184;
  assign _EVAL_74 = _EVAL_147 & _EVAL_163;
  assign _EVAL_166 = _EVAL_14 ? _EVAL_193 : _EVAL_122;
  assign _EVAL_2 = expander__EVAL_0;
  assign _EVAL_44 = _EVAL_87 <= _EVAL_217;
  assign _EVAL_42 = ~_EVAL_118;
  assign _EVAL_20 = _EVAL_55;
  assign _EVAL_169 = _EVAL_58 & _EVAL_162;
  assign _EVAL_90 = _EVAL_13[1];
  assign _EVAL_244 = _EVAL_0[31:16];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_25 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_38 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_43 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_55 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_66 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_75 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_87 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_92 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_101 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_115 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_118 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_122 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_128 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_185 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_188 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_190 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_196 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_201 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_209 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_210 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_211 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_212 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_213 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_218 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_238 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_12) begin
    if (_EVAL_152) begin
      if (_EVAL_62) begin
        if (_EVAL_220) begin
          _EVAL_25 <= _EVAL_225;
        end else begin
          _EVAL_25 <= _EVAL_244;
        end
      end else if (_EVAL_93) begin
        if (_EVAL_220) begin
          _EVAL_25 <= _EVAL_155;
        end else begin
          _EVAL_25 <= _EVAL_245;
        end
      end else if (_EVAL_52) begin
        if (_EVAL_148) begin
          _EVAL_25 <= _EVAL_101;
        end else if (_EVAL_74) begin
          _EVAL_25 <= _EVAL_115;
        end
      end
    end else if (_EVAL_52) begin
      if (_EVAL_148) begin
        _EVAL_25 <= _EVAL_101;
      end else if (_EVAL_74) begin
        _EVAL_25 <= _EVAL_115;
      end
    end
    if (_EVAL_152) begin
      if (_EVAL_27) begin
        if (_EVAL_220) begin
          _EVAL_38 <= _EVAL_225;
        end else begin
          _EVAL_38 <= _EVAL_244;
        end
      end else if (_EVAL_62) begin
        if (_EVAL_220) begin
          _EVAL_38 <= _EVAL_155;
        end else begin
          _EVAL_38 <= _EVAL_245;
        end
      end else if (_EVAL_52) begin
        if (_EVAL_186) begin
          _EVAL_38 <= _EVAL_115;
        end else if (_EVAL_31) begin
          _EVAL_38 <= _EVAL_25;
        end
      end
    end else if (_EVAL_52) begin
      if (_EVAL_186) begin
        _EVAL_38 <= _EVAL_115;
      end else if (_EVAL_31) begin
        _EVAL_38 <= _EVAL_25;
      end
    end
    if (_EVAL_152) begin
      if (_EVAL_27) begin
        if (_EVAL_220) begin
          _EVAL_43 <= _EVAL_212;
        end else begin
          _EVAL_43 <= _EVAL_5;
        end
      end else if (_EVAL_62) begin
        if (_EVAL_220) begin
          _EVAL_43 <= _EVAL_212;
        end else begin
          _EVAL_43 <= _EVAL_5;
        end
      end else if (_EVAL_52) begin
        if (_EVAL_186) begin
          _EVAL_43 <= _EVAL_92;
        end else if (_EVAL_31) begin
          _EVAL_43 <= _EVAL_196;
        end
      end
    end else if (_EVAL_52) begin
      if (_EVAL_186) begin
        _EVAL_43 <= _EVAL_92;
      end else if (_EVAL_31) begin
        _EVAL_43 <= _EVAL_196;
      end
    end
    if (_EVAL_240) begin
      _EVAL_55 <= _EVAL_216;
    end else if (_EVAL_124) begin
      _EVAL_55 <= _EVAL_216;
    end
    if (_EVAL_152) begin
      if (_EVAL_144) begin
        if (_EVAL_220) begin
          _EVAL_66 <= _EVAL_225;
        end else begin
          _EVAL_66 <= _EVAL_244;
        end
      end else if (_EVAL_27) begin
        if (_EVAL_220) begin
          _EVAL_66 <= _EVAL_155;
        end else begin
          _EVAL_66 <= _EVAL_245;
        end
      end else if (_EVAL_52) begin
        if (_EVAL_184) begin
          _EVAL_66 <= _EVAL_25;
        end else if (_EVAL_163) begin
          _EVAL_66 <= _EVAL_38;
        end
      end
    end else if (_EVAL_52) begin
      if (_EVAL_184) begin
        _EVAL_66 <= _EVAL_25;
      end else if (_EVAL_163) begin
        _EVAL_66 <= _EVAL_38;
      end
    end
    if (_EVAL_240) begin
      if (_EVAL_55) begin
        _EVAL_75 <= _EVAL_202;
      end else if (_EVAL_19) begin
        _EVAL_75 <= 3'h2;
      end else if (_EVAL_124) begin
        if (_EVAL_55) begin
          _EVAL_75 <= _EVAL_123;
        end
      end
    end else if (_EVAL_19) begin
      _EVAL_75 <= 3'h2;
    end else if (_EVAL_124) begin
      if (_EVAL_55) begin
        _EVAL_75 <= _EVAL_123;
      end
    end
    if (_EVAL_23) begin
      _EVAL_87 <= 3'h0;
    end else if (_EVAL_19) begin
      _EVAL_87 <= 3'h0;
    end else begin
      _EVAL_87 <= _EVAL_98;
    end
    if (_EVAL_152) begin
      if (_EVAL_93) begin
        if (_EVAL_220) begin
          _EVAL_92 <= _EVAL_212;
        end else begin
          _EVAL_92 <= _EVAL_5;
        end
      end else if (_EVAL_194) begin
        if (_EVAL_220) begin
          _EVAL_92 <= _EVAL_212;
        end else begin
          _EVAL_92 <= _EVAL_5;
        end
      end else if (_EVAL_52) begin
        if (_EVAL_78) begin
          _EVAL_92 <= _EVAL_213;
        end else if (_EVAL_168) begin
          _EVAL_92 <= _EVAL_188;
        end
      end
    end else if (_EVAL_52) begin
      if (_EVAL_78) begin
        _EVAL_92 <= _EVAL_213;
      end else if (_EVAL_168) begin
        _EVAL_92 <= _EVAL_188;
      end
    end
    if (_EVAL_152) begin
      if (_EVAL_194) begin
        if (_EVAL_220) begin
          _EVAL_101 <= _EVAL_225;
        end else begin
          _EVAL_101 <= _EVAL_244;
        end
      end else if (_EVAL_79) begin
        if (_EVAL_220) begin
          _EVAL_101 <= _EVAL_155;
        end else begin
          _EVAL_101 <= _EVAL_245;
        end
      end else if (_EVAL_52) begin
        if (_EVAL_85) begin
          _EVAL_101 <= _EVAL_211;
        end else if (_EVAL_247) begin
          _EVAL_101 <= _EVAL_209;
        end
      end
    end else if (_EVAL_52) begin
      if (_EVAL_85) begin
        _EVAL_101 <= _EVAL_211;
      end else if (_EVAL_247) begin
        _EVAL_101 <= _EVAL_209;
      end
    end
    if (_EVAL_152) begin
      if (_EVAL_93) begin
        _EVAL_115 <= _EVAL_54;
      end else if (_EVAL_194) begin
        _EVAL_115 <= _EVAL_207;
      end else if (_EVAL_52) begin
        if (_EVAL_78) begin
          _EVAL_115 <= _EVAL_209;
        end else if (_EVAL_168) begin
          _EVAL_115 <= _EVAL_101;
        end
      end
    end else if (_EVAL_52) begin
      if (_EVAL_78) begin
        _EVAL_115 <= _EVAL_209;
      end else if (_EVAL_168) begin
        _EVAL_115 <= _EVAL_101;
      end
    end
    if (_EVAL_23) begin
      _EVAL_118 <= 1'h0;
    end else begin
      _EVAL_118 <= _EVAL_204;
    end
    if (_EVAL_23) begin
      _EVAL_122 <= 1'h0;
    end else if (_EVAL_240) begin
      _EVAL_122 <= _EVAL_142;
    end else if (_EVAL_124) begin
      _EVAL_122 <= _EVAL_206;
    end else if (_EVAL_14) begin
      if (~_EVAL_18) begin
        _EVAL_122 <= 1'h0;
      end
    end
    if (_EVAL_175) begin
      _EVAL_128 <= _EVAL_0;
    end
    if (_EVAL_175) begin
      _EVAL_185 <= _EVAL_18;
    end
    if (_EVAL_152) begin
      if (_EVAL_194) begin
        _EVAL_188 <= _EVAL_132;
      end else if (_EVAL_79) begin
        _EVAL_188 <= _EVAL_132;
      end else if (_EVAL_52) begin
        if (_EVAL_85) begin
          _EVAL_188 <= _EVAL_218;
        end else if (_EVAL_247) begin
          _EVAL_188 <= _EVAL_213;
        end
      end
    end else if (_EVAL_52) begin
      if (_EVAL_85) begin
        _EVAL_188 <= _EVAL_218;
      end else if (_EVAL_247) begin
        _EVAL_188 <= _EVAL_213;
      end
    end
    if (_EVAL_240) begin
      if (~_EVAL_55) begin
        _EVAL_190 <= _EVAL_202;
      end else if (_EVAL_19) begin
        _EVAL_190 <= 3'h2;
      end else if (_EVAL_124) begin
        if (~_EVAL_55) begin
          _EVAL_190 <= _EVAL_123;
        end
      end
    end else if (_EVAL_19) begin
      _EVAL_190 <= 3'h2;
    end else if (_EVAL_124) begin
      if (~_EVAL_55) begin
        _EVAL_190 <= _EVAL_123;
      end
    end
    if (_EVAL_152) begin
      if (_EVAL_62) begin
        _EVAL_196 <= _EVAL_132;
      end else if (_EVAL_93) begin
        _EVAL_196 <= _EVAL_132;
      end else if (_EVAL_52) begin
        if (_EVAL_148) begin
          _EVAL_196 <= _EVAL_188;
        end else if (_EVAL_74) begin
          _EVAL_196 <= _EVAL_92;
        end
      end
    end else if (_EVAL_52) begin
      if (_EVAL_148) begin
        _EVAL_196 <= _EVAL_188;
      end else if (_EVAL_74) begin
        _EVAL_196 <= _EVAL_92;
      end
    end
    if (_EVAL_23) begin
      _EVAL_201 <= 1'h0;
    end else if (_EVAL_240) begin
      _EVAL_201 <= _EVAL_164;
    end else if (_EVAL_124) begin
      _EVAL_201 <= _EVAL_141;
    end else if (_EVAL_14) begin
      if (_EVAL_18) begin
        _EVAL_201 <= 1'h0;
      end
    end
    if (_EVAL_152) begin
      if (_EVAL_79) begin
        _EVAL_209 <= _EVAL_54;
      end else if (_EVAL_105) begin
        _EVAL_209 <= _EVAL_207;
      end else if (_EVAL_52) begin
        if (_EVAL_119) begin
          _EVAL_209 <= _EVAL_211;
        end
      end
    end else if (_EVAL_52) begin
      if (_EVAL_119) begin
        _EVAL_209 <= _EVAL_211;
      end
    end
    if (_EVAL_23) begin
      _EVAL_210 <= 1'h0;
    end else begin
      _EVAL_210 <= 1'h1;
    end
    if (_EVAL_152) begin
      if (_EVAL_105) begin
        _EVAL_211 <= _EVAL_54;
      end
    end
    if (_EVAL_175) begin
      _EVAL_212 <= _EVAL_5;
    end
    if (_EVAL_152) begin
      if (_EVAL_79) begin
        _EVAL_213 <= _EVAL_132;
      end else if (_EVAL_105) begin
        _EVAL_213 <= _EVAL_132;
      end else if (_EVAL_52) begin
        if (_EVAL_119) begin
          _EVAL_213 <= _EVAL_218;
        end
      end
    end else if (_EVAL_52) begin
      if (_EVAL_119) begin
        _EVAL_213 <= _EVAL_218;
      end
    end
    if (_EVAL_152) begin
      if (_EVAL_105) begin
        _EVAL_218 <= _EVAL_132;
      end
    end
    if (_EVAL_152) begin
      if (_EVAL_144) begin
        _EVAL_238 <= _EVAL_132;
      end else if (_EVAL_27) begin
        _EVAL_238 <= _EVAL_132;
      end else if (_EVAL_52) begin
        if (_EVAL_184) begin
          _EVAL_238 <= _EVAL_196;
        end else if (_EVAL_163) begin
          _EVAL_238 <= _EVAL_43;
        end
      end
    end else if (_EVAL_52) begin
      if (_EVAL_184) begin
        _EVAL_238 <= _EVAL_196;
      end else if (_EVAL_163) begin
        _EVAL_238 <= _EVAL_43;
      end
    end
  end
endmodule
