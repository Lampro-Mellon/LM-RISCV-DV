//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_63(
  output [2:0]  _EVAL,
  output        _EVAL_0,
  input  [31:0] _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [1:0]  _EVAL_3,
  output [25:0] _EVAL_4,
  input         _EVAL_5,
  output [31:0] _EVAL_6,
  input         _EVAL_7,
  input  [2:0]  _EVAL_8,
  output [3:0]  _EVAL_9,
  output        _EVAL_10,
  input  [1:0]  _EVAL_11,
  input  [3:0]  _EVAL_12,
  output        _EVAL_13,
  input  [2:0]  _EVAL_14,
  output [13:0] _EVAL_15,
  output [2:0]  _EVAL_16,
  input         _EVAL_17,
  output        _EVAL_18,
  input  [2:0]  _EVAL_19,
  input         _EVAL_20,
  input  [2:0]  _EVAL_21,
  input         _EVAL_22,
  output [31:0] _EVAL_23,
  output        _EVAL_24,
  output [2:0]  _EVAL_25,
  output [31:0] _EVAL_26,
  output        _EVAL_27,
  input  [2:0]  _EVAL_28,
  output        _EVAL_29,
  input         _EVAL_30,
  output        _EVAL_31,
  output [1:0]  _EVAL_32,
  output        _EVAL_33,
  output [1:0]  _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36,
  input  [3:0]  _EVAL_37,
  output [3:0]  _EVAL_38,
  input  [2:0]  _EVAL_39,
  input         _EVAL_40,
  output [29:0] _EVAL_41,
  output [3:0]  _EVAL_42,
  output [14:0] _EVAL_43,
  output [2:0]  _EVAL_44,
  input  [2:0]  _EVAL_45,
  input  [1:0]  _EVAL_46,
  output [2:0]  _EVAL_47,
  output        _EVAL_48,
  output [31:0] _EVAL_49,
  output [1:0]  _EVAL_50,
  output        _EVAL_51,
  input  [1:0]  _EVAL_52,
  input         _EVAL_53,
  output [3:0]  _EVAL_54,
  input  [31:0] _EVAL_55,
  output [2:0]  _EVAL_56,
  input         _EVAL_57,
  input         _EVAL_58,
  output [3:0]  _EVAL_59,
  input  [29:0] _EVAL_60,
  input         _EVAL_61,
  input  [31:0] _EVAL_62,
  input         _EVAL_63,
  output        _EVAL_64,
  output        _EVAL_65,
  output        _EVAL_66,
  output [11:0] _EVAL_67,
  output [2:0]  _EVAL_68,
  output        _EVAL_69,
  input  [2:0]  _EVAL_70,
  input         _EVAL_71,
  output        _EVAL_72,
  input  [2:0]  _EVAL_73,
  output        _EVAL_74,
  output [2:0]  _EVAL_75,
  output [2:0]  _EVAL_76,
  input  [1:0]  _EVAL_77,
  output [2:0]  _EVAL_78,
  input         _EVAL_79,
  input         _EVAL_80,
  output        _EVAL_81,
  output        _EVAL_82,
  output [3:0]  _EVAL_83,
  output        _EVAL_84,
  output [2:0]  _EVAL_85,
  input         _EVAL_86,
  input         _EVAL_87,
  output [1:0]  _EVAL_88,
  output [3:0]  _EVAL_89,
  input  [3:0]  _EVAL_90,
  input         _EVAL_91,
  output [2:0]  _EVAL_92,
  output [2:0]  _EVAL_93,
  output [1:0]  _EVAL_94,
  input  [31:0] _EVAL_95,
  input         _EVAL_96,
  output [31:0] _EVAL_97,
  input  [2:0]  _EVAL_98,
  input  [1:0]  _EVAL_99,
  input  [2:0]  _EVAL_100,
  input         _EVAL_101,
  output        _EVAL_102,
  output [2:0]  _EVAL_103,
  input  [31:0] _EVAL_104,
  output        _EVAL_105,
  input         _EVAL_106,
  input         _EVAL_107,
  input         _EVAL_108,
  output [2:0]  _EVAL_109,
  input  [2:0]  _EVAL_110,
  output        _EVAL_111,
  output [2:0]  _EVAL_112,
  output [2:0]  _EVAL_113,
  input  [31:0] _EVAL_114,
  output        _EVAL_115
);
  wire  _EVAL_116;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire [46:0] _EVAL_120;
  wire [8:0] _EVAL_121;
  wire [30:0] _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire [4:0] _EVAL_125;
  wire  _EVAL_127;
  wire [4:0] _EVAL_128;
  wire [4:0] _EVAL_129;
  wire [3:0] _EVAL_130;
  wire [5:0] _EVAL_131;
  wire [46:0] _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire [30:0] _EVAL_138;
  wire  _EVAL_140;
  wire [6:0] _EVAL_141;
  wire [7:0] _EVAL_142;
  wire [4:0] _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire [46:0] _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire [6:0] _EVAL_153;
  wire [9:0] _EVAL_154;
  wire  _EVAL_155;
  wire [46:0] _EVAL_156;
  wire [5:0] _EVAL_157;
  wire [4:0] _EVAL_158;
  wire [9:0] _EVAL_159;
  wire  _EVAL_161;
  wire [29:0] _EVAL_162;
  wire [7:0] _EVAL_163;
  reg  _EVAL_164;
  reg [31:0] _RAND_0;
  wire [46:0] _EVAL_165;
  wire  _EVAL_166;
  wire [5:0] _EVAL_167;
  wire  _EVAL_168;
  wire [30:0] _EVAL_169;
  reg [5:0] _EVAL_171;
  reg [31:0] _RAND_1;
  wire  _EVAL_174;
  wire [4:0] _EVAL_175;
  wire [30:0] _EVAL_176;
  wire [22:0] _EVAL_177;
  wire [9:0] _EVAL_178;
  wire [4:0] _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire [9:0] _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire [29:0] _EVAL_187;
  wire [30:0] _EVAL_189;
  wire [4:0] _EVAL_190;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire [4:0] _EVAL_194;
  wire [46:0] _EVAL_195;
  wire [30:0] _EVAL_196;
  wire [9:0] _EVAL_197;
  wire [4:0] _EVAL_198;
  wire  _EVAL_200;
  wire [8:0] _EVAL_201;
  wire  _EVAL_202;
  wire [4:0] _EVAL_203;
  wire [8:0] _EVAL_204;
  wire [9:0] _EVAL_205;
  wire [46:0] _EVAL_206;
  wire [30:0] _EVAL_207;
  wire  _EVAL_208;
  wire [9:0] _EVAL_209;
  wire [5:0] _EVAL_210;
  wire [30:0] _EVAL_211;
  reg  _EVAL_212;
  reg [31:0] _RAND_2;
  wire [3:0] _EVAL_213;
  wire  _EVAL_215;
  wire [4:0] _EVAL_217;
  wire [30:0] _EVAL_218;
  wire  _EVAL_222;
  wire [46:0] _EVAL_223;
  wire [30:0] _EVAL_224;
  wire [46:0] _EVAL_225;
  wire  _EVAL_226;
  wire [3:0] _EVAL_227;
  wire [4:0] _EVAL_228;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire [46:0] _EVAL_235;
  wire  _EVAL_237;
  wire [30:0] _EVAL_238;
  wire  _EVAL_240;
  reg  _EVAL_241;
  reg [31:0] _RAND_3;
  wire  _EVAL_242;
  wire [3:0] _EVAL_243;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire [9:0] _EVAL_247;
  reg  _EVAL_248;
  reg [31:0] _RAND_4;
  wire  _EVAL_250;
  wire  _EVAL_251;
  reg  _EVAL_252;
  reg [31:0] _RAND_5;
  reg [4:0] _EVAL_253;
  reg [31:0] _RAND_6;
  wire [46:0] _EVAL_254;
  wire [30:0] _EVAL_255;
  wire [5:0] _EVAL_256;
  wire [46:0] _EVAL_257;
  wire [30:0] _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire [7:0] _EVAL_262;
  wire [4:0] _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire [29:0] _EVAL_266;
  wire [9:0] _EVAL_267;
  wire [29:0] _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire [30:0] _EVAL_271;
  wire [46:0] _EVAL_272;
  wire [46:0] _EVAL_274;
  wire  _EVAL_275;
  wire [30:0] _EVAL_276;
  wire [9:0] _EVAL_279;
  assign _EVAL_254 = _EVAL_136 ? _EVAL_272 : 47'h0;
  assign _EVAL_242 = _EVAL_234 & _EVAL_96;
  assign _EVAL_81 = _EVAL_235[0];
  assign _EVAL_68 = _EVAL_39;
  assign _EVAL_161 = _EVAL_118 & _EVAL_106;
  assign _EVAL_154 = {_EVAL_198,_EVAL_80,_EVAL_106,_EVAL_71,_EVAL_96,_EVAL_107};
  assign _EVAL_127 = $signed(_EVAL_169) == 31'sh0;
  assign _EVAL_226 = _EVAL_171 == 6'h0;
  assign _EVAL_74 = _EVAL_235[33];
  assign _EVAL_78 = _EVAL_110;
  assign _EVAL_44 = _EVAL_235[46:44];
  assign _EVAL_211 = $signed(_EVAL_122) & 31'sh22000000;
  assign _EVAL_15 = _EVAL_60[13:0];
  assign _EVAL_26 = _EVAL_95;
  assign _EVAL_25 = _EVAL_110;
  assign _EVAL_201 = {_EVAL_175, 4'h0};
  assign _EVAL_166 = _EVAL_123 | _EVAL_182;
  assign _EVAL_42 = _EVAL_12;
  assign _EVAL_82 = _EVAL_36;
  assign _EVAL_4 = _EVAL_60[25:0];
  assign _EVAL_245 = _EVAL_140 & _EVAL_80;
  assign _EVAL_228 = _EVAL_201[4:0];
  assign _EVAL_128 = _EVAL_175 | _EVAL_228;
  assign _EVAL_237 = _EVAL_260 & _EVAL_107;
  assign _EVAL_112 = _EVAL_235[37:35];
  assign _EVAL_72 = _EVAL_22;
  assign _EVAL_247 = {{1'd0}, _EVAL_121};
  assign _EVAL_205 = _EVAL_183 | _EVAL_197;
  assign _EVAL_120 = _EVAL_134 ? _EVAL_223 : 47'h0;
  assign _EVAL_102 = _EVAL_40 & _EVAL_144;
  assign _EVAL_125 = _EVAL_256[4:0];
  assign _EVAL_6 = _EVAL_235[32:1];
  assign _EVAL_190 = _EVAL_194 & _EVAL_129;
  assign _EVAL_129 = _EVAL_209[4:0];
  assign _EVAL_133 = _EVAL_226 ? _EVAL_251 : _EVAL_164;
  assign _EVAL_94 = _EVAL_90[1:0];
  assign _EVAL_23 = _EVAL_95;
  assign _EVAL_75 = _EVAL_70;
  assign _EVAL_225 = _EVAL_195 | _EVAL_156;
  assign _EVAL_268 = _EVAL_60 ^ 30'h2000;
  assign _EVAL_272 = {_EVAL_8,2'h0,_EVAL_130,_EVAL_100,2'h0,_EVAL_62,1'h0};
  assign _EVAL_177 = 23'hff << _EVAL_37;
  assign _EVAL_119 = _EVAL_264 | _EVAL_240;
  assign _EVAL_105 = _EVAL_7;
  assign _EVAL_141 = _EVAL_171 - _EVAL_131;
  assign _EVAL_123 = _EVAL_168 | _EVAL_200;
  assign _EVAL_276 = _EVAL_224;
  assign _EVAL_88 = _EVAL_90[1:0];
  assign _EVAL_93 = _EVAL_110;
  assign _EVAL_67 = _EVAL_60[11:0];
  assign _EVAL_261 = _EVAL_149 | _EVAL_259;
  assign _EVAL_187 = _EVAL_60 ^ 30'h4000;
  assign _EVAL_165 = _EVAL_233 ? _EVAL_132 : 47'h0;
  assign _EVAL_136 = _EVAL_226 ? _EVAL_245 : _EVAL_212;
  assign _EVAL_274 = {_EVAL_73,2'h0,_EVAL_243,_EVAL_98,2'h0,_EVAL_55,1'h0};
  assign _EVAL_178 = _EVAL_205 | _EVAL_279;
  assign _EVAL_89 = _EVAL_12;
  assign _EVAL_203 = _EVAL_153[4:0];
  assign _EVAL_206 = _EVAL_275 ? _EVAL_148 : 47'h0;
  assign _EVAL_9 = _EVAL_90;
  assign _EVAL_113 = _EVAL_39;
  assign _EVAL_149 = _EVAL_241 & _EVAL_107;
  assign _EVAL_69 = _EVAL_235[34];
  assign _EVAL_76 = _EVAL_39;
  assign _EVAL_197 = {{2'd0}, _EVAL_262};
  assign _EVAL_215 = _EVAL_185 & _EVAL_155;
  assign _EVAL_233 = _EVAL_226 ? _EVAL_242 : _EVAL_248;
  assign _EVAL_111 = _EVAL_61 & _EVAL_146;
  assign _EVAL_262 = _EVAL_183[9:2];
  assign _EVAL_59 = _EVAL_12;
  assign _EVAL_138 = $signed(_EVAL_255) & 31'sh22006000;
  assign _EVAL_49 = _EVAL_95;
  assign _EVAL_153 = {_EVAL_179, 2'h0};
  assign _EVAL_174 = _EVAL_40 & _EVAL_137;
  assign _EVAL_51 = _EVAL_61 & _EVAL_246;
  assign _EVAL_152 = _EVAL_212 & _EVAL_80;
  assign _EVAL_92 = _EVAL_70;
  assign _EVAL_150 = _EVAL_184 | _EVAL_80;
  assign _EVAL_66 = _EVAL_166 | _EVAL_208;
  assign _EVAL_194 = _EVAL_209[9:5];
  assign _EVAL_140 = _EVAL_158[4];
  assign _EVAL_122 = {1'b0,$signed(_EVAL_162)};
  assign _EVAL_47 = _EVAL_70;
  assign _EVAL_246 = $signed(_EVAL_258) == 31'sh0;
  assign _EVAL_115 = _EVAL_7;
  assign _EVAL_263 = _EVAL_158 & _EVAL_217;
  assign _EVAL_162 = _EVAL_60 ^ 30'h2000000;
  assign _EVAL_13 = _EVAL_40 & _EVAL_270;
  assign _EVAL_56 = _EVAL_39;
  assign _EVAL_198 = _EVAL_217 & _EVAL_143;
  assign _EVAL_175 = _EVAL_179 | _EVAL_203;
  assign _EVAL_64 = _EVAL_7;
  assign _EVAL_257 = _EVAL_225 | _EVAL_206;
  assign _EVAL_243 = {{2'd0}, _EVAL_46};
  assign _EVAL_85 = _EVAL_70;
  assign _EVAL_38 = _EVAL_235[41:38];
  assign _EVAL_167 = _EVAL_205[9:4];
  assign _EVAL_202 = $signed(_EVAL_176) == 31'sh0;
  assign _EVAL_184 = _EVAL_124 | _EVAL_106;
  assign _EVAL_255 = {1'b0,$signed(_EVAL_266)};
  assign _EVAL_217 = {_EVAL_80,_EVAL_106,_EVAL_71,_EVAL_96,_EVAL_107};
  assign _EVAL_250 = _EVAL_158[2];
  assign _EVAL_84 = _EVAL_40 & _EVAL_147;
  assign _EVAL_208 = _EVAL_193 & _EVAL_30;
  assign _EVAL_159 = {{1'd0}, _EVAL_204};
  assign _EVAL_227 = {{2'd0}, _EVAL_11};
  assign _EVAL_209 = _EVAL_159 | _EVAL_267;
  assign _EVAL_156 = _EVAL_133 ? _EVAL_274 : 47'h0;
  assign _EVAL_185 = _EVAL_226 & _EVAL_40;
  assign _EVAL_163 = ~_EVAL_142;
  assign _EVAL_16 = _EVAL_110;
  assign _EVAL_168 = _EVAL_192 | _EVAL_222;
  assign _EVAL_223 = {_EVAL_28,_EVAL_3,_EVAL_37,_EVAL_2,_EVAL_57,_EVAL_17,_EVAL_104,_EVAL_5};
  assign _EVAL_181 = _EVAL_226 ? _EVAL_118 : _EVAL_252;
  assign _EVAL_269 = _EVAL_107 | _EVAL_96;
  assign _EVAL_148 = {_EVAL_21,_EVAL_52,_EVAL_227,_EVAL_45,_EVAL_91,_EVAL_58,_EVAL_1,_EVAL_63};
  assign _EVAL_238 = {1'b0,$signed(_EVAL_187)};
  assign _EVAL_144 = _EVAL_226 ? _EVAL_250 : _EVAL_164;
  assign _EVAL_131 = {{5'd0}, _EVAL_174};
  assign _EVAL = _EVAL_70;
  assign _EVAL_271 = {1'b0,$signed(_EVAL_60)};
  assign _EVAL_195 = _EVAL_120 | _EVAL_165;
  assign _EVAL_180 = _EVAL_226 ? _EVAL_260 : _EVAL_241;
  assign _EVAL_118 = _EVAL_158[3];
  assign _EVAL_121 = _EVAL_154[9:1];
  assign _EVAL_235 = _EVAL_257 | _EVAL_254;
  assign _EVAL_0 = _EVAL_61 & _EVAL_127;
  assign _EVAL_240 = _EVAL_252 & _EVAL_106;
  assign _EVAL_130 = {{2'd0}, _EVAL_99};
  assign _EVAL_33 = _EVAL_7;
  assign _EVAL_189 = $signed(_EVAL_207) & 31'sh22006000;
  assign _EVAL_196 = $signed(_EVAL_271) & 31'sh22006000;
  assign _EVAL_265 = _EVAL_119 | _EVAL_152;
  assign _EVAL_109 = _EVAL_39;
  assign _EVAL_193 = $signed(_EVAL_276) == 31'sh0;
  assign _EVAL_54 = _EVAL_12;
  assign _EVAL_134 = _EVAL_226 ? _EVAL_237 : _EVAL_241;
  assign _EVAL_146 = $signed(_EVAL_218) == 31'sh0;
  assign _EVAL_270 = _EVAL_226 ? _EVAL_234 : _EVAL_248;
  assign _EVAL_158 = ~_EVAL_190;
  assign _EVAL_218 = _EVAL_189;
  assign _EVAL_24 = _EVAL_7;
  assign _EVAL_143 = ~_EVAL_253;
  assign _EVAL_207 = {1'b0,$signed(_EVAL_268)};
  assign _EVAL_234 = _EVAL_158[1];
  assign _EVAL_182 = _EVAL_127 & _EVAL_101;
  assign _EVAL_29 = _EVAL_40 & _EVAL_181;
  assign _EVAL_258 = _EVAL_196;
  assign _EVAL_124 = _EVAL_269 | _EVAL_71;
  assign _EVAL_27 = _EVAL_61 & _EVAL_202;
  assign _EVAL_264 = _EVAL_261 | _EVAL_116;
  assign _EVAL_31 = _EVAL_20;
  assign _EVAL_32 = _EVAL_90[1:0];
  assign _EVAL_183 = _EVAL_154 | _EVAL_247;
  assign _EVAL_147 = _EVAL_226 ? _EVAL_140 : _EVAL_212;
  assign _EVAL_256 = {_EVAL_263, 1'h0};
  assign _EVAL_169 = _EVAL_138;
  assign _EVAL_224 = $signed(_EVAL_238) & 31'sh22006000;
  assign _EVAL_48 = _EVAL_108;
  assign _EVAL_157 = _EVAL_141[5:0];
  assign _EVAL_132 = {_EVAL_14,2'h0,_EVAL_213,_EVAL_19,2'h0,_EVAL_114,1'h0};
  assign _EVAL_43 = _EVAL_60[14:0];
  assign _EVAL_210 = _EVAL_163[7:2];
  assign _EVAL_10 = _EVAL_226 ? _EVAL_150 : _EVAL_265;
  assign _EVAL_251 = _EVAL_250 & _EVAL_71;
  assign _EVAL_155 = _EVAL_217 != 5'h0;
  assign _EVAL_259 = _EVAL_248 & _EVAL_96;
  assign _EVAL_213 = {{2'd0}, _EVAL_77};
  assign _EVAL_142 = _EVAL_177[7:0];
  assign _EVAL_176 = _EVAL_211;
  assign _EVAL_260 = _EVAL_158[0];
  assign _EVAL_204 = _EVAL_178[9:1];
  assign _EVAL_192 = _EVAL_146 & _EVAL_35;
  assign _EVAL_18 = _EVAL_61 & _EVAL_193;
  assign _EVAL_137 = _EVAL_226 ? _EVAL_150 : _EVAL_265;
  assign _EVAL_97 = _EVAL_95;
  assign _EVAL_41 = _EVAL_60;
  assign _EVAL_83 = _EVAL_12;
  assign _EVAL_65 = _EVAL_40 & _EVAL_180;
  assign _EVAL_267 = {_EVAL_253, 5'h0};
  assign _EVAL_34 = _EVAL_90[1:0];
  assign _EVAL_266 = _EVAL_60 ^ 30'h20000000;
  assign _EVAL_50 = _EVAL_235[43:42];
  assign _EVAL_279 = {{4'd0}, _EVAL_167};
  assign _EVAL_151 = _EVAL_28[0];
  assign _EVAL_116 = _EVAL_164 & _EVAL_71;
  assign _EVAL_222 = _EVAL_202 & _EVAL_53;
  assign _EVAL_179 = _EVAL_263 | _EVAL_125;
  assign _EVAL_200 = _EVAL_246 & _EVAL_87;
  assign _EVAL_103 = _EVAL_110;
  assign _EVAL_275 = _EVAL_226 ? _EVAL_161 : _EVAL_252;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_164 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_171 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_212 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_241 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_248 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_252 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_253 = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_79) begin
    if (_EVAL_86) begin
      _EVAL_164 <= 1'h0;
    end else if (_EVAL_226) begin
      _EVAL_164 <= _EVAL_251;
    end
    if (_EVAL_86) begin
      _EVAL_171 <= 6'h0;
    end else if (_EVAL_185) begin
      if (_EVAL_237) begin
        if (_EVAL_151) begin
          _EVAL_171 <= _EVAL_210;
        end else begin
          _EVAL_171 <= 6'h0;
        end
      end else begin
        _EVAL_171 <= 6'h0;
      end
    end else begin
      _EVAL_171 <= _EVAL_157;
    end
    if (_EVAL_86) begin
      _EVAL_212 <= 1'h0;
    end else if (_EVAL_226) begin
      _EVAL_212 <= _EVAL_245;
    end
    if (_EVAL_86) begin
      _EVAL_241 <= 1'h0;
    end else if (_EVAL_226) begin
      _EVAL_241 <= _EVAL_237;
    end
    if (_EVAL_86) begin
      _EVAL_248 <= 1'h0;
    end else if (_EVAL_226) begin
      _EVAL_248 <= _EVAL_242;
    end
    if (_EVAL_86) begin
      _EVAL_252 <= 1'h0;
    end else if (_EVAL_226) begin
      _EVAL_252 <= _EVAL_161;
    end
    if (_EVAL_86) begin
      _EVAL_253 <= 5'h1f;
    end else if (_EVAL_215) begin
      _EVAL_253 <= _EVAL_128;
    end
  end
endmodule
