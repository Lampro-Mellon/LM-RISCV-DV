//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_161_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [31:0] _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [3:0]  _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [1:0]  _EVAL_13,
  input         _EVAL_14,
  input  [3:0]  _EVAL_15,
  input         _EVAL_16,
  input  [2:0]  _EVAL_17,
  input  [3:0]  _EVAL_18
);
  wire  _EVAL_19;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire [6:0] _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire [5:0] _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire [32:0] _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire [7:0] _EVAL_46;
  wire  _EVAL_47;
  wire [6:0] _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire [32:0] _EVAL_56;
  wire [32:0] _EVAL_57;
  wire  _EVAL_58;
  wire [5:0] _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_62;
  wire [31:0] _EVAL_63;
  wire  _EVAL_64;
  wire [7:0] _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire [1:0] _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  reg [5:0] _EVAL_81;
  reg [31:0] _RAND_0;
  wire  _EVAL_82;
  wire [22:0] _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  reg [5:0] _EVAL_89;
  reg [31:0] _RAND_1;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire [32:0] _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire [31:0] _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  reg [5:0] _EVAL_103;
  reg [31:0] _RAND_2;
  wire [1:0] _EVAL_105;
  wire  _EVAL_107;
  wire  _EVAL_108;
  reg [5:0] _EVAL_109;
  reg [31:0] _RAND_3;
  wire [32:0] _EVAL_110;
  wire [31:0] _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  reg [2:0] _EVAL_118;
  reg [31:0] _RAND_4;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  reg [2:0] _EVAL_127;
  reg [31:0] _RAND_5;
  wire [1:0] _EVAL_128;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire [3:0] _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire [1:0] _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [5:0] _EVAL_143;
  reg [3:0] _EVAL_144;
  reg [31:0] _RAND_6;
  wire  _EVAL_145;
  wire [32:0] _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire [32:0] _EVAL_151;
  wire  _EVAL_152;
  wire [32:0] _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire [1:0] _EVAL_157;
  wire  _EVAL_158;
  reg  _EVAL_159;
  reg [31:0] _RAND_7;
  wire  _EVAL_160;
  wire  _EVAL_161;
  reg [31:0] _EVAL_162;
  reg [31:0] _RAND_8;
  wire [7:0] _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire [32:0] _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire [32:0] _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire [3:0] _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  reg [2:0] _EVAL_181;
  reg [31:0] _RAND_9;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire [7:0] _EVAL_186;
  wire [32:0] _EVAL_187;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire [5:0] _EVAL_198;
  reg  _EVAL_199;
  reg [31:0] _RAND_10;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire [1:0] _EVAL_202;
  reg [1:0] _EVAL_203;
  reg [31:0] _RAND_11;
  wire [1:0] _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire [5:0] _EVAL_216;
  wire  _EVAL_217;
  reg  _EVAL_218;
  reg [31:0] _RAND_12;
  wire  _EVAL_219;
  wire [5:0] _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire [32:0] _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire [6:0] _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire [1:0] _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire [31:0] _EVAL_238;
  wire [31:0] _EVAL_239;
  wire  _EVAL_240;
  wire [32:0] _EVAL_242;
  wire [6:0] _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  reg [1:0] _EVAL_246;
  reg [31:0] _RAND_13;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire [32:0] _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  reg  _EVAL_253;
  reg [31:0] _RAND_14;
  wire  _EVAL_254;
  wire [1:0] _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire [31:0] _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire [3:0] _EVAL_268;
  wire [31:0] _EVAL_269;
  wire  _EVAL_270;
  wire [32:0] _EVAL_271;
  wire  _EVAL_272;
  wire [32:0] _EVAL_273;
  wire  _EVAL_274;
  reg [3:0] _EVAL_275;
  reg [31:0] _RAND_15;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire [31:0] _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire [22:0] _EVAL_283;
  wire  _EVAL_284;
  wire [32:0] _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_288;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire [32:0] _EVAL_296;
  wire [1:0] _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire [1:0] _EVAL_301;
  reg [31:0] _EVAL_302;
  reg [31:0] _RAND_16;
  wire  _EVAL_303;
  wire [1:0] _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_314;
  wire [3:0] _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire  _EVAL_321;
  wire  _EVAL_322;
  wire  _EVAL_323;
  wire  _EVAL_324;
  wire [32:0] _EVAL_325;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_116 = _EVAL_18 == _EVAL_275;
  assign _EVAL_191 = ~_EVAL_130;
  assign _EVAL_23 = $signed(_EVAL_296) == 33'sh0;
  assign _EVAL_69 = _EVAL_17 == _EVAL_181;
  assign _EVAL_170 = _EVAL_12 == 3'h1;
  assign _EVAL_40 = _EVAL_277 | _EVAL_14;
  assign _EVAL_145 = _EVAL_209 | _EVAL_29;
  assign _EVAL_76 = 2'h1 << _EVAL_7;
  assign _EVAL_38 = ~_EVAL_185;
  assign _EVAL_78 = _EVAL_8 & _EVAL_147;
  assign _EVAL_83 = 23'hff << _EVAL_18;
  assign _EVAL_138 = _EVAL_12 == 3'h0;
  assign _EVAL_90 = _EVAL_55 & _EVAL_149;
  assign _EVAL_142 = ~_EVAL_88;
  assign _EVAL_262 = _EVAL_5 ^ 32'h80000000;
  assign _EVAL_284 = ~_EVAL_49;
  assign _EVAL_205 = ~_EVAL_293;
  assign _EVAL_140 = _EVAL_148 | _EVAL_14;
  assign _EVAL_163 = _EVAL_83[7:0];
  assign _EVAL_292 = _EVAL_8 & _EVAL_231;
  assign _EVAL_155 = _EVAL_81 == 6'h0;
  assign _EVAL_52 = _EVAL_101 | _EVAL_299;
  assign _EVAL_168 = {1'b0,$signed(_EVAL_269)};
  assign _EVAL_268 = ~_EVAL_134;
  assign _EVAL_270 = _EVAL_255 != 2'h0;
  assign _EVAL_84 = _EVAL_161 | _EVAL_14;
  assign _EVAL_86 = ~_EVAL_31;
  assign _EVAL_94 = _EVAL_103 == 6'h0;
  assign _EVAL_294 = _EVAL_190 | _EVAL_14;
  assign _EVAL_227 = _EVAL_17 != 3'h0;
  assign _EVAL_222 = _EVAL_315 == 4'h0;
  assign _EVAL_122 = ~_EVAL_221;
  assign _EVAL_33 = _EVAL_244 & _EVAL_95;
  assign _EVAL_34 = ~_EVAL_120;
  assign _EVAL_248 = _EVAL_1 == _EVAL_199;
  assign _EVAL_58 = ~_EVAL_306;
  assign _EVAL_190 = _EVAL == _EVAL_253;
  assign _EVAL_258 = _EVAL_322 | _EVAL_90;
  assign _EVAL_318 = _EVAL_139 & _EVAL_155;
  assign _EVAL_66 = ~_EVAL_260;
  assign _EVAL_215 = ~_EVAL_172;
  assign _EVAL_228 = _EVAL_10 == _EVAL_134;
  assign _EVAL_288 = ~_EVAL_240;
  assign _EVAL_264 = ~_EVAL_40;
  assign _EVAL_75 = _EVAL_301[0];
  assign _EVAL_240 = _EVAL_80 | _EVAL_14;
  assign _EVAL_143 = _EVAL_243[5:0];
  assign _EVAL_308 = ~_EVAL_272;
  assign _EVAL_166 = _EVAL_7 == _EVAL_218;
  assign _EVAL_153 = $signed(_EVAL_285) & -33'sh1000000;
  assign _EVAL_151 = {1'b0,$signed(_EVAL_262)};
  assign _EVAL_255 = _EVAL_169 ? _EVAL_76 : 2'h0;
  assign _EVAL_124 = ~_EVAL_87;
  assign _EVAL_283 = 23'hff << _EVAL_15;
  assign _EVAL_232 = _EVAL_13 == _EVAL_203;
  assign _EVAL_236 = _EVAL_112 | _EVAL_14;
  assign _EVAL_311 = _EVAL_18 >= 4'h2;
  assign _EVAL_179 = _EVAL_9 == 3'h4;
  assign _EVAL_114 = _EVAL_115 & _EVAL_108;
  assign _EVAL_206 = _EVAL_246 != 2'h0;
  assign _EVAL_24 = _EVAL_67 & _EVAL_35;
  assign _EVAL_224 = _EVAL_116 | _EVAL_14;
  assign _EVAL_323 = ~_EVAL_99;
  assign _EVAL_167 = _EVAL_180 | _EVAL_90;
  assign _EVAL_93 = ~_EVAL_14;
  assign _EVAL_73 = _EVAL_0 & _EVAL_249;
  assign _EVAL_42 = ~_EVAL_140;
  assign _EVAL_107 = _EVAL_15 >= 4'h2;
  assign _EVAL_303 = _EVAL_0 & _EVAL_320;
  assign _EVAL_172 = _EVAL_9[2];
  assign _EVAL_47 = _EVAL_41 | _EVAL_214;
  assign _EVAL_67 = _EVAL_15 <= 4'h2;
  assign _EVAL_319 = _EVAL_207 | _EVAL_114;
  assign _EVAL_156 = _EVAL_109 == 6'h0;
  assign _EVAL_59 = _EVAL_48[5:0];
  assign _EVAL_296 = _EVAL_271;
  assign _EVAL_197 = _EVAL_8 & _EVAL_251;
  assign _EVAL_146 = _EVAL_173;
  assign _EVAL_50 = _EVAL_227 | _EVAL_14;
  assign _EVAL_37 = _EVAL_58 | _EVAL_14;
  assign _EVAL_272 = _EVAL_126 | _EVAL_14;
  assign _EVAL_247 = _EVAL_26 | _EVAL_14;
  assign _EVAL_314 = ~_EVAL_224;
  assign _EVAL_97 = $signed(_EVAL_56) & -33'sh2000;
  assign _EVAL_226 = _EVAL_0 & _EVAL_43;
  assign _EVAL_117 = _EVAL_13 <= 2'h2;
  assign _EVAL_290 = _EVAL_67 & _EVAL_145;
  assign _EVAL_41 = _EVAL_255 != _EVAL_297;
  assign _EVAL_157 = _EVAL_246 >> _EVAL_7;
  assign _EVAL_325 = {1'b0,$signed(_EVAL_5)};
  assign _EVAL_48 = _EVAL_109 - 6'h1;
  assign _EVAL_276 = $signed(_EVAL_250) == 33'sh0;
  assign _EVAL_271 = $signed(_EVAL_168) & -33'sh2000;
  assign _EVAL_279 = _EVAL_167 | _EVAL_14;
  assign _EVAL_249 = _EVAL_12 == 3'h2;
  assign _EVAL_266 = _EVAL_15 <= 4'h6;
  assign _EVAL_126 = _EVAL_211 | _EVAL_177;
  assign _EVAL_244 = _EVAL_204[1];
  assign _EVAL_238 = _EVAL_5 ^ 32'h2000000;
  assign _EVAL_291 = ~_EVAL_30;
  assign _EVAL_115 = _EVAL_204[0];
  assign _EVAL_105 = _EVAL_255 | _EVAL_246;
  assign _EVAL_149 = $signed(_EVAL_36) == 33'sh0;
  assign _EVAL_219 = ~_EVAL_37;
  assign _EVAL_280 = _EVAL_110[31:0];
  assign _EVAL_137 = _EVAL_246 | _EVAL_255;
  assign _EVAL_200 = _EVAL_82 | _EVAL_276;
  assign _EVAL_49 = _EVAL_12 == 3'h6;
  assign _EVAL_27 = _EVAL_89 - 6'h1;
  assign _EVAL_178 = _EVAL_10 & _EVAL_268;
  assign _EVAL_254 = _EVAL_8 & _EVAL_176;
  assign _EVAL_193 = _EVAL_17 <= 3'h1;
  assign _EVAL_79 = _EVAL_274 | _EVAL_189;
  assign _EVAL_147 = _EVAL_9 == 3'h1;
  assign _EVAL_261 = ~_EVAL_95;
  assign _EVAL_301 = _EVAL_105 >> _EVAL_1;
  assign _EVAL_43 = _EVAL_12 == 3'h5;
  assign _EVAL_112 = _EVAL_15 == _EVAL_144;
  assign _EVAL_134 = {_EVAL_79,_EVAL_39,_EVAL_319,_EVAL_237};
  assign _EVAL_324 = _EVAL_3 == _EVAL_159;
  assign _EVAL_312 = ~_EVAL_132;
  assign _EVAL_282 = ~_EVAL_307;
  assign _EVAL_91 = _EVAL_9 == 3'h2;
  assign _EVAL_243 = _EVAL_103 - 6'h1;
  assign _EVAL_251 = _EVAL_9 == 3'h6;
  assign _EVAL_185 = _EVAL_228 | _EVAL_14;
  assign _EVAL_164 = _EVAL_15[0];
  assign _EVAL_53 = _EVAL_8 & _EVAL_265;
  assign _EVAL_141 = _EVAL_152 | _EVAL_14;
  assign _EVAL_285 = {1'b0,$signed(_EVAL_238)};
  assign _EVAL_242 = $signed(_EVAL_273) & -33'sh1000;
  assign _EVAL_87 = _EVAL_311 | _EVAL_14;
  assign _EVAL_225 = _EVAL_97;
  assign _EVAL_305 = ~_EVAL_11;
  assign _EVAL_55 = _EVAL_15 <= 4'h8;
  assign _EVAL_44 = ~_EVAL_155;
  assign _EVAL_123 = _EVAL_5 == _EVAL_302;
  assign _EVAL_177 = _EVAL_67 & _EVAL_29;
  assign _EVAL_201 = _EVAL_111 == 32'h0;
  assign _EVAL_131 = _EVAL_266 & _EVAL_23;
  assign _EVAL_158 = _EVAL_8 & _EVAL_44;
  assign _EVAL_92 = _EVAL_123 | _EVAL_14;
  assign _EVAL_121 = _EVAL_54 | _EVAL_14;
  assign _EVAL_102 = ~_EVAL_235;
  assign _EVAL_45 = ~_EVAL_156;
  assign _EVAL_88 = _EVAL_258 | _EVAL_14;
  assign _EVAL_277 = _EVAL_212 | _EVAL_11;
  assign _EVAL_196 = ~_EVAL_252;
  assign _EVAL_304 = 2'h1 << _EVAL_1;
  assign _EVAL_250 = _EVAL_187;
  assign _EVAL_120 = _EVAL_193 | _EVAL_14;
  assign _EVAL_25 = ~_EVAL_195;
  assign _EVAL_119 = ~_EVAL_300;
  assign _EVAL_194 = _EVAL_28 & _EVAL_284;
  assign _EVAL_70 = _EVAL_8 & _EVAL_91;
  assign _EVAL_300 = _EVAL_222 | _EVAL_14;
  assign _EVAL_315 = ~_EVAL_10;
  assign _EVAL_204 = _EVAL_234 | 2'h1;
  assign _EVAL_216 = _EVAL_27[5:0];
  assign _EVAL_202 = ~_EVAL_297;
  assign _EVAL_26 = _EVAL_178 == 4'h0;
  assign _EVAL_223 = _EVAL_139 | _EVAL_68;
  assign _EVAL_128 = _EVAL_137 & _EVAL_202;
  assign _EVAL_135 = ~_EVAL_236;
  assign _EVAL_316 = ~_EVAL_84;
  assign _EVAL_111 = _EVAL_5 & _EVAL_63;
  assign _EVAL_154 = _EVAL_0 & _EVAL_170;
  assign _EVAL_175 = $signed(_EVAL_146) == 33'sh0;
  assign _EVAL_214 = ~_EVAL_270;
  assign _EVAL_99 = _EVAL_305 | _EVAL_14;
  assign _EVAL_256 = _EVAL_115 & _EVAL_267;
  assign _EVAL_306 = _EVAL_157[0];
  assign _EVAL_184 = _EVAL_9 == 3'h5;
  assign _EVAL_307 = _EVAL_75 | _EVAL_14;
  assign _EVAL_207 = _EVAL_107 | _EVAL_245;
  assign _EVAL_310 = _EVAL_0 & _EVAL_49;
  assign _EVAL_65 = ~_EVAL_46;
  assign _EVAL_320 = _EVAL_12 == 3'h4;
  assign _EVAL_317 = ~_EVAL_247;
  assign _EVAL_110 = _EVAL_162 + 32'h1;
  assign _EVAL_72 = _EVAL_17 == 3'h0;
  assign _EVAL_169 = _EVAL_139 & _EVAL_60;
  assign _EVAL_210 = _EVAL_212 | _EVAL_14;
  assign _EVAL_220 = _EVAL_65[7:2];
  assign _EVAL_35 = _EVAL_200 | _EVAL_29;
  assign _EVAL_195 = _EVAL_107 | _EVAL_14;
  assign _EVAL_63 = {{24'd0}, _EVAL_65};
  assign _EVAL_260 = _EVAL_248 | _EVAL_14;
  assign _EVAL_237 = _EVAL_207 | _EVAL_256;
  assign _EVAL_113 = ~_EVAL_121;
  assign _EVAL_180 = _EVAL_67 & _EVAL_200;
  assign _EVAL_183 = _EVAL_47 | _EVAL_14;
  assign _EVAL_60 = _EVAL_89 == 6'h0;
  assign _EVAL_108 = _EVAL_261 & _EVAL_233;
  assign _EVAL_160 = ~_EVAL_183;
  assign _EVAL_321 = _EVAL_115 & _EVAL_259;
  assign _EVAL_85 = ~_EVAL_294;
  assign _EVAL_161 = _EVAL_17 <= 3'h2;
  assign _EVAL_267 = _EVAL_261 & _EVAL_182;
  assign _EVAL_100 = _EVAL_5 ^ 32'h20000000;
  assign _EVAL_96 = ~_EVAL_217;
  assign _EVAL_187 = $signed(_EVAL_325) & -33'sh5000;
  assign _EVAL_245 = _EVAL_244 & _EVAL_261;
  assign _EVAL_71 = _EVAL_95 & _EVAL_233;
  assign _EVAL_173 = $signed(_EVAL_151) & -33'shc000;
  assign _EVAL_186 = ~_EVAL_163;
  assign _EVAL_132 = _EVAL_69 | _EVAL_14;
  assign _EVAL_322 = _EVAL_24 | _EVAL_131;
  assign _EVAL_252 = _EVAL_166 | _EVAL_14;
  assign _EVAL_101 = ~_EVAL_206;
  assign _EVAL_217 = _EVAL_117 | _EVAL_14;
  assign _EVAL_56 = {1'b0,$signed(_EVAL_100)};
  assign _EVAL_234 = 2'h1 << _EVAL_164;
  assign _EVAL_31 = _EVAL_72 | _EVAL_14;
  assign _EVAL_139 = _EVAL_4 & _EVAL_8;
  assign _EVAL_269 = _EVAL_5 ^ 32'h40000000;
  assign _EVAL_239 = _EVAL_5 ^ 32'h3000;
  assign _EVAL_278 = ~_EVAL_210;
  assign _EVAL_22 = _EVAL_162 < plusarg_reader_out;
  assign _EVAL_192 = _EVAL_0 & _EVAL_138;
  assign _EVAL_51 = _EVAL_8 & _EVAL_184;
  assign _EVAL_230 = _EVAL_81 - 6'h1;
  assign _EVAL_281 = _EVAL_229 | _EVAL_14;
  assign _EVAL_30 = _EVAL_290 | _EVAL_14;
  assign _EVAL_229 = _EVAL_17 <= 3'h3;
  assign _EVAL_36 = _EVAL_242;
  assign _EVAL_29 = $signed(_EVAL_225) == 33'sh0;
  assign _EVAL_57 = _EVAL_153;
  assign _EVAL_176 = _EVAL_9 == 3'h7;
  assign _EVAL_259 = _EVAL_95 & _EVAL_182;
  assign _EVAL_263 = ~_EVAL_281;
  assign _EVAL_82 = _EVAL_175 | _EVAL_21;
  assign _EVAL_231 = _EVAL_9 == 3'h0;
  assign _EVAL_309 = ~_EVAL_50;
  assign _EVAL_293 = _EVAL_232 | _EVAL_14;
  assign _EVAL_171 = ~_EVAL_279;
  assign _EVAL_257 = _EVAL_13 != 2'h2;
  assign _EVAL_152 = _EVAL_17 <= 3'h4;
  assign _EVAL_286 = _EVAL_12 <= 3'h6;
  assign _EVAL_297 = _EVAL_194 ? _EVAL_304 : 2'h0;
  assign _EVAL_189 = _EVAL_115 & _EVAL_71;
  assign _EVAL_221 = _EVAL_298 | _EVAL_14;
  assign _EVAL_21 = $signed(_EVAL_57) == 33'sh0;
  assign _EVAL_265 = _EVAL_9 == 3'h3;
  assign _EVAL_148 = _EVAL_9 == _EVAL_118;
  assign _EVAL_136 = _EVAL_201 | _EVAL_14;
  assign _EVAL_299 = plusarg_reader_out == 32'h0;
  assign _EVAL_74 = ~_EVAL_92;
  assign _EVAL_95 = _EVAL_5[1];
  assign _EVAL_165 = _EVAL_149 | _EVAL_21;
  assign _EVAL_77 = _EVAL_8 & _EVAL_179;
  assign _EVAL_298 = _EVAL_13 == 2'h0;
  assign _EVAL_274 = _EVAL_107 | _EVAL_33;
  assign _EVAL_174 = ~_EVAL_141;
  assign _EVAL_19 = _EVAL_68 & _EVAL_156;
  assign _EVAL_46 = _EVAL_283[7:0];
  assign _EVAL_208 = _EVAL_125 | _EVAL_14;
  assign _EVAL_28 = _EVAL_68 & _EVAL_94;
  assign _EVAL_198 = _EVAL_186[7:2];
  assign _EVAL_62 = ~_EVAL_98;
  assign _EVAL_273 = {1'b0,$signed(_EVAL_239)};
  assign _EVAL_295 = ~_EVAL_208;
  assign _EVAL_130 = _EVAL_324 | _EVAL_14;
  assign _EVAL_39 = _EVAL_274 | _EVAL_321;
  assign _EVAL_233 = _EVAL_5[0];
  assign _EVAL_68 = _EVAL_2 & _EVAL_0;
  assign _EVAL_212 = ~_EVAL;
  assign _EVAL_182 = ~_EVAL_233;
  assign _EVAL_32 = _EVAL_230[5:0];
  assign _EVAL_54 = _EVAL_52 | _EVAL_22;
  assign _EVAL_150 = ~_EVAL_136;
  assign _EVAL_80 = ~_EVAL_16;
  assign _EVAL_209 = _EVAL_165 | _EVAL_276;
  assign _EVAL_235 = _EVAL_257 | _EVAL_14;
  assign _EVAL_213 = _EVAL_12[0];
  assign _EVAL_98 = _EVAL_286 | _EVAL_14;
  assign _EVAL_125 = _EVAL_12 == _EVAL_127;
  assign _EVAL_211 = _EVAL_131 | _EVAL_90;
  assign _EVAL_64 = _EVAL_0 & _EVAL_45;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_81 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_89 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_103 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_109 = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_118 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_127 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_144 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_159 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_162 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_181 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_199 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_203 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_218 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_246 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_253 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_275 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_302 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_6) begin
    if (_EVAL_14) begin
      _EVAL_81 <= 6'h0;
    end else if (_EVAL_139) begin
      if (_EVAL_155) begin
        if (_EVAL_215) begin
          _EVAL_81 <= _EVAL_220;
        end else begin
          _EVAL_81 <= 6'h0;
        end
      end else begin
        _EVAL_81 <= _EVAL_32;
      end
    end
    if (_EVAL_14) begin
      _EVAL_89 <= 6'h0;
    end else if (_EVAL_139) begin
      if (_EVAL_60) begin
        if (_EVAL_215) begin
          _EVAL_89 <= _EVAL_220;
        end else begin
          _EVAL_89 <= 6'h0;
        end
      end else begin
        _EVAL_89 <= _EVAL_216;
      end
    end
    if (_EVAL_14) begin
      _EVAL_103 <= 6'h0;
    end else if (_EVAL_68) begin
      if (_EVAL_94) begin
        if (_EVAL_213) begin
          _EVAL_103 <= _EVAL_198;
        end else begin
          _EVAL_103 <= 6'h0;
        end
      end else begin
        _EVAL_103 <= _EVAL_143;
      end
    end
    if (_EVAL_14) begin
      _EVAL_109 <= 6'h0;
    end else if (_EVAL_68) begin
      if (_EVAL_156) begin
        if (_EVAL_213) begin
          _EVAL_109 <= _EVAL_198;
        end else begin
          _EVAL_109 <= 6'h0;
        end
      end else begin
        _EVAL_109 <= _EVAL_59;
      end
    end
    if (_EVAL_318) begin
      _EVAL_118 <= _EVAL_9;
    end
    if (_EVAL_19) begin
      _EVAL_127 <= _EVAL_12;
    end
    if (_EVAL_318) begin
      _EVAL_144 <= _EVAL_15;
    end
    if (_EVAL_19) begin
      _EVAL_159 <= _EVAL_3;
    end
    if (_EVAL_14) begin
      _EVAL_162 <= 32'h0;
    end else if (_EVAL_223) begin
      _EVAL_162 <= 32'h0;
    end else begin
      _EVAL_162 <= _EVAL_280;
    end
    if (_EVAL_318) begin
      _EVAL_181 <= _EVAL_17;
    end
    if (_EVAL_19) begin
      _EVAL_199 <= _EVAL_1;
    end
    if (_EVAL_19) begin
      _EVAL_203 <= _EVAL_13;
    end
    if (_EVAL_318) begin
      _EVAL_218 <= _EVAL_7;
    end
    if (_EVAL_14) begin
      _EVAL_246 <= 2'h0;
    end else begin
      _EVAL_246 <= _EVAL_128;
    end
    if (_EVAL_19) begin
      _EVAL_253 <= _EVAL;
    end
    if (_EVAL_19) begin
      _EVAL_275 <= _EVAL_18;
    end
    if (_EVAL_318) begin
      _EVAL_302 <= _EVAL_5;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_323) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed1fcdfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_288) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10395d21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_264) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f97f1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53f8b4ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54808202)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d323eef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_288) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7564c20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_323) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47d75383)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4869d365)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_308) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7640474b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_288) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4050bbf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_323) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8cac592)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(593ff283)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88f11629)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4193e8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3696a1e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_264) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e12309fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_323) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_264) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ec71618)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5eb026e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a860211b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d62da4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_308) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a472c296)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d35a190)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_288) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f37d84f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(297a8647)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_66) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_288) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1321e6b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6144ae9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8229ad03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53fae094)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bddd3c54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3936610)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d2a867c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_316) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_323) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55e6db90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c8aeb85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb0df290)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcbcaa3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e27a348)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3654ec09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1b5953b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_323) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c864f23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a13428c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5227d799)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(585c2b5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_66) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c53a0894)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5026ce7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9eda665)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3706179c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d206fd38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e15394a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d564188)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6e43cee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_323) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63f2648d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdeb743d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29cb37b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_288) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_264) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84d6f74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_316) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13d71d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8b3ba16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(641f1a03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_314) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_323) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9a6a59c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(beb51ed5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aeffdf1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbed5faf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8f2b7c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_316) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_316) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e128f09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5aa9e9f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_314) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90398261)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bae9eb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ca9913)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc11972)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43ec951)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_288) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d20ae72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_288) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2edaeba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d45c47e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(474cdd12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4033b189)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe5c0c36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b0630a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
