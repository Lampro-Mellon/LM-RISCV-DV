//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module SiFive_CoreIPSubsystem(
  input          clock,
  input          reset,
  output         halt_from_tile_0,
  output         wfi_from_tile_0,
  output         cease_from_tile_0,
  input          psd_test_clock_enable,
  input          meip_0,
  input          resetctrl_hartIsInReset_0,
  input          debug_clock,
  input          debug_reset,
  input          debug_systemjtag_jtag_TCK,
  input          debug_systemjtag_jtag_TMS,
  input          debug_systemjtag_jtag_TDI,
  output         debug_systemjtag_jtag_TDO_data,
  output         debug_systemjtag_jtag_TDO_driven,
  input          debug_systemjtag_reset,
  input  [10:0]  debug_systemjtag_mfr_id,
  input  [15:0]  debug_systemjtag_part_number,
  input  [3:0]   debug_systemjtag_version,
  output         debug_ndreset,
  output         debug_dmactive,
  input          debug_dmactiveAck,
  input  [31:0]  reset_vector_0,
  input          rtc_toggle,
  input  [126:0] local_interrupts_0,
  output         sys_port_ahb_0_hmastlock,
  input          sys_port_ahb_0_hready,
  output [1:0]   sys_port_ahb_0_htrans,
  output [2:0]   sys_port_ahb_0_hsize,
  output [2:0]   sys_port_ahb_0_hburst,
  output         sys_port_ahb_0_hwrite,
  output [3:0]   sys_port_ahb_0_hprot,
  output [30:0]  sys_port_ahb_0_haddr,
  output [31:0]  sys_port_ahb_0_hwdata,
  input          sys_port_ahb_0_hresp,
  input  [31:0]  sys_port_ahb_0_hrdata,
  output         periph_port_ahb_0_hmastlock,
  input          periph_port_ahb_0_hready,
  output [1:0]   periph_port_ahb_0_htrans,
  output [2:0]   periph_port_ahb_0_hsize,
  output [2:0]   periph_port_ahb_0_hburst,
  output         periph_port_ahb_0_hwrite,
  output [3:0]   periph_port_ahb_0_hprot,
  output [29:0]  periph_port_ahb_0_haddr,
  output [31:0]  periph_port_ahb_0_hwdata,
  input          periph_port_ahb_0_hresp,
  input  [31:0]  periph_port_ahb_0_hrdata,
  input          front_port_ahb_0_hmastlock,
  input          front_port_ahb_0_hsel,
  input          front_port_ahb_0_hready,
  output         front_port_ahb_0_hreadyout,
  input  [1:0]   front_port_ahb_0_htrans,
  input  [2:0]   front_port_ahb_0_hsize,
  input  [2:0]   front_port_ahb_0_hburst,
  input          front_port_ahb_0_hwrite,
  input  [3:0]   front_port_ahb_0_hprot,
  input  [31:0]  front_port_ahb_0_haddr,
  input  [31:0]  front_port_ahb_0_hwdata,
  output         front_port_ahb_0_hresp,
  output [31:0]  front_port_ahb_0_hrdata
);
  wire  testIndicator_auto_control_xing_in_a_ready;
  wire  testIndicator_auto_control_xing_in_a_valid;
  wire [2:0] testIndicator_auto_control_xing_in_a_bits_opcode;
  wire [2:0] testIndicator_auto_control_xing_in_a_bits_param;
  wire [1:0] testIndicator_auto_control_xing_in_a_bits_size;
  wire [2:0] testIndicator_auto_control_xing_in_a_bits_source;
  wire [14:0] testIndicator_auto_control_xing_in_a_bits_address;
  wire [3:0] testIndicator_auto_control_xing_in_a_bits_mask;
  wire [31:0] testIndicator_auto_control_xing_in_a_bits_data;
  wire  testIndicator_auto_control_xing_in_a_bits_corrupt;
  wire  testIndicator_auto_control_xing_in_d_ready;
  wire  testIndicator_auto_control_xing_in_d_valid;
  wire [2:0] testIndicator_auto_control_xing_in_d_bits_opcode;
  wire [1:0] testIndicator_auto_control_xing_in_d_bits_size;
  wire [2:0] testIndicator_auto_control_xing_in_d_bits_source;
  wire [31:0] testIndicator_auto_control_xing_in_d_bits_data;
  wire  testIndicator_clock;
  wire  testIndicator_reset;
  wire  xbar_1__EVAL;
  wire  xbar_1__EVAL_0;
  wire  xbar_2__EVAL;
  wire  xbar_2__EVAL_0;
  wire  _EVAL;
  wire  island__EVAL;
  wire [1:0] island__EVAL_0;
  wire [31:0] island__EVAL_1;
  wire  island__EVAL_2;
  wire  island__EVAL_3;
  wire  island__EVAL_4;
  wire [3:0] island__EVAL_5;
  wire  island__EVAL_6;
  wire  island__EVAL_7;
  wire [1:0] island__EVAL_8;
  wire [2:0] island__EVAL_9;
  wire [2:0] island__EVAL_10;
  wire [31:0] island__EVAL_11;
  wire  island__EVAL_12;
  wire [2:0] island__EVAL_13;
  wire [31:0] island__EVAL_14;
  wire [2:0] island__EVAL_15;
  wire [2:0] island__EVAL_16;
  wire  sbus__EVAL;
  wire  sbus__EVAL_0;
  wire [30:0] sbus__EVAL_1;
  wire [31:0] sbus__EVAL_2;
  wire [3:0] sbus__EVAL_3;
  wire [3:0] sbus__EVAL_4;
  wire [1:0] sbus__EVAL_5;
  wire [2:0] sbus__EVAL_6;
  wire  sbus__EVAL_7;
  wire  sbus__EVAL_8;
  wire  sbus__EVAL_9;
  wire [1:0] sbus__EVAL_10;
  wire [3:0] sbus__EVAL_11;
  wire [2:0] sbus__EVAL_12;
  wire [1:0] sbus__EVAL_13;
  wire  sbus__EVAL_14;
  wire [31:0] sbus__EVAL_15;
  wire  sbus__EVAL_16;
  wire  sbus__EVAL_17;
  wire  sbus__EVAL_18;
  wire  sbus__EVAL_19;
  wire  sbus__EVAL_20;
  wire [2:0] sbus__EVAL_21;
  wire  sbus__EVAL_23;
  wire  sbus__EVAL_24;
  wire [2:0] sbus__EVAL_25;
  wire [1:0] sbus__EVAL_26;
  wire [3:0] sbus__EVAL_27;
  wire  sbus__EVAL_28;
  wire  sbus__EVAL_29;
  wire [31:0] sbus__EVAL_30;
  wire  sbus__EVAL_31;
  wire [3:0] sbus__EVAL_32;
  wire [2:0] sbus__EVAL_33;
  wire  sbus__EVAL_34;
  wire  sbus__EVAL_36;
  wire  sbus__EVAL_37;
  wire [2:0] sbus__EVAL_38;
  wire  sbus__EVAL_39;
  wire [1:0] sbus__EVAL_41;
  wire [31:0] sbus__EVAL_42;
  wire  sbus__EVAL_43;
  wire [2:0] sbus__EVAL_44;
  wire  sbus__EVAL_45;
  wire  sbus__EVAL_46;
  wire [2:0] sbus__EVAL_47;
  wire  sbus__EVAL_48;
  wire  sbus__EVAL_50;
  wire  sbus__EVAL_51;
  wire [2:0] sbus__EVAL_52;
  wire  sbus__EVAL_53;
  wire  sbus__EVAL_54;
  wire  sbus__EVAL_55;
  wire [31:0] sbus__EVAL_56;
  wire [3:0] sbus__EVAL_57;
  wire [2:0] sbus__EVAL_58;
  wire  sbus__EVAL_59;
  wire  sbus__EVAL_60;
  wire  sbus__EVAL_61;
  wire  sbus__EVAL_62;
  wire  sbus__EVAL_63;
  wire [2:0] sbus__EVAL_64;
  wire [3:0] sbus__EVAL_65;
  wire [2:0] sbus__EVAL_66;
  wire [3:0] sbus__EVAL_67;
  wire  sbus__EVAL_68;
  wire  sbus__EVAL_69;
  wire [2:0] sbus__EVAL_70;
  wire  sbus__EVAL_71;
  wire  sbus__EVAL_72;
  wire [31:0] sbus__EVAL_73;
  wire  sbus__EVAL_74;
  wire  sbus__EVAL_76;
  wire  sbus__EVAL_77;
  wire  sbus__EVAL_78;
  wire [31:0] sbus__EVAL_79;
  wire [3:0] sbus__EVAL_80;
  wire  sbus__EVAL_81;
  wire  sbus__EVAL_82;
  wire  sbus__EVAL_83;
  wire  sbus__EVAL_84;
  wire  sbus__EVAL_85;
  wire [3:0] sbus__EVAL_86;
  wire [31:0] sbus__EVAL_87;
  wire [1:0] sbus__EVAL_89;
  wire [2:0] sbus__EVAL_90;
  wire  sbus__EVAL_91;
  wire  sbus__EVAL_92;
  wire  sbus__EVAL_93;
  wire [2:0] sbus__EVAL_94;
  wire  sbus__EVAL_95;
  wire  sbus__EVAL_96;
  wire  sbus__EVAL_97;
  wire [3:0] sbus__EVAL_98;
  wire [29:0] sbus__EVAL_99;
  wire  sbus__EVAL_100;
  wire  sbus__EVAL_101;
  wire [3:0] sbus__EVAL_102;
  wire  sbus__EVAL_103;
  wire [31:0] sbus__EVAL_104;
  wire  sbus__EVAL_105;
  wire [31:0] sbus__EVAL_106;
  wire  sbus__EVAL_107;
  wire [31:0] sbus__EVAL_108;
  wire [1:0] sbus__EVAL_109;
  wire  sbus__EVAL_110;
  wire [31:0] sbus__EVAL_111;
  wire [2:0] sbus__EVAL_112;
  wire  sbus__EVAL_113;
  wire  sbus__EVAL_114;
  wire [31:0] sbus__EVAL_115;
  wire [2:0] sbus__EVAL_116;
  wire  sbus__EVAL_117;
  wire [2:0] sbus__EVAL_118;
  wire [2:0] sbus__EVAL_119;
  wire  sbus__EVAL_120;
  wire  sbus__EVAL_121;
  wire  sbus__EVAL_122;
  wire [2:0] sbus__EVAL_123;
  wire [3:0] sbus__EVAL_124;
  wire [2:0] sbus__EVAL_125;
  wire [2:0] sbus__EVAL_126;
  wire [1:0] sbus__EVAL_128;
  wire  sbus__EVAL_129;
  wire  sbus__EVAL_130;
  wire  sbus__EVAL_131;
  wire [3:0] sbus__EVAL_132;
  wire  sbus__EVAL_133;
  wire  sbus__EVAL_134;
  wire  sbus__EVAL_135;
  wire  sbus__EVAL_136;
  wire  sbus__EVAL_137;
  wire  sbus__EVAL_138;
  wire  sbus__EVAL_139;
  wire  sbus__EVAL_140;
  wire  sbus__EVAL_141;
  wire  sbus__EVAL_142;
  wire  sbus__EVAL_143;
  wire  sbus__EVAL_144;
  wire [2:0] sbus__EVAL_146;
  wire [31:0] sbus__EVAL_147;
  wire [31:0] sbus__EVAL_148;
  wire [31:0] sbus__EVAL_150;
  wire [3:0] sbus__EVAL_151;
  wire [2:0] sbus__EVAL_152;
  wire  sbus__EVAL_153;
  wire [31:0] sbus__EVAL_154;
  wire  sbus__EVAL_156;
  wire  sbus__EVAL_157;
  wire  sbus__EVAL_158;
  wire  sbus__EVAL_159;
  wire  sbus__EVAL_160;
  wire [31:0] sbus__EVAL_161;
  wire [1:0] sbus__EVAL_162;
  wire [31:0] sbus__EVAL_164;
  wire  sbus__EVAL_165;
  wire [2:0] sbus__EVAL_167;
  wire [2:0] sbus__EVAL_168;
  wire  sbus__EVAL_169;
  wire  sbus__EVAL_170;
  wire  sbus__EVAL_171;
  reg  _EVAL_0;
  reg [31:0] _RAND_0;
  wire  SynchronizerShiftReg_w1_d3__EVAL;
  wire  SynchronizerShiftReg_w1_d3__EVAL_0;
  wire  SynchronizerShiftReg_w1_d3__EVAL_1;
  wire  _EVAL_1;
  wire [31:0] cbus__EVAL;
  wire  cbus__EVAL_0;
  wire [3:0] cbus__EVAL_1;
  wire [2:0] cbus__EVAL_2;
  wire  cbus__EVAL_3;
  wire  cbus__EVAL_4;
  wire [31:0] cbus__EVAL_7;
  wire [31:0] cbus__EVAL_8;
  wire [1:0] cbus__EVAL_9;
  wire [31:0] cbus__EVAL_10;
  wire  cbus__EVAL_11;
  wire  cbus__EVAL_12;
  wire [29:0] cbus__EVAL_13;
  wire [2:0] cbus__EVAL_14;
  wire [2:0] cbus__EVAL_15;
  wire  cbus__EVAL_16;
  wire [1:0] cbus__EVAL_17;
  wire  cbus__EVAL_18;
  wire [2:0] cbus__EVAL_19;
  wire [3:0] cbus__EVAL_20;
  wire [2:0] cbus__EVAL_21;
  wire [11:0] cbus__EVAL_22;
  wire  cbus__EVAL_23;
  wire  cbus__EVAL_24;
  wire [31:0] cbus__EVAL_25;
  wire [1:0] cbus__EVAL_26;
  wire [1:0] cbus__EVAL_27;
  wire  cbus__EVAL_28;
  wire [2:0] cbus__EVAL_29;
  wire [1:0] cbus__EVAL_30;
  wire  cbus__EVAL_31;
  wire [31:0] cbus__EVAL_32;
  wire [1:0] cbus__EVAL_34;
  wire  cbus__EVAL_35;
  wire  cbus__EVAL_36;
  wire [2:0] cbus__EVAL_37;
  wire  cbus__EVAL_38;
  wire  cbus__EVAL_39;
  wire  cbus__EVAL_40;
  wire [31:0] cbus__EVAL_41;
  wire  cbus__EVAL_42;
  wire  cbus__EVAL_43;
  wire [25:0] cbus__EVAL_44;
  wire [3:0] cbus__EVAL_45;
  wire [2:0] cbus__EVAL_46;
  wire [2:0] cbus__EVAL_47;
  wire [2:0] cbus__EVAL_48;
  wire [3:0] cbus__EVAL_49;
  wire [2:0] cbus__EVAL_50;
  wire [3:0] cbus__EVAL_51;
  wire  cbus__EVAL_52;
  wire [2:0] cbus__EVAL_54;
  wire [31:0] cbus__EVAL_55;
  wire  cbus__EVAL_56;
  wire  cbus__EVAL_57;
  wire [31:0] cbus__EVAL_58;
  wire  cbus__EVAL_59;
  wire  cbus__EVAL_60;
  wire [31:0] cbus__EVAL_61;
  wire [3:0] cbus__EVAL_62;
  wire  cbus__EVAL_63;
  wire [14:0] cbus__EVAL_64;
  wire [2:0] cbus__EVAL_65;
  wire [29:0] cbus__EVAL_66;
  wire  cbus__EVAL_67;
  wire [1:0] cbus__EVAL_68;
  wire [2:0] cbus__EVAL_69;
  wire  cbus__EVAL_70;
  wire  cbus__EVAL_71;
  wire [2:0] cbus__EVAL_72;
  wire  cbus__EVAL_73;
  wire [2:0] cbus__EVAL_74;
  wire  cbus__EVAL_75;
  wire [2:0] cbus__EVAL_76;
  wire  cbus__EVAL_77;
  wire  cbus__EVAL_78;
  wire [3:0] cbus__EVAL_79;
  wire  cbus__EVAL_80;
  wire [2:0] cbus__EVAL_81;
  wire [2:0] cbus__EVAL_82;
  wire  cbus__EVAL_83;
  wire  cbus__EVAL_84;
  wire [1:0] cbus__EVAL_85;
  wire  cbus__EVAL_86;
  wire [2:0] cbus__EVAL_87;
  wire  cbus__EVAL_88;
  wire [2:0] cbus__EVAL_89;
  wire  cbus__EVAL_90;
  wire  tile__EVAL;
  wire  tile__EVAL_0;
  wire [2:0] tile__EVAL_1;
  wire  tile__EVAL_2;
  wire  tile__EVAL_3;
  wire [7:0] tile__EVAL_4;
  wire [31:0] tile__EVAL_5;
  wire  tile__EVAL_6;
  wire  tile__EVAL_7;
  wire [31:0] tile__EVAL_8;
  wire  tile__EVAL_9;
  wire  tile__EVAL_10;
  wire  tile__EVAL_11;
  wire [3:0] tile__EVAL_12;
  wire  tile__EVAL_13;
  wire [7:0] tile__EVAL_14;
  wire  tile__EVAL_15;
  wire  tile__EVAL_16;
  wire [2:0] tile__EVAL_17;
  wire  tile__EVAL_18;
  wire  tile__EVAL_19;
  wire [31:0] tile__EVAL_20;
  wire  tile__EVAL_21;
  wire [3:0] tile__EVAL_22;
  wire  tile__EVAL_23;
  wire  tile__EVAL_24;
  wire  tile__EVAL_25;
  wire [31:0] tile__EVAL_26;
  wire  tile__EVAL_27;
  wire  tile__EVAL_28;
  wire  tile__EVAL_29;
  wire  tile__EVAL_30;
  wire  tile__EVAL_31;
  wire  tile__EVAL_32;
  wire  tile__EVAL_33;
  wire [2:0] tile__EVAL_34;
  wire  tile__EVAL_35;
  wire  tile__EVAL_36;
  wire  tile__EVAL_37;
  wire  tile__EVAL_38;
  wire [1:0] tile__EVAL_39;
  wire  tile__EVAL_40;
  wire  tile__EVAL_41;
  wire  tile__EVAL_42;
  wire [31:0] tile__EVAL_43;
  wire [1:0] tile__EVAL_44;
  wire [3:0] tile__EVAL_45;
  wire  tile__EVAL_46;
  wire [2:0] tile__EVAL_47;
  wire  tile__EVAL_48;
  wire [2:0] tile__EVAL_49;
  wire  tile__EVAL_50;
  wire  tile__EVAL_51;
  wire  tile__EVAL_52;
  wire  tile__EVAL_53;
  wire  tile__EVAL_54;
  wire  tile__EVAL_55;
  wire  tile__EVAL_56;
  wire  tile__EVAL_57;
  wire [3:0] tile__EVAL_58;
  wire [31:0] tile__EVAL_59;
  wire [3:0] tile__EVAL_60;
  wire [3:0] tile__EVAL_61;
  wire [2:0] tile__EVAL_62;
  wire  tile__EVAL_63;
  wire  tile__EVAL_64;
  wire  tile__EVAL_65;
  wire [31:0] tile__EVAL_66;
  wire  tile__EVAL_67;
  reg  _EVAL_2;
  reg [31:0] _RAND_1;
  wire  dummyClockGroupSourceNode__EVAL;
  wire  dummyClockGroupSourceNode__EVAL_0;
  wire  dummyClockGroupSourceNode__EVAL_1;
  wire  dummyClockGroupSourceNode__EVAL_2;
  wire  dummyClockGroupSourceNode__EVAL_3;
  wire  dummyClockGroupSourceNode__EVAL_8;
  wire  dummyClockGroupSourceNode__EVAL_11;
  wire  dummyClockGroupSourceNode__EVAL_12;
  wire [31:0] island_1__EVAL;
  wire [31:0] island_1__EVAL_0;
  wire [2:0] island_1__EVAL_1;
  wire [31:0] island_1__EVAL_2;
  wire  island_1__EVAL_3;
  wire  island_1__EVAL_4;
  wire  island_1__EVAL_5;
  wire  island_1__EVAL_6;
  wire  island_1__EVAL_7;
  wire [2:0] island_1__EVAL_8;
  wire [2:0] island_1__EVAL_9;
  wire [1:0] island_1__EVAL_10;
  wire [3:0] island_1__EVAL_11;
  wire [1:0] island_1__EVAL_12;
  wire [2:0] island_1__EVAL_13;
  wire  island_1__EVAL_14;
  wire [2:0] island_1__EVAL_15;
  wire  island_1__EVAL_16;
  wire  xbar__EVAL;
  wire  xbar__EVAL_0;
  wire [1:0] _EVAL_3;
  wire  dtm__EVAL;
  wire  dtm__EVAL_0;
  wire [6:0] dtm__EVAL_1;
  wire  dtm__EVAL_2;
  wire [31:0] dtm__EVAL_3;
  wire  dtm__EVAL_4;
  wire [3:0] dtm__EVAL_5;
  wire [15:0] dtm__EVAL_6;
  wire  dtm__EVAL_7;
  wire  dtm__EVAL_8;
  wire  dtm__EVAL_9;
  wire  dtm__EVAL_10;
  wire [1:0] dtm__EVAL_11;
  wire [31:0] dtm__EVAL_12;
  wire [10:0] dtm__EVAL_13;
  wire  dtm__EVAL_14;
  wire [1:0] dtm__EVAL_15;
  wire  dtm__EVAL_16;
  wire [2:0] debug_1__EVAL;
  wire  debug_1__EVAL_0;
  wire [6:0] debug_1__EVAL_1;
  wire [31:0] debug_1__EVAL_2;
  wire  debug_1__EVAL_3;
  wire [11:0] debug_1__EVAL_4;
  wire  debug_1__EVAL_5;
  wire  debug_1__EVAL_6;
  wire [1:0] debug_1__EVAL_7;
  wire  debug_1__EVAL_8;
  wire  debug_1__EVAL_9;
  wire [3:0] debug_1__EVAL_10;
  wire [31:0] debug_1__EVAL_11;
  wire [2:0] debug_1__EVAL_12;
  wire  debug_1__EVAL_13;
  wire  debug_1__EVAL_14;
  wire [2:0] debug_1__EVAL_15;
  wire [31:0] debug_1__EVAL_16;
  wire [1:0] debug_1__EVAL_17;
  wire  debug_1__EVAL_18;
  wire  debug_1__EVAL_19;
  wire [1:0] debug_1__EVAL_20;
  wire  debug_1__EVAL_21;
  wire  debug_1__EVAL_22;
  wire  debug_1__EVAL_23;
  wire  debug_1__EVAL_24;
  wire [2:0] debug_1__EVAL_25;
  wire [1:0] debug_1__EVAL_26;
  wire  debug_1__EVAL_27;
  wire [31:0] debug_1__EVAL_28;
  wire [2:0] debug_1__EVAL_29;
  wire  debug_1__EVAL_30;
  wire  debug_1__EVAL_31;
  wire  debug_1__EVAL_32;
  wire  _EVAL_4;
  wire [3:0] fbus__EVAL;
  wire  fbus__EVAL_0;
  wire  fbus__EVAL_1;
  wire  fbus__EVAL_2;
  wire [31:0] fbus__EVAL_3;
  wire [31:0] fbus__EVAL_4;
  wire  fbus__EVAL_5;
  wire [1:0] fbus__EVAL_6;
  wire  fbus__EVAL_7;
  wire  fbus__EVAL_8;
  wire [31:0] fbus__EVAL_9;
  wire  fbus__EVAL_10;
  wire  fbus__EVAL_11;
  wire  fbus__EVAL_12;
  wire [2:0] fbus__EVAL_13;
  wire [2:0] fbus__EVAL_14;
  wire [2:0] fbus__EVAL_15;
  wire  fbus__EVAL_16;
  wire  fbus__EVAL_17;
  wire  fbus__EVAL_18;
  wire  fbus__EVAL_19;
  wire [3:0] fbus__EVAL_20;
  wire  fbus__EVAL_21;
  wire  fbus__EVAL_22;
  wire  fbus__EVAL_23;
  wire [1:0] fbus__EVAL_24;
  wire  fbus__EVAL_25;
  wire  fbus__EVAL_26;
  wire [2:0] fbus__EVAL_27;
  wire [31:0] fbus__EVAL_28;
  wire [31:0] fbus__EVAL_29;
  wire [3:0] fbus__EVAL_30;
  wire [3:0] fbus__EVAL_31;
  wire  fbus__EVAL_32;
  wire  fbus__EVAL_33;
  wire  fbus__EVAL_34;
  wire [31:0] fbus__EVAL_35;
  wire [2:0] fbus__EVAL_36;
  wire  fbus__EVAL_37;
  wire  fbus__EVAL_38;
  wire  clic__EVAL;
  wire  clic__EVAL_0;
  wire  clic__EVAL_1;
  wire  clic__EVAL_2;
  wire  clic__EVAL_3;
  wire  clic__EVAL_4;
  wire  clic__EVAL_5;
  wire  clic__EVAL_6;
  wire  clic__EVAL_7;
  wire  clic__EVAL_8;
  wire  clic__EVAL_9;
  wire  clic__EVAL_10;
  wire  clic__EVAL_11;
  wire  clic__EVAL_12;
  wire  clic__EVAL_13;
  wire  clic__EVAL_14;
  wire [7:0] clic__EVAL_15;
  wire  clic__EVAL_16;
  wire  clic__EVAL_17;
  wire  clic__EVAL_18;
  wire  clic__EVAL_19;
  wire  clic__EVAL_20;
  wire  clic__EVAL_21;
  wire  clic__EVAL_22;
  wire  clic__EVAL_23;
  wire  clic__EVAL_24;
  wire [2:0] clic__EVAL_25;
  wire [1:0] clic__EVAL_26;
  wire  clic__EVAL_27;
  wire  clic__EVAL_28;
  wire  clic__EVAL_29;
  wire  clic__EVAL_30;
  wire  clic__EVAL_31;
  wire  clic__EVAL_32;
  wire  clic__EVAL_33;
  wire  clic__EVAL_34;
  wire  clic__EVAL_35;
  wire  clic__EVAL_36;
  wire  clic__EVAL_37;
  wire  clic__EVAL_38;
  wire  clic__EVAL_39;
  wire  clic__EVAL_40;
  wire  clic__EVAL_41;
  wire  clic__EVAL_42;
  wire  clic__EVAL_43;
  wire  clic__EVAL_44;
  wire  clic__EVAL_45;
  wire  clic__EVAL_46;
  wire  clic__EVAL_47;
  wire  clic__EVAL_48;
  wire  clic__EVAL_49;
  wire  clic__EVAL_50;
  wire  clic__EVAL_51;
  wire  clic__EVAL_52;
  wire  clic__EVAL_53;
  wire  clic__EVAL_54;
  wire  clic__EVAL_55;
  wire  clic__EVAL_56;
  wire  clic__EVAL_57;
  wire  clic__EVAL_58;
  wire  clic__EVAL_59;
  wire  clic__EVAL_60;
  wire  clic__EVAL_61;
  wire  clic__EVAL_62;
  wire  clic__EVAL_63;
  wire  clic__EVAL_64;
  wire  clic__EVAL_65;
  wire  clic__EVAL_66;
  wire [31:0] clic__EVAL_67;
  wire [2:0] clic__EVAL_68;
  wire  clic__EVAL_69;
  wire  clic__EVAL_70;
  wire  clic__EVAL_71;
  wire  clic__EVAL_72;
  wire  clic__EVAL_73;
  wire  clic__EVAL_74;
  wire  clic__EVAL_75;
  wire  clic__EVAL_76;
  wire [2:0] clic__EVAL_77;
  wire  clic__EVAL_78;
  wire  clic__EVAL_79;
  wire  clic__EVAL_80;
  wire  clic__EVAL_81;
  wire  clic__EVAL_82;
  wire  clic__EVAL_83;
  wire  clic__EVAL_84;
  wire  clic__EVAL_85;
  wire [7:0] clic__EVAL_86;
  wire  clic__EVAL_87;
  wire [2:0] clic__EVAL_88;
  wire  clic__EVAL_89;
  wire  clic__EVAL_90;
  wire  clic__EVAL_91;
  wire  clic__EVAL_92;
  wire  clic__EVAL_93;
  wire  clic__EVAL_94;
  wire  clic__EVAL_95;
  wire  clic__EVAL_96;
  wire  clic__EVAL_97;
  wire  clic__EVAL_98;
  wire  clic__EVAL_99;
  wire  clic__EVAL_100;
  wire  clic__EVAL_101;
  wire  clic__EVAL_102;
  wire  clic__EVAL_103;
  wire  clic__EVAL_104;
  wire  clic__EVAL_105;
  wire  clic__EVAL_106;
  wire  clic__EVAL_107;
  wire  clic__EVAL_108;
  wire  clic__EVAL_109;
  wire  clic__EVAL_110;
  wire  clic__EVAL_111;
  wire  clic__EVAL_112;
  wire  clic__EVAL_113;
  wire  clic__EVAL_114;
  wire  clic__EVAL_115;
  wire  clic__EVAL_116;
  wire  clic__EVAL_117;
  wire  clic__EVAL_118;
  wire  clic__EVAL_119;
  wire [1:0] clic__EVAL_120;
  wire  clic__EVAL_121;
  wire  clic__EVAL_122;
  wire  clic__EVAL_123;
  wire [3:0] clic__EVAL_124;
  wire  clic__EVAL_125;
  wire  clic__EVAL_126;
  wire  clic__EVAL_127;
  wire  clic__EVAL_128;
  wire  clic__EVAL_129;
  wire  clic__EVAL_130;
  wire [25:0] clic__EVAL_131;
  wire  clic__EVAL_132;
  wire  clic__EVAL_133;
  wire  clic__EVAL_134;
  wire  clic__EVAL_135;
  wire  clic__EVAL_136;
  wire  clic__EVAL_137;
  wire [2:0] clic__EVAL_138;
  wire  clic__EVAL_139;
  wire [31:0] clic__EVAL_140;
  wire  clic__EVAL_141;
  wire  clic__EVAL_142;
  wire  clic__EVAL_143;
  wire  clic__EVAL_144;
  wire  clic__EVAL_145;
  wire  clic__EVAL_146;
  wire  clic__EVAL_147;
  wire  clic__EVAL_148;
  wire  clic__EVAL_149;
  wire  clic__EVAL_150;
  wire  clic__EVAL_151;
  wire  clic__EVAL_152;
  wire  clic__EVAL_153;
  SiFive_TLTestIndicator testIndicator (
    .auto_control_xing_in_a_ready(testIndicator_auto_control_xing_in_a_ready),
    .auto_control_xing_in_a_valid(testIndicator_auto_control_xing_in_a_valid),
    .auto_control_xing_in_a_bits_opcode(testIndicator_auto_control_xing_in_a_bits_opcode),
    .auto_control_xing_in_a_bits_param(testIndicator_auto_control_xing_in_a_bits_param),
    .auto_control_xing_in_a_bits_size(testIndicator_auto_control_xing_in_a_bits_size),
    .auto_control_xing_in_a_bits_source(testIndicator_auto_control_xing_in_a_bits_source),
    .auto_control_xing_in_a_bits_address(testIndicator_auto_control_xing_in_a_bits_address),
    .auto_control_xing_in_a_bits_mask(testIndicator_auto_control_xing_in_a_bits_mask),
    .auto_control_xing_in_a_bits_data(testIndicator_auto_control_xing_in_a_bits_data),
    .auto_control_xing_in_a_bits_corrupt(testIndicator_auto_control_xing_in_a_bits_corrupt),
    .auto_control_xing_in_d_ready(testIndicator_auto_control_xing_in_d_ready),
    .auto_control_xing_in_d_valid(testIndicator_auto_control_xing_in_d_valid),
    .auto_control_xing_in_d_bits_opcode(testIndicator_auto_control_xing_in_d_bits_opcode),
    .auto_control_xing_in_d_bits_size(testIndicator_auto_control_xing_in_d_bits_size),
    .auto_control_xing_in_d_bits_source(testIndicator_auto_control_xing_in_d_bits_source),
    .auto_control_xing_in_d_bits_data(testIndicator_auto_control_xing_in_d_bits_data),
    .clock(testIndicator_clock),
    .reset(testIndicator_reset)
  );
  _EVAL_110 xbar_1 (
    ._EVAL(xbar_1__EVAL),
    ._EVAL_0(xbar_1__EVAL_0)
  );
  _EVAL_110 xbar_2 (
    ._EVAL(xbar_2__EVAL),
    ._EVAL_0(xbar_2__EVAL_0)
  );
  _EVAL_170 island (
    ._EVAL(island__EVAL),
    ._EVAL_0(island__EVAL_0),
    ._EVAL_1(island__EVAL_1),
    ._EVAL_2(island__EVAL_2),
    ._EVAL_3(island__EVAL_3),
    ._EVAL_4(island__EVAL_4),
    ._EVAL_5(island__EVAL_5),
    ._EVAL_6(island__EVAL_6),
    ._EVAL_7(island__EVAL_7),
    ._EVAL_8(island__EVAL_8),
    ._EVAL_9(island__EVAL_9),
    ._EVAL_10(island__EVAL_10),
    ._EVAL_11(island__EVAL_11),
    ._EVAL_12(island__EVAL_12),
    ._EVAL_13(island__EVAL_13),
    ._EVAL_14(island__EVAL_14),
    ._EVAL_15(island__EVAL_15),
    ._EVAL_16(island__EVAL_16)
  );
  _EVAL_37 sbus (
    ._EVAL(sbus__EVAL),
    ._EVAL_0(sbus__EVAL_0),
    ._EVAL_1(sbus__EVAL_1),
    ._EVAL_2(sbus__EVAL_2),
    ._EVAL_3(sbus__EVAL_3),
    ._EVAL_4(sbus__EVAL_4),
    ._EVAL_5(sbus__EVAL_5),
    ._EVAL_6(sbus__EVAL_6),
    ._EVAL_7(sbus__EVAL_7),
    ._EVAL_8(sbus__EVAL_8),
    ._EVAL_9(sbus__EVAL_9),
    ._EVAL_10(sbus__EVAL_10),
    ._EVAL_11(sbus__EVAL_11),
    ._EVAL_12(sbus__EVAL_12),
    ._EVAL_13(sbus__EVAL_13),
    ._EVAL_14(sbus__EVAL_14),
    ._EVAL_15(sbus__EVAL_15),
    ._EVAL_16(sbus__EVAL_16),
    ._EVAL_17(sbus__EVAL_17),
    ._EVAL_18(sbus__EVAL_18),
    ._EVAL_19(sbus__EVAL_19),
    ._EVAL_20(sbus__EVAL_20),
    ._EVAL_21(sbus__EVAL_21),
    ._EVAL_23(sbus__EVAL_23),
    ._EVAL_24(sbus__EVAL_24),
    ._EVAL_25(sbus__EVAL_25),
    ._EVAL_26(sbus__EVAL_26),
    ._EVAL_27(sbus__EVAL_27),
    ._EVAL_28(sbus__EVAL_28),
    ._EVAL_29(sbus__EVAL_29),
    ._EVAL_30(sbus__EVAL_30),
    ._EVAL_31(sbus__EVAL_31),
    ._EVAL_32(sbus__EVAL_32),
    ._EVAL_33(sbus__EVAL_33),
    ._EVAL_34(sbus__EVAL_34),
    ._EVAL_36(sbus__EVAL_36),
    ._EVAL_37(sbus__EVAL_37),
    ._EVAL_38(sbus__EVAL_38),
    ._EVAL_39(sbus__EVAL_39),
    ._EVAL_41(sbus__EVAL_41),
    ._EVAL_42(sbus__EVAL_42),
    ._EVAL_43(sbus__EVAL_43),
    ._EVAL_44(sbus__EVAL_44),
    ._EVAL_45(sbus__EVAL_45),
    ._EVAL_46(sbus__EVAL_46),
    ._EVAL_47(sbus__EVAL_47),
    ._EVAL_48(sbus__EVAL_48),
    ._EVAL_50(sbus__EVAL_50),
    ._EVAL_51(sbus__EVAL_51),
    ._EVAL_52(sbus__EVAL_52),
    ._EVAL_53(sbus__EVAL_53),
    ._EVAL_54(sbus__EVAL_54),
    ._EVAL_55(sbus__EVAL_55),
    ._EVAL_56(sbus__EVAL_56),
    ._EVAL_57(sbus__EVAL_57),
    ._EVAL_58(sbus__EVAL_58),
    ._EVAL_59(sbus__EVAL_59),
    ._EVAL_60(sbus__EVAL_60),
    ._EVAL_61(sbus__EVAL_61),
    ._EVAL_62(sbus__EVAL_62),
    ._EVAL_63(sbus__EVAL_63),
    ._EVAL_64(sbus__EVAL_64),
    ._EVAL_65(sbus__EVAL_65),
    ._EVAL_66(sbus__EVAL_66),
    ._EVAL_67(sbus__EVAL_67),
    ._EVAL_68(sbus__EVAL_68),
    ._EVAL_69(sbus__EVAL_69),
    ._EVAL_70(sbus__EVAL_70),
    ._EVAL_71(sbus__EVAL_71),
    ._EVAL_72(sbus__EVAL_72),
    ._EVAL_73(sbus__EVAL_73),
    ._EVAL_74(sbus__EVAL_74),
    ._EVAL_76(sbus__EVAL_76),
    ._EVAL_77(sbus__EVAL_77),
    ._EVAL_78(sbus__EVAL_78),
    ._EVAL_79(sbus__EVAL_79),
    ._EVAL_80(sbus__EVAL_80),
    ._EVAL_81(sbus__EVAL_81),
    ._EVAL_82(sbus__EVAL_82),
    ._EVAL_83(sbus__EVAL_83),
    ._EVAL_84(sbus__EVAL_84),
    ._EVAL_85(sbus__EVAL_85),
    ._EVAL_86(sbus__EVAL_86),
    ._EVAL_87(sbus__EVAL_87),
    ._EVAL_89(sbus__EVAL_89),
    ._EVAL_90(sbus__EVAL_90),
    ._EVAL_91(sbus__EVAL_91),
    ._EVAL_92(sbus__EVAL_92),
    ._EVAL_93(sbus__EVAL_93),
    ._EVAL_94(sbus__EVAL_94),
    ._EVAL_95(sbus__EVAL_95),
    ._EVAL_96(sbus__EVAL_96),
    ._EVAL_97(sbus__EVAL_97),
    ._EVAL_98(sbus__EVAL_98),
    ._EVAL_99(sbus__EVAL_99),
    ._EVAL_100(sbus__EVAL_100),
    ._EVAL_101(sbus__EVAL_101),
    ._EVAL_102(sbus__EVAL_102),
    ._EVAL_103(sbus__EVAL_103),
    ._EVAL_104(sbus__EVAL_104),
    ._EVAL_105(sbus__EVAL_105),
    ._EVAL_106(sbus__EVAL_106),
    ._EVAL_107(sbus__EVAL_107),
    ._EVAL_108(sbus__EVAL_108),
    ._EVAL_109(sbus__EVAL_109),
    ._EVAL_110(sbus__EVAL_110),
    ._EVAL_111(sbus__EVAL_111),
    ._EVAL_112(sbus__EVAL_112),
    ._EVAL_113(sbus__EVAL_113),
    ._EVAL_114(sbus__EVAL_114),
    ._EVAL_115(sbus__EVAL_115),
    ._EVAL_116(sbus__EVAL_116),
    ._EVAL_117(sbus__EVAL_117),
    ._EVAL_118(sbus__EVAL_118),
    ._EVAL_119(sbus__EVAL_119),
    ._EVAL_120(sbus__EVAL_120),
    ._EVAL_121(sbus__EVAL_121),
    ._EVAL_122(sbus__EVAL_122),
    ._EVAL_123(sbus__EVAL_123),
    ._EVAL_124(sbus__EVAL_124),
    ._EVAL_125(sbus__EVAL_125),
    ._EVAL_126(sbus__EVAL_126),
    ._EVAL_128(sbus__EVAL_128),
    ._EVAL_129(sbus__EVAL_129),
    ._EVAL_130(sbus__EVAL_130),
    ._EVAL_131(sbus__EVAL_131),
    ._EVAL_132(sbus__EVAL_132),
    ._EVAL_133(sbus__EVAL_133),
    ._EVAL_134(sbus__EVAL_134),
    ._EVAL_135(sbus__EVAL_135),
    ._EVAL_136(sbus__EVAL_136),
    ._EVAL_137(sbus__EVAL_137),
    ._EVAL_138(sbus__EVAL_138),
    ._EVAL_139(sbus__EVAL_139),
    ._EVAL_140(sbus__EVAL_140),
    ._EVAL_141(sbus__EVAL_141),
    ._EVAL_142(sbus__EVAL_142),
    ._EVAL_143(sbus__EVAL_143),
    ._EVAL_144(sbus__EVAL_144),
    ._EVAL_146(sbus__EVAL_146),
    ._EVAL_147(sbus__EVAL_147),
    ._EVAL_148(sbus__EVAL_148),
    ._EVAL_150(sbus__EVAL_150),
    ._EVAL_151(sbus__EVAL_151),
    ._EVAL_152(sbus__EVAL_152),
    ._EVAL_153(sbus__EVAL_153),
    ._EVAL_154(sbus__EVAL_154),
    ._EVAL_156(sbus__EVAL_156),
    ._EVAL_157(sbus__EVAL_157),
    ._EVAL_158(sbus__EVAL_158),
    ._EVAL_159(sbus__EVAL_159),
    ._EVAL_160(sbus__EVAL_160),
    ._EVAL_161(sbus__EVAL_161),
    ._EVAL_162(sbus__EVAL_162),
    ._EVAL_164(sbus__EVAL_164),
    ._EVAL_165(sbus__EVAL_165),
    ._EVAL_167(sbus__EVAL_167),
    ._EVAL_168(sbus__EVAL_168),
    ._EVAL_169(sbus__EVAL_169),
    ._EVAL_170(sbus__EVAL_170),
    ._EVAL_171(sbus__EVAL_171)
  );
  _EVAL_190 SynchronizerShiftReg_w1_d3 (
    ._EVAL(SynchronizerShiftReg_w1_d3__EVAL),
    ._EVAL_0(SynchronizerShiftReg_w1_d3__EVAL_0),
    ._EVAL_1(SynchronizerShiftReg_w1_d3__EVAL_1)
  );
  _EVAL_107 cbus (
    ._EVAL(cbus__EVAL),
    ._EVAL_0(cbus__EVAL_0),
    ._EVAL_1(cbus__EVAL_1),
    ._EVAL_2(cbus__EVAL_2),
    ._EVAL_3(cbus__EVAL_3),
    ._EVAL_4(cbus__EVAL_4),
    ._EVAL_7(cbus__EVAL_7),
    ._EVAL_8(cbus__EVAL_8),
    ._EVAL_9(cbus__EVAL_9),
    ._EVAL_10(cbus__EVAL_10),
    ._EVAL_11(cbus__EVAL_11),
    ._EVAL_12(cbus__EVAL_12),
    ._EVAL_13(cbus__EVAL_13),
    ._EVAL_14(cbus__EVAL_14),
    ._EVAL_15(cbus__EVAL_15),
    ._EVAL_16(cbus__EVAL_16),
    ._EVAL_17(cbus__EVAL_17),
    ._EVAL_18(cbus__EVAL_18),
    ._EVAL_19(cbus__EVAL_19),
    ._EVAL_20(cbus__EVAL_20),
    ._EVAL_21(cbus__EVAL_21),
    ._EVAL_22(cbus__EVAL_22),
    ._EVAL_23(cbus__EVAL_23),
    ._EVAL_24(cbus__EVAL_24),
    ._EVAL_25(cbus__EVAL_25),
    ._EVAL_26(cbus__EVAL_26),
    ._EVAL_27(cbus__EVAL_27),
    ._EVAL_28(cbus__EVAL_28),
    ._EVAL_29(cbus__EVAL_29),
    ._EVAL_30(cbus__EVAL_30),
    ._EVAL_31(cbus__EVAL_31),
    ._EVAL_32(cbus__EVAL_32),
    ._EVAL_34(cbus__EVAL_34),
    ._EVAL_35(cbus__EVAL_35),
    ._EVAL_36(cbus__EVAL_36),
    ._EVAL_37(cbus__EVAL_37),
    ._EVAL_38(cbus__EVAL_38),
    ._EVAL_39(cbus__EVAL_39),
    ._EVAL_40(cbus__EVAL_40),
    ._EVAL_41(cbus__EVAL_41),
    ._EVAL_42(cbus__EVAL_42),
    ._EVAL_43(cbus__EVAL_43),
    ._EVAL_44(cbus__EVAL_44),
    ._EVAL_45(cbus__EVAL_45),
    ._EVAL_46(cbus__EVAL_46),
    ._EVAL_47(cbus__EVAL_47),
    ._EVAL_48(cbus__EVAL_48),
    ._EVAL_49(cbus__EVAL_49),
    ._EVAL_50(cbus__EVAL_50),
    ._EVAL_51(cbus__EVAL_51),
    ._EVAL_52(cbus__EVAL_52),
    ._EVAL_54(cbus__EVAL_54),
    ._EVAL_55(cbus__EVAL_55),
    ._EVAL_56(cbus__EVAL_56),
    ._EVAL_57(cbus__EVAL_57),
    ._EVAL_58(cbus__EVAL_58),
    ._EVAL_59(cbus__EVAL_59),
    ._EVAL_60(cbus__EVAL_60),
    ._EVAL_61(cbus__EVAL_61),
    ._EVAL_62(cbus__EVAL_62),
    ._EVAL_63(cbus__EVAL_63),
    ._EVAL_64(cbus__EVAL_64),
    ._EVAL_65(cbus__EVAL_65),
    ._EVAL_66(cbus__EVAL_66),
    ._EVAL_67(cbus__EVAL_67),
    ._EVAL_68(cbus__EVAL_68),
    ._EVAL_69(cbus__EVAL_69),
    ._EVAL_70(cbus__EVAL_70),
    ._EVAL_71(cbus__EVAL_71),
    ._EVAL_72(cbus__EVAL_72),
    ._EVAL_73(cbus__EVAL_73),
    ._EVAL_74(cbus__EVAL_74),
    ._EVAL_75(cbus__EVAL_75),
    ._EVAL_76(cbus__EVAL_76),
    ._EVAL_77(cbus__EVAL_77),
    ._EVAL_78(cbus__EVAL_78),
    ._EVAL_79(cbus__EVAL_79),
    ._EVAL_80(cbus__EVAL_80),
    ._EVAL_81(cbus__EVAL_81),
    ._EVAL_82(cbus__EVAL_82),
    ._EVAL_83(cbus__EVAL_83),
    ._EVAL_84(cbus__EVAL_84),
    ._EVAL_85(cbus__EVAL_85),
    ._EVAL_86(cbus__EVAL_86),
    ._EVAL_87(cbus__EVAL_87),
    ._EVAL_88(cbus__EVAL_88),
    ._EVAL_89(cbus__EVAL_89),
    ._EVAL_90(cbus__EVAL_90)
  );
  _EVAL_165 tile (
    ._EVAL(tile__EVAL),
    ._EVAL_0(tile__EVAL_0),
    ._EVAL_1(tile__EVAL_1),
    ._EVAL_2(tile__EVAL_2),
    ._EVAL_3(tile__EVAL_3),
    ._EVAL_4(tile__EVAL_4),
    ._EVAL_5(tile__EVAL_5),
    ._EVAL_6(tile__EVAL_6),
    ._EVAL_7(tile__EVAL_7),
    ._EVAL_8(tile__EVAL_8),
    ._EVAL_9(tile__EVAL_9),
    ._EVAL_10(tile__EVAL_10),
    ._EVAL_11(tile__EVAL_11),
    ._EVAL_12(tile__EVAL_12),
    ._EVAL_13(tile__EVAL_13),
    ._EVAL_14(tile__EVAL_14),
    ._EVAL_15(tile__EVAL_15),
    ._EVAL_16(tile__EVAL_16),
    ._EVAL_17(tile__EVAL_17),
    ._EVAL_18(tile__EVAL_18),
    ._EVAL_19(tile__EVAL_19),
    ._EVAL_20(tile__EVAL_20),
    ._EVAL_21(tile__EVAL_21),
    ._EVAL_22(tile__EVAL_22),
    ._EVAL_23(tile__EVAL_23),
    ._EVAL_24(tile__EVAL_24),
    ._EVAL_25(tile__EVAL_25),
    ._EVAL_26(tile__EVAL_26),
    ._EVAL_27(tile__EVAL_27),
    ._EVAL_28(tile__EVAL_28),
    ._EVAL_29(tile__EVAL_29),
    ._EVAL_30(tile__EVAL_30),
    ._EVAL_31(tile__EVAL_31),
    ._EVAL_32(tile__EVAL_32),
    ._EVAL_33(tile__EVAL_33),
    ._EVAL_34(tile__EVAL_34),
    ._EVAL_35(tile__EVAL_35),
    ._EVAL_36(tile__EVAL_36),
    ._EVAL_37(tile__EVAL_37),
    ._EVAL_38(tile__EVAL_38),
    ._EVAL_39(tile__EVAL_39),
    ._EVAL_40(tile__EVAL_40),
    ._EVAL_41(tile__EVAL_41),
    ._EVAL_42(tile__EVAL_42),
    ._EVAL_43(tile__EVAL_43),
    ._EVAL_44(tile__EVAL_44),
    ._EVAL_45(tile__EVAL_45),
    ._EVAL_46(tile__EVAL_46),
    ._EVAL_47(tile__EVAL_47),
    ._EVAL_48(tile__EVAL_48),
    ._EVAL_49(tile__EVAL_49),
    ._EVAL_50(tile__EVAL_50),
    ._EVAL_51(tile__EVAL_51),
    ._EVAL_52(tile__EVAL_52),
    ._EVAL_53(tile__EVAL_53),
    ._EVAL_54(tile__EVAL_54),
    ._EVAL_55(tile__EVAL_55),
    ._EVAL_56(tile__EVAL_56),
    ._EVAL_57(tile__EVAL_57),
    ._EVAL_58(tile__EVAL_58),
    ._EVAL_59(tile__EVAL_59),
    ._EVAL_60(tile__EVAL_60),
    ._EVAL_61(tile__EVAL_61),
    ._EVAL_62(tile__EVAL_62),
    ._EVAL_63(tile__EVAL_63),
    ._EVAL_64(tile__EVAL_64),
    ._EVAL_65(tile__EVAL_65),
    ._EVAL_66(tile__EVAL_66),
    ._EVAL_67(tile__EVAL_67)
  );
  _EVAL_108 dummyClockGroupSourceNode (
    ._EVAL(dummyClockGroupSourceNode__EVAL),
    ._EVAL_0(dummyClockGroupSourceNode__EVAL_0),
    ._EVAL_1(dummyClockGroupSourceNode__EVAL_1),
    ._EVAL_2(dummyClockGroupSourceNode__EVAL_2),
    ._EVAL_3(dummyClockGroupSourceNode__EVAL_3),
    ._EVAL_8(dummyClockGroupSourceNode__EVAL_8),
    ._EVAL_11(dummyClockGroupSourceNode__EVAL_11),
    ._EVAL_12(dummyClockGroupSourceNode__EVAL_12)
  );
  _EVAL_175 island_1 (
    ._EVAL(island_1__EVAL),
    ._EVAL_0(island_1__EVAL_0),
    ._EVAL_1(island_1__EVAL_1),
    ._EVAL_2(island_1__EVAL_2),
    ._EVAL_3(island_1__EVAL_3),
    ._EVAL_4(island_1__EVAL_4),
    ._EVAL_5(island_1__EVAL_5),
    ._EVAL_6(island_1__EVAL_6),
    ._EVAL_7(island_1__EVAL_7),
    ._EVAL_8(island_1__EVAL_8),
    ._EVAL_9(island_1__EVAL_9),
    ._EVAL_10(island_1__EVAL_10),
    ._EVAL_11(island_1__EVAL_11),
    ._EVAL_12(island_1__EVAL_12),
    ._EVAL_13(island_1__EVAL_13),
    ._EVAL_14(island_1__EVAL_14),
    ._EVAL_15(island_1__EVAL_15),
    ._EVAL_16(island_1__EVAL_16)
  );
  _EVAL_110 xbar (
    ._EVAL(xbar__EVAL),
    ._EVAL_0(xbar__EVAL_0)
  );
  _EVAL_187 dtm (
    ._EVAL(dtm__EVAL),
    ._EVAL_0(dtm__EVAL_0),
    ._EVAL_1(dtm__EVAL_1),
    ._EVAL_2(dtm__EVAL_2),
    ._EVAL_3(dtm__EVAL_3),
    ._EVAL_4(dtm__EVAL_4),
    ._EVAL_5(dtm__EVAL_5),
    ._EVAL_6(dtm__EVAL_6),
    ._EVAL_7(dtm__EVAL_7),
    ._EVAL_8(dtm__EVAL_8),
    ._EVAL_9(dtm__EVAL_9),
    ._EVAL_10(dtm__EVAL_10),
    ._EVAL_11(dtm__EVAL_11),
    ._EVAL_12(dtm__EVAL_12),
    ._EVAL_13(dtm__EVAL_13),
    ._EVAL_14(dtm__EVAL_14),
    ._EVAL_15(dtm__EVAL_15),
    ._EVAL_16(dtm__EVAL_16)
  );
  _EVAL_149 debug_1 (
    ._EVAL(debug_1__EVAL),
    ._EVAL_0(debug_1__EVAL_0),
    ._EVAL_1(debug_1__EVAL_1),
    ._EVAL_2(debug_1__EVAL_2),
    ._EVAL_3(debug_1__EVAL_3),
    ._EVAL_4(debug_1__EVAL_4),
    ._EVAL_5(debug_1__EVAL_5),
    ._EVAL_6(debug_1__EVAL_6),
    ._EVAL_7(debug_1__EVAL_7),
    ._EVAL_8(debug_1__EVAL_8),
    ._EVAL_9(debug_1__EVAL_9),
    ._EVAL_10(debug_1__EVAL_10),
    ._EVAL_11(debug_1__EVAL_11),
    ._EVAL_12(debug_1__EVAL_12),
    ._EVAL_13(debug_1__EVAL_13),
    ._EVAL_14(debug_1__EVAL_14),
    ._EVAL_15(debug_1__EVAL_15),
    ._EVAL_16(debug_1__EVAL_16),
    ._EVAL_17(debug_1__EVAL_17),
    ._EVAL_18(debug_1__EVAL_18),
    ._EVAL_19(debug_1__EVAL_19),
    ._EVAL_20(debug_1__EVAL_20),
    ._EVAL_21(debug_1__EVAL_21),
    ._EVAL_22(debug_1__EVAL_22),
    ._EVAL_23(debug_1__EVAL_23),
    ._EVAL_24(debug_1__EVAL_24),
    ._EVAL_25(debug_1__EVAL_25),
    ._EVAL_26(debug_1__EVAL_26),
    ._EVAL_27(debug_1__EVAL_27),
    ._EVAL_28(debug_1__EVAL_28),
    ._EVAL_29(debug_1__EVAL_29),
    ._EVAL_30(debug_1__EVAL_30),
    ._EVAL_31(debug_1__EVAL_31),
    ._EVAL_32(debug_1__EVAL_32)
  );
  _EVAL_55 fbus (
    ._EVAL(fbus__EVAL),
    ._EVAL_0(fbus__EVAL_0),
    ._EVAL_1(fbus__EVAL_1),
    ._EVAL_2(fbus__EVAL_2),
    ._EVAL_3(fbus__EVAL_3),
    ._EVAL_4(fbus__EVAL_4),
    ._EVAL_5(fbus__EVAL_5),
    ._EVAL_6(fbus__EVAL_6),
    ._EVAL_7(fbus__EVAL_7),
    ._EVAL_8(fbus__EVAL_8),
    ._EVAL_9(fbus__EVAL_9),
    ._EVAL_10(fbus__EVAL_10),
    ._EVAL_11(fbus__EVAL_11),
    ._EVAL_12(fbus__EVAL_12),
    ._EVAL_13(fbus__EVAL_13),
    ._EVAL_14(fbus__EVAL_14),
    ._EVAL_15(fbus__EVAL_15),
    ._EVAL_16(fbus__EVAL_16),
    ._EVAL_17(fbus__EVAL_17),
    ._EVAL_18(fbus__EVAL_18),
    ._EVAL_19(fbus__EVAL_19),
    ._EVAL_20(fbus__EVAL_20),
    ._EVAL_21(fbus__EVAL_21),
    ._EVAL_22(fbus__EVAL_22),
    ._EVAL_23(fbus__EVAL_23),
    ._EVAL_24(fbus__EVAL_24),
    ._EVAL_25(fbus__EVAL_25),
    ._EVAL_26(fbus__EVAL_26),
    ._EVAL_27(fbus__EVAL_27),
    ._EVAL_28(fbus__EVAL_28),
    ._EVAL_29(fbus__EVAL_29),
    ._EVAL_30(fbus__EVAL_30),
    ._EVAL_31(fbus__EVAL_31),
    ._EVAL_32(fbus__EVAL_32),
    ._EVAL_33(fbus__EVAL_33),
    ._EVAL_34(fbus__EVAL_34),
    ._EVAL_35(fbus__EVAL_35),
    ._EVAL_36(fbus__EVAL_36),
    ._EVAL_37(fbus__EVAL_37),
    ._EVAL_38(fbus__EVAL_38)
  );
  _EVAL_116 clic (
    ._EVAL(clic__EVAL),
    ._EVAL_0(clic__EVAL_0),
    ._EVAL_1(clic__EVAL_1),
    ._EVAL_2(clic__EVAL_2),
    ._EVAL_3(clic__EVAL_3),
    ._EVAL_4(clic__EVAL_4),
    ._EVAL_5(clic__EVAL_5),
    ._EVAL_6(clic__EVAL_6),
    ._EVAL_7(clic__EVAL_7),
    ._EVAL_8(clic__EVAL_8),
    ._EVAL_9(clic__EVAL_9),
    ._EVAL_10(clic__EVAL_10),
    ._EVAL_11(clic__EVAL_11),
    ._EVAL_12(clic__EVAL_12),
    ._EVAL_13(clic__EVAL_13),
    ._EVAL_14(clic__EVAL_14),
    ._EVAL_15(clic__EVAL_15),
    ._EVAL_16(clic__EVAL_16),
    ._EVAL_17(clic__EVAL_17),
    ._EVAL_18(clic__EVAL_18),
    ._EVAL_19(clic__EVAL_19),
    ._EVAL_20(clic__EVAL_20),
    ._EVAL_21(clic__EVAL_21),
    ._EVAL_22(clic__EVAL_22),
    ._EVAL_23(clic__EVAL_23),
    ._EVAL_24(clic__EVAL_24),
    ._EVAL_25(clic__EVAL_25),
    ._EVAL_26(clic__EVAL_26),
    ._EVAL_27(clic__EVAL_27),
    ._EVAL_28(clic__EVAL_28),
    ._EVAL_29(clic__EVAL_29),
    ._EVAL_30(clic__EVAL_30),
    ._EVAL_31(clic__EVAL_31),
    ._EVAL_32(clic__EVAL_32),
    ._EVAL_33(clic__EVAL_33),
    ._EVAL_34(clic__EVAL_34),
    ._EVAL_35(clic__EVAL_35),
    ._EVAL_36(clic__EVAL_36),
    ._EVAL_37(clic__EVAL_37),
    ._EVAL_38(clic__EVAL_38),
    ._EVAL_39(clic__EVAL_39),
    ._EVAL_40(clic__EVAL_40),
    ._EVAL_41(clic__EVAL_41),
    ._EVAL_42(clic__EVAL_42),
    ._EVAL_43(clic__EVAL_43),
    ._EVAL_44(clic__EVAL_44),
    ._EVAL_45(clic__EVAL_45),
    ._EVAL_46(clic__EVAL_46),
    ._EVAL_47(clic__EVAL_47),
    ._EVAL_48(clic__EVAL_48),
    ._EVAL_49(clic__EVAL_49),
    ._EVAL_50(clic__EVAL_50),
    ._EVAL_51(clic__EVAL_51),
    ._EVAL_52(clic__EVAL_52),
    ._EVAL_53(clic__EVAL_53),
    ._EVAL_54(clic__EVAL_54),
    ._EVAL_55(clic__EVAL_55),
    ._EVAL_56(clic__EVAL_56),
    ._EVAL_57(clic__EVAL_57),
    ._EVAL_58(clic__EVAL_58),
    ._EVAL_59(clic__EVAL_59),
    ._EVAL_60(clic__EVAL_60),
    ._EVAL_61(clic__EVAL_61),
    ._EVAL_62(clic__EVAL_62),
    ._EVAL_63(clic__EVAL_63),
    ._EVAL_64(clic__EVAL_64),
    ._EVAL_65(clic__EVAL_65),
    ._EVAL_66(clic__EVAL_66),
    ._EVAL_67(clic__EVAL_67),
    ._EVAL_68(clic__EVAL_68),
    ._EVAL_69(clic__EVAL_69),
    ._EVAL_70(clic__EVAL_70),
    ._EVAL_71(clic__EVAL_71),
    ._EVAL_72(clic__EVAL_72),
    ._EVAL_73(clic__EVAL_73),
    ._EVAL_74(clic__EVAL_74),
    ._EVAL_75(clic__EVAL_75),
    ._EVAL_76(clic__EVAL_76),
    ._EVAL_77(clic__EVAL_77),
    ._EVAL_78(clic__EVAL_78),
    ._EVAL_79(clic__EVAL_79),
    ._EVAL_80(clic__EVAL_80),
    ._EVAL_81(clic__EVAL_81),
    ._EVAL_82(clic__EVAL_82),
    ._EVAL_83(clic__EVAL_83),
    ._EVAL_84(clic__EVAL_84),
    ._EVAL_85(clic__EVAL_85),
    ._EVAL_86(clic__EVAL_86),
    ._EVAL_87(clic__EVAL_87),
    ._EVAL_88(clic__EVAL_88),
    ._EVAL_89(clic__EVAL_89),
    ._EVAL_90(clic__EVAL_90),
    ._EVAL_91(clic__EVAL_91),
    ._EVAL_92(clic__EVAL_92),
    ._EVAL_93(clic__EVAL_93),
    ._EVAL_94(clic__EVAL_94),
    ._EVAL_95(clic__EVAL_95),
    ._EVAL_96(clic__EVAL_96),
    ._EVAL_97(clic__EVAL_97),
    ._EVAL_98(clic__EVAL_98),
    ._EVAL_99(clic__EVAL_99),
    ._EVAL_100(clic__EVAL_100),
    ._EVAL_101(clic__EVAL_101),
    ._EVAL_102(clic__EVAL_102),
    ._EVAL_103(clic__EVAL_103),
    ._EVAL_104(clic__EVAL_104),
    ._EVAL_105(clic__EVAL_105),
    ._EVAL_106(clic__EVAL_106),
    ._EVAL_107(clic__EVAL_107),
    ._EVAL_108(clic__EVAL_108),
    ._EVAL_109(clic__EVAL_109),
    ._EVAL_110(clic__EVAL_110),
    ._EVAL_111(clic__EVAL_111),
    ._EVAL_112(clic__EVAL_112),
    ._EVAL_113(clic__EVAL_113),
    ._EVAL_114(clic__EVAL_114),
    ._EVAL_115(clic__EVAL_115),
    ._EVAL_116(clic__EVAL_116),
    ._EVAL_117(clic__EVAL_117),
    ._EVAL_118(clic__EVAL_118),
    ._EVAL_119(clic__EVAL_119),
    ._EVAL_120(clic__EVAL_120),
    ._EVAL_121(clic__EVAL_121),
    ._EVAL_122(clic__EVAL_122),
    ._EVAL_123(clic__EVAL_123),
    ._EVAL_124(clic__EVAL_124),
    ._EVAL_125(clic__EVAL_125),
    ._EVAL_126(clic__EVAL_126),
    ._EVAL_127(clic__EVAL_127),
    ._EVAL_128(clic__EVAL_128),
    ._EVAL_129(clic__EVAL_129),
    ._EVAL_130(clic__EVAL_130),
    ._EVAL_131(clic__EVAL_131),
    ._EVAL_132(clic__EVAL_132),
    ._EVAL_133(clic__EVAL_133),
    ._EVAL_134(clic__EVAL_134),
    ._EVAL_135(clic__EVAL_135),
    ._EVAL_136(clic__EVAL_136),
    ._EVAL_137(clic__EVAL_137),
    ._EVAL_138(clic__EVAL_138),
    ._EVAL_139(clic__EVAL_139),
    ._EVAL_140(clic__EVAL_140),
    ._EVAL_141(clic__EVAL_141),
    ._EVAL_142(clic__EVAL_142),
    ._EVAL_143(clic__EVAL_143),
    ._EVAL_144(clic__EVAL_144),
    ._EVAL_145(clic__EVAL_145),
    ._EVAL_146(clic__EVAL_146),
    ._EVAL_147(clic__EVAL_147),
    ._EVAL_148(clic__EVAL_148),
    ._EVAL_149(clic__EVAL_149),
    ._EVAL_150(clic__EVAL_150),
    ._EVAL_151(clic__EVAL_151),
    ._EVAL_152(clic__EVAL_152),
    ._EVAL_153(clic__EVAL_153)
  );
  assign debug_1__EVAL_8 = dtm__EVAL_14;
  assign cbus__EVAL_61 = sbus__EVAL_164;
  assign clic__EVAL_46 = local_interrupts_0[9];
  assign clic__EVAL_118 = local_interrupts_0[81];
  assign debug_1__EVAL_22 = debug_systemjtag_reset;
  assign clic__EVAL_97 = local_interrupts_0[120];
  assign sys_port_ahb_0_hprot = sbus__EVAL_124;
  assign clic__EVAL_91 = local_interrupts_0[54];
  assign sbus__EVAL_169 = tile__EVAL_50;
  assign fbus__EVAL_30 = front_port_ahb_0_hprot;
  assign sbus__EVAL_170 = tile__EVAL_23;
  assign cbus__EVAL_9 = testIndicator_auto_control_xing_in_d_bits_size;
  assign clic__EVAL_151 = local_interrupts_0[117];
  assign tile__EVAL_1 = sbus__EVAL_167;
  assign island_1__EVAL_7 = sbus__EVAL_165;
  assign sbus__EVAL_98 = tile__EVAL_60;
  assign sbus__EVAL_36 = cbus__EVAL_60;
  assign tile__EVAL_54 = sbus__EVAL_54;
  assign debug_1__EVAL_25 = cbus__EVAL_87;
  assign sbus__EVAL_139 = tile__EVAL_48;
  assign clic__EVAL_23 = local_interrupts_0[87];
  assign sbus__EVAL_115 = fbus__EVAL_4;
  assign clic__EVAL = local_interrupts_0[77];
  assign fbus__EVAL_28 = front_port_ahb_0_hwdata;
  assign sbus__EVAL_134 = tile__EVAL_16;
  assign debug_1__EVAL_19 = cbus__EVAL_18;
  assign clic__EVAL_135 = local_interrupts_0[14];
  assign clic__EVAL_140 = cbus__EVAL_32;
  assign clic__EVAL_95 = local_interrupts_0[40];
  assign testIndicator_auto_control_xing_in_a_bits_size = cbus__EVAL_26;
  assign testIndicator_auto_control_xing_in_a_bits_opcode = cbus__EVAL_2;
  assign tile__EVAL_39 = sbus__EVAL_26;
  assign clic__EVAL_58 = local_interrupts_0[90];
  assign fbus__EVAL_11 = sbus__EVAL_131;
  assign clic__EVAL_115 = local_interrupts_0[85];
  assign sbus__EVAL_85 = fbus__EVAL_19;
  assign dtm__EVAL_6 = debug_systemjtag_part_number;
  assign sbus__EVAL_113 = tile__EVAL_13;
  assign sbus__EVAL_77 = tile__EVAL_25;
  assign tile__EVAL_53 = sbus__EVAL;
  assign debug_1__EVAL_18 = cbus__EVAL_73;
  assign clic__EVAL_39 = local_interrupts_0[25];
  assign sbus__EVAL_10 = island__EVAL_0;
  assign tile__EVAL_18 = sbus__EVAL_7;
  assign sbus__EVAL_102 = tile__EVAL_22;
  assign clic__EVAL_103 = local_interrupts_0[43];
  assign sbus__EVAL_9 = fbus__EVAL_16;
  assign _EVAL_4 = _EVAL & _EVAL_1;
  assign clic__EVAL_146 = local_interrupts_0[22];
  assign clic__EVAL_100 = local_interrupts_0[104];
  assign clic__EVAL_70 = local_interrupts_0[23];
  assign clic__EVAL_16 = local_interrupts_0[53];
  assign island_1__EVAL = sbus__EVAL_150;
  assign clic__EVAL_9 = local_interrupts_0[94];
  assign sbus__EVAL_93 = tile__EVAL_41;
  assign clic__EVAL_6 = local_interrupts_0[84];
  assign sbus__EVAL_101 = fbus__EVAL_8;
  assign cbus__EVAL_88 = periph_port_ahb_0_hready;
  assign debug_1__EVAL_17 = dtm__EVAL_15;
  assign fbus__EVAL_6 = front_port_ahb_0_htrans;
  assign clic__EVAL_74 = local_interrupts_0[70];
  assign clic__EVAL_119 = local_interrupts_0[47];
  assign clic__EVAL_75 = local_interrupts_0[35];
  assign sbus__EVAL_63 = dummyClockGroupSourceNode__EVAL_11;
  assign sbus__EVAL_73 = cbus__EVAL_55;
  assign fbus__EVAL_36 = front_port_ahb_0_hsize;
  assign clic__EVAL_88 = cbus__EVAL_46;
  assign cbus__EVAL_17 = clic__EVAL_120;
  assign clic__EVAL_104 = local_interrupts_0[102];
  assign sbus__EVAL_143 = tile__EVAL_46;
  assign tile__EVAL_35 = clic__EVAL_145;
  assign periph_port_ahb_0_hwrite = cbus__EVAL_77;
  assign sbus__EVAL_11 = fbus__EVAL_31;
  assign testIndicator_auto_control_xing_in_a_bits_source = cbus__EVAL_21;
  assign clic__EVAL_132 = local_interrupts_0[93];
  assign sbus__EVAL_68 = cbus__EVAL_56;
  assign cbus__EVAL_34 = debug_1__EVAL_26;
  assign clic__EVAL_28 = local_interrupts_0[39];
  assign cbus__EVAL_50 = sbus__EVAL_52;
  assign periph_port_ahb_0_hburst = 3'h0;
  assign cbus__EVAL_49 = sbus__EVAL_80;
  assign sbus__EVAL_64 = fbus__EVAL_15;
  assign clic__EVAL_148 = local_interrupts_0[65];
  assign clic__EVAL_110 = local_interrupts_0[69];
  assign debug_1__EVAL_1 = dtm__EVAL_1;
  assign clic__EVAL_19 = local_interrupts_0[67];
  assign sbus__EVAL_6 = tile__EVAL_62;
  assign dtm__EVAL_11 = debug_1__EVAL_20;
  assign fbus__EVAL_38 = front_port_ahb_0_hready;
  assign clic__EVAL_12 = local_interrupts_0[106];
  assign island__EVAL_11 = sbus__EVAL_154;
  assign clic__EVAL_30 = local_interrupts_0[103];
  assign periph_port_ahb_0_haddr = cbus__EVAL_13;
  assign clic__EVAL_102 = local_interrupts_0[60];
  assign clic__EVAL_64 = local_interrupts_0[17];
  assign clic__EVAL_62 = local_interrupts_0[107];
  assign clic__EVAL_99 = local_interrupts_0[19];
  assign fbus__EVAL_27 = sbus__EVAL_58;
  assign clic__EVAL_83 = local_interrupts_0[26];
  assign clic__EVAL_65 = local_interrupts_0[2];
  assign clic__EVAL_5 = local_interrupts_0[55];
  assign clic__EVAL_127 = local_interrupts_0[79];
  assign cbus__EVAL_74 = testIndicator_auto_control_xing_in_d_bits_source;
  assign debug_1__EVAL_4 = cbus__EVAL_22;
  assign testIndicator_clock = cbus__EVAL_78;
  assign fbus__EVAL_17 = sbus__EVAL_140;
  assign clic__EVAL_133 = local_interrupts_0[0];
  assign clic__EVAL_82 = local_interrupts_0[86];
  assign clic__EVAL_122 = local_interrupts_0[113];
  assign tile__EVAL_66 = reset_vector_0;
  assign clic__EVAL_84 = local_interrupts_0[4];
  assign debug_1__EVAL_32 = debug_dmactiveAck;
  assign clic__EVAL_44 = local_interrupts_0[13];
  assign cbus__EVAL_69 = sbus__EVAL_168;
  assign sbus__EVAL_39 = cbus__EVAL_11;
  assign island__EVAL_16 = sbus__EVAL_118;
  assign sbus__EVAL_111 = tile__EVAL_8;
  assign testIndicator_auto_control_xing_in_d_ready = cbus__EVAL_39;
  assign clic__EVAL_129 = local_interrupts_0[110];
  assign debug_1__EVAL_30 = debug_reset;
  assign fbus__EVAL_1 = front_port_ahb_0_hwrite;
  assign tile__EVAL_43 = sbus__EVAL_15;
  assign sbus__EVAL_106 = tile__EVAL_26;
  assign cbus__EVAL_19 = debug_1__EVAL_15;
  assign fbus__EVAL_7 = sbus__EVAL_122;
  assign fbus__EVAL_23 = front_port_ahb_0_hsel;
  assign sys_port_ahb_0_hburst = sbus__EVAL_66;
  assign dtm__EVAL_16 = debug_systemjtag_jtag_TMS;
  assign clic__EVAL_53 = local_interrupts_0[124];
  assign clic__EVAL_48 = local_interrupts_0[108];
  assign fbus__EVAL_21 = sbus__EVAL_24;
  assign sbus__EVAL_126 = island_1__EVAL_15;
  assign sbus__EVAL_8 = fbus__EVAL_32;
  assign clic__EVAL_137 = local_interrupts_0[27];
  assign sbus__EVAL_137 = fbus__EVAL_5;
  assign tile__EVAL_15 = sbus__EVAL_136;
  assign clic__EVAL_114 = local_interrupts_0[12];
  assign clic__EVAL_108 = local_interrupts_0[59];
  assign sbus__EVAL_125 = tile__EVAL_34;
  assign cbus__EVAL = debug_1__EVAL_11;
  assign clic__EVAL_101 = _EVAL_0;
  assign cbus__EVAL_84 = periph_port_ahb_0_hresp;
  assign cbus__EVAL_80 = sbus__EVAL_130;
  assign testIndicator_auto_control_xing_in_a_bits_data = cbus__EVAL_8;
  assign clic__EVAL_96 = local_interrupts_0[96];
  assign clic__EVAL_121 = local_interrupts_0[92];
  assign debug_systemjtag_jtag_TDO_driven = dtm__EVAL_10;
  assign tile__EVAL_14 = clic__EVAL_86;
  assign sbus__EVAL_55 = dummyClockGroupSourceNode__EVAL;
  assign island_1__EVAL_14 = sbus__EVAL_157;
  assign clic__EVAL_144 = local_interrupts_0[64];
  assign clic__EVAL_123 = local_interrupts_0[21];
  assign clic__EVAL_71 = local_interrupts_0[8];
  assign debug_1__EVAL_13 = dtm__EVAL;
  assign debug_systemjtag_jtag_TDO_data = dtm__EVAL_4;
  assign sys_port_ahb_0_haddr = sbus__EVAL_1;
  assign island_1__EVAL_9 = sbus__EVAL_12;
  assign sbus__EVAL_112 = fbus__EVAL_13;
  assign island_1__EVAL_13 = sbus__EVAL_119;
  assign island__EVAL_15 = sbus__EVAL_70;
  assign clic__EVAL_153 = local_interrupts_0[115];
  assign clic__EVAL_13 = local_interrupts_0[116];
  assign periph_port_ahb_0_hsize = cbus__EVAL_72;
  assign cbus__EVAL_41 = testIndicator_auto_control_xing_in_d_bits_data;
  assign clic__EVAL_1 = local_interrupts_0[100];
  assign sbus__EVAL_33 = island__EVAL_9;
  assign clic__EVAL_21 = local_interrupts_0[88];
  assign clic__EVAL_76 = local_interrupts_0[66];
  assign clic__EVAL_85 = local_interrupts_0[91];
  assign clic__EVAL_54 = local_interrupts_0[58];
  assign cbus__EVAL_16 = sbus__EVAL_156;
  assign clic__EVAL_43 = local_interrupts_0[126];
  assign clic__EVAL_32 = local_interrupts_0[118];
  assign periph_port_ahb_0_hprot = cbus__EVAL_79;
  assign island__EVAL_8 = sbus__EVAL_89;
  assign island__EVAL_2 = sbus__EVAL_60;
  assign cbus__EVAL_10 = periph_port_ahb_0_hrdata;
  assign sbus__EVAL_141 = island_1__EVAL_16;
  assign clic__EVAL_111 = local_interrupts_0[32];
  assign clic__EVAL_14 = local_interrupts_0[62];
  assign debug_1__EVAL_7 = cbus__EVAL_30;
  assign clic__EVAL_50 = local_interrupts_0[71];
  assign clic__EVAL_41 = local_interrupts_0[95];
  assign clic__EVAL_112 = cbus__EVAL_86;
  assign sys_port_ahb_0_htrans = sbus__EVAL_162;
  assign dtm__EVAL_7 = debug_1__EVAL_27;
  assign island__EVAL_14 = sbus__EVAL_147;
  assign sbus__EVAL_38 = tile__EVAL_47;
  assign dummyClockGroupSourceNode__EVAL_2 = clock;
  assign clic__EVAL_25 = cbus__EVAL_76;
  assign testIndicator_auto_control_xing_in_a_bits_corrupt = cbus__EVAL_31;
  assign clic__EVAL_116 = local_interrupts_0[101];
  assign tile__EVAL_4 = clic__EVAL_15;
  assign front_port_ahb_0_hreadyout = fbus__EVAL_33;
  assign dtm__EVAL_0 = debug_systemjtag_reset;
  assign tile__EVAL_10 = psd_test_clock_enable;
  assign tile__EVAL_51 = clic__EVAL_49;
  assign sbus__EVAL_65 = tile__EVAL_12;
  assign clic__EVAL_61 = local_interrupts_0[10];
  assign tile__EVAL_58 = sbus__EVAL_67;
  assign debug_1__EVAL_12 = cbus__EVAL_82;
  assign tile__EVAL_63 = _EVAL_3[0];
  assign sbus__EVAL_31 = fbus__EVAL_2;
  assign clic__EVAL_36 = local_interrupts_0[75];
  assign debug_1__EVAL_10 = cbus__EVAL_51;
  assign tile__EVAL_27 = sbus__EVAL_100;
  assign halt_from_tile_0 = xbar__EVAL;
  assign sbus__EVAL_74 = island__EVAL_7;
  assign dtm__EVAL_12 = debug_1__EVAL_16;
  assign xbar_2__EVAL_0 = tile__EVAL_55;
  assign cbus__EVAL_35 = sbus__EVAL_19;
  assign sbus__EVAL_158 = dummyClockGroupSourceNode__EVAL_1;
  assign fbus__EVAL = sbus__EVAL_132;
  assign clic__EVAL_152 = local_interrupts_0[42];
  assign sbus__EVAL_146 = cbus__EVAL_29;
  assign sbus__EVAL_121 = tile__EVAL_2;
  assign tile__EVAL_28 = sbus__EVAL_37;
  assign clic__EVAL_56 = local_interrupts_0[44];
  assign SynchronizerShiftReg_w1_d3__EVAL_0 = clock;
  assign sbus__EVAL_103 = tile__EVAL_57;
  assign dtm__EVAL_2 = debug_systemjtag_jtag_TCK;
  assign island__EVAL_4 = sbus__EVAL_144;
  assign clic__EVAL_69 = local_interrupts_0[51];
  assign fbus__EVAL_25 = sbus__EVAL_28;
  assign sbus__EVAL_25 = island_1__EVAL_1;
  assign clic__EVAL_45 = local_interrupts_0[114];
  assign sbus__EVAL_48 = tile__EVAL_40;
  assign SynchronizerShiftReg_w1_d3__EVAL_1 = rtc_toggle;
  assign clic__EVAL_35 = local_interrupts_0[68];
  assign island__EVAL = sbus__EVAL_29;
  assign debug_1__EVAL_0 = debug_clock;
  assign debug_1__EVAL_28 = dtm__EVAL_3;
  assign tile__EVAL_37 = sbus__EVAL_69;
  assign cbus__EVAL_0 = sbus__EVAL_81;
  assign clic__EVAL_147 = local_interrupts_0[122];
  assign clic__EVAL_2 = local_interrupts_0[76];
  assign front_port_ahb_0_hrdata = fbus__EVAL_9;
  assign clic__EVAL_134 = local_interrupts_0[112];
  assign sbus__EVAL_91 = fbus__EVAL_12;
  assign sbus__EVAL_51 = sys_port_ahb_0_hresp;
  assign sbus__EVAL_114 = tile__EVAL_19;
  assign tile__EVAL_56 = sbus__EVAL_18;
  assign sbus__EVAL_129 = fbus__EVAL_37;
  assign clic__EVAL_93 = local_interrupts_0[98];
  assign clic__EVAL_0 = local_interrupts_0[52];
  assign clic__EVAL_20 = local_interrupts_0[38];
  assign testIndicator_reset = cbus__EVAL_70;
  assign clic__EVAL_59 = local_interrupts_0[119];
  assign cease_from_tile_0 = xbar_2__EVAL;
  assign clic__EVAL_130 = local_interrupts_0[36];
  assign clic__EVAL_139 = local_interrupts_0[28];
  assign clic__EVAL_81 = local_interrupts_0[46];
  assign clic__EVAL_73 = local_interrupts_0[89];
  assign island_1__EVAL_0 = sbus__EVAL_30;
  assign clic__EVAL_31 = local_interrupts_0[5];
  assign clic__EVAL_11 = cbus__EVAL_90;
  assign clic__EVAL_26 = cbus__EVAL_68;
  assign clic__EVAL_106 = clock;
  assign sbus__EVAL_87 = tile__EVAL_5;
  assign fbus__EVAL_29 = sbus__EVAL_2;
  assign clic__EVAL_117 = local_interrupts_0[45];
  assign clic__EVAL_94 = local_interrupts_0[78];
  assign sbus__EVAL_95 = fbus__EVAL_10;
  assign cbus__EVAL_89 = clic__EVAL_138;
  assign tile__EVAL_29 = sbus__EVAL_14;
  assign island__EVAL_12 = sbus__EVAL_17;
  assign clic__EVAL_7 = local_interrupts_0[123];
  assign periph_port_ahb_0_hmastlock = 1'h0;
  assign tile__EVAL_3 = clic__EVAL_47;
  assign sbus__EVAL_71 = tile__EVAL_31;
  assign fbus__EVAL_35 = front_port_ahb_0_haddr;
  assign cbus__EVAL_48 = clic__EVAL_68;
  assign tile__EVAL_9 = sbus__EVAL_138;
  assign clic__EVAL_143 = local_interrupts_0[37];
  assign clic__EVAL_87 = local_interrupts_0[20];
  assign tile__EVAL = clic__EVAL_78;
  assign sbus__EVAL_97 = sys_port_ahb_0_hready;
  assign tile__EVAL_17 = sbus__EVAL_47;
  assign clic__EVAL_17 = local_interrupts_0[56];
  assign sbus__EVAL_171 = tile__EVAL_65;
  assign sbus__EVAL_56 = island__EVAL_1;
  assign sbus__EVAL_108 = island_1__EVAL_2;
  assign sbus__EVAL_94 = island__EVAL_13;
  assign clic__EVAL_92 = local_interrupts_0[111];
  assign clic__EVAL_22 = local_interrupts_0[61];
  assign debug_ndreset = debug_1__EVAL_21;
  assign sbus__EVAL_109 = island_1__EVAL_10;
  assign clic__EVAL_90 = local_interrupts_0[41];
  assign tile__EVAL_61 = sbus__EVAL_86;
  assign sbus__EVAL_107 = tile__EVAL_64;
  assign clic__EVAL_33 = local_interrupts_0[7];
  assign debug_dmactive = debug_1__EVAL_23;
  assign clic__EVAL_141 = local_interrupts_0[15];
  assign dummyClockGroupSourceNode__EVAL_12 = reset;
  assign sbus__EVAL_78 = cbus__EVAL_52;
  assign sbus__EVAL_4 = tile__EVAL_45;
  assign clic__EVAL_80 = local_interrupts_0[121];
  assign clic__EVAL_34 = cbus__EVAL_36;
  assign sbus__EVAL_0 = fbus__EVAL_18;
  assign clic__EVAL_29 = local_interrupts_0[30];
  assign clic__EVAL_8 = local_interrupts_0[97];
  assign front_port_ahb_0_hresp = fbus__EVAL_22;
  assign sbus__EVAL_32 = cbus__EVAL_45;
  assign tile__EVAL_44 = sbus__EVAL_5;
  assign island_1__EVAL_11 = sbus__EVAL_27;
  assign clic__EVAL_126 = local_interrupts_0[105];
  assign cbus__EVAL_7 = clic__EVAL_67;
  assign xbar_1__EVAL_0 = tile__EVAL_33;
  assign clic__EVAL_40 = local_interrupts_0[11];
  assign cbus__EVAL_15 = testIndicator_auto_control_xing_in_d_bits_opcode;
  assign clic__EVAL_52 = local_interrupts_0[34];
  assign sys_port_ahb_0_hwrite = sbus__EVAL_76;
  assign clic__EVAL_42 = local_interrupts_0[99];
  assign tile__EVAL_52 = clic__EVAL_113;
  assign fbus__EVAL_24 = sbus__EVAL_128;
  assign cbus__EVAL_12 = sbus__EVAL_83;
  assign dtm__EVAL_13 = debug_systemjtag_mfr_id;
  assign testIndicator_auto_control_xing_in_a_bits_mask = cbus__EVAL_20;
  assign clic__EVAL_63 = local_interrupts_0[49];
  assign xbar__EVAL_0 = tile__EVAL_7;
  assign sbus__EVAL_44 = cbus__EVAL_37;
  assign periph_port_ahb_0_hwdata = cbus__EVAL_25;
  assign dtm__EVAL_9 = debug_1__EVAL_3;
  assign sys_port_ahb_0_hwdata = sbus__EVAL_79;
  assign clic__EVAL_98 = local_interrupts_0[1];
  assign tile__EVAL_59 = sbus__EVAL_148;
  assign debug_1__EVAL_5 = cbus__EVAL_28;
  assign cbus__EVAL_14 = sbus__EVAL_21;
  assign sys_port_ahb_0_hmastlock = 1'h0;
  assign island_1__EVAL_8 = sbus__EVAL_116;
  assign sbus__EVAL_53 = tile__EVAL_11;
  assign tile__EVAL_32 = reset;
  assign clic__EVAL_128 = local_interrupts_0[3];
  assign island_1__EVAL_12 = sbus__EVAL_13;
  assign cbus__EVAL_42 = clic__EVAL_18;
  assign tile__EVAL_6 = sbus__EVAL_61;
  assign clic__EVAL_38 = local_interrupts_0[109];
  assign cbus__EVAL_75 = debug_1__EVAL_24;
  assign sbus__EVAL_110 = island__EVAL_3;
  assign testIndicator_auto_control_xing_in_a_bits_param = cbus__EVAL_81;
  assign sbus__EVAL_104 = tile__EVAL_20;
  assign sbus__EVAL_41 = cbus__EVAL_27;
  assign clic__EVAL_51 = local_interrupts_0[16];
  assign clic__EVAL_105 = local_interrupts_0[18];
  assign sbus__EVAL_153 = dummyClockGroupSourceNode__EVAL_8;
  assign tile__EVAL_21 = clock;
  assign periph_port_ahb_0_htrans = cbus__EVAL_85;
  assign island__EVAL_6 = sbus__EVAL_34;
  assign sbus__EVAL_43 = tile__EVAL_0;
  assign sbus__EVAL_152 = tile__EVAL_49;
  assign sbus__EVAL_45 = island_1__EVAL_5;
  assign wfi_from_tile_0 = xbar_1__EVAL;
  assign clic__EVAL_27 = local_interrupts_0[83];
  assign cbus__EVAL_4 = sbus__EVAL_20;
  assign fbus__EVAL_26 = sbus__EVAL_120;
  assign cbus__EVAL_38 = clic__EVAL_142;
  assign _EVAL_1 = ~_EVAL_2;
  assign sbus__EVAL_161 = sys_port_ahb_0_hrdata;
  assign cbus__EVAL_67 = sbus__EVAL_16;
  assign clic__EVAL_37 = local_interrupts_0[31];
  assign cbus__EVAL_83 = testIndicator_auto_control_xing_in_a_ready;
  assign sbus__EVAL_82 = tile__EVAL_38;
  assign clic__EVAL_66 = local_interrupts_0[57];
  assign island__EVAL_5 = sbus__EVAL_57;
  assign sbus__EVAL_117 = tile__EVAL_42;
  assign cbus__EVAL_23 = sbus__EVAL_135;
  assign clic__EVAL_79 = local_interrupts_0[33];
  assign sbus__EVAL_42 = fbus__EVAL_3;
  assign clic__EVAL_55 = local_interrupts_0[80];
  assign _EVAL_3 = 2'h0;
  assign _EVAL = SynchronizerShiftReg_w1_d3__EVAL;
  assign cbus__EVAL_43 = sbus__EVAL_62;
  assign sys_port_ahb_0_hsize = sbus__EVAL_123;
  assign testIndicator_auto_control_xing_in_a_bits_address = cbus__EVAL_64;
  assign cbus__EVAL_40 = sbus__EVAL_160;
  assign clic__EVAL_150 = local_interrupts_0[29];
  assign testIndicator_auto_control_xing_in_a_valid = cbus__EVAL_71;
  assign cbus__EVAL_62 = sbus__EVAL_3;
  assign sbus__EVAL_159 = fbus__EVAL_0;
  assign clic__EVAL_60 = debug_1__EVAL_14;
  assign cbus__EVAL_57 = testIndicator_auto_control_xing_in_d_valid;
  assign clic__EVAL_57 = local_interrupts_0[24];
  assign dtm__EVAL_8 = debug_systemjtag_jtag_TDI;
  assign island__EVAL_10 = sbus__EVAL_90;
  assign clic__EVAL_10 = local_interrupts_0[72];
  assign debug_1__EVAL_2 = cbus__EVAL_58;
  assign island_1__EVAL_3 = sbus__EVAL_34;
  assign clic__EVAL_125 = local_interrupts_0[82];
  assign tile__EVAL_36 = sbus__EVAL_96;
  assign clic__EVAL_124 = cbus__EVAL_1;
  assign dtm__EVAL_5 = debug_systemjtag_version;
  assign cbus__EVAL_63 = sbus__EVAL_142;
  assign fbus__EVAL_14 = front_port_ahb_0_hburst;
  assign cbus__EVAL_59 = sbus__EVAL_105;
  assign island_1__EVAL_4 = sbus__EVAL_17;
  assign debug_1__EVAL_6 = resetctrl_hartIsInReset_0;
  assign debug_1__EVAL_31 = debug_systemjtag_jtag_TCK;
  assign clic__EVAL_24 = reset;
  assign fbus__EVAL_34 = sbus__EVAL_50;
  assign clic__EVAL_72 = local_interrupts_0[48];
  assign clic__EVAL_3 = local_interrupts_0[50];
  assign debug_1__EVAL_29 = cbus__EVAL_47;
  assign clic__EVAL_131 = cbus__EVAL_44;
  assign clic__EVAL_136 = local_interrupts_0[6];
  assign clic__EVAL_89 = local_interrupts_0[63];
  assign sbus__EVAL_92 = tile__EVAL_24;
  assign clic__EVAL_4 = local_interrupts_0[73];
  assign cbus__EVAL_3 = debug_1__EVAL_9;
  assign cbus__EVAL_66 = sbus__EVAL_99;
  assign clic__EVAL_77 = cbus__EVAL_65;
  assign sbus__EVAL_84 = dummyClockGroupSourceNode__EVAL_0;
  assign clic__EVAL_109 = local_interrupts_0[125];
  assign clic__EVAL_107 = meip_0;
  assign sbus__EVAL_72 = cbus__EVAL_24;
  assign sbus__EVAL_46 = tile__EVAL_67;
  assign sbus__EVAL_133 = dummyClockGroupSourceNode__EVAL_3;
  assign sbus__EVAL_59 = tile__EVAL_30;
  assign sbus__EVAL_151 = fbus__EVAL_20;
  assign island_1__EVAL_6 = sbus__EVAL_23;
  assign cbus__EVAL_54 = debug_1__EVAL;
  assign clic__EVAL_149 = local_interrupts_0[74];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_2 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _EVAL_0 <= 1'h0;
    end else begin
      _EVAL_0 <= _EVAL_4;
    end
    if (reset) begin
      _EVAL_2 <= 1'h0;
    end else begin
      _EVAL_2 <= _EVAL;
    end
  end
endmodule
