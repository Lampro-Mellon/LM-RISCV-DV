//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_70_assert(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input  [3:0]  _EVAL_4,
  input         _EVAL_5,
  input  [3:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [13:0] _EVAL_10,
  input  [3:0]  _EVAL_11,
  input         _EVAL_12,
  input  [2:0]  _EVAL_13,
  input  [2:0]  _EVAL_14,
  input  [2:0]  _EVAL_15
);
  wire [4:0] _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire [22:0] _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  reg [2:0] _EVAL_26;
  reg [31:0] _RAND_0;
  wire  _EVAL_27;
  wire [1:0] _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire [13:0] _EVAL_31;
  wire  _EVAL_32;
  wire [31:0] _EVAL_33;
  wire  _EVAL_34;
  wire [5:0] _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  reg [5:0] _EVAL_43;
  reg [31:0] _RAND_1;
  wire  _EVAL_44;
  wire  _EVAL_45;
  reg [31:0] _EVAL_46;
  reg [31:0] _RAND_2;
  reg [5:0] _EVAL_47;
  reg [31:0] _RAND_3;
  reg [2:0] _EVAL_48;
  reg [31:0] _RAND_4;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire [3:0] _EVAL_57;
  wire  _EVAL_58;
  wire [6:0] _EVAL_59;
  wire  _EVAL_60;
  wire [5:0] _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  reg [2:0] _EVAL_69;
  reg [31:0] _RAND_5;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire [13:0] _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire [1:0] _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire [22:0] _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire [4:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire [14:0] _EVAL_108;
  wire  _EVAL_110;
  wire [7:0] _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire [1:0] _EVAL_123;
  wire [7:0] _EVAL_124;
  wire  _EVAL_126;
  wire [14:0] _EVAL_127;
  wire  _EVAL_128;
  wire [32:0] _EVAL_129;
  wire [7:0] _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire [13:0] _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire [6:0] _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire [5:0] _EVAL_154;
  wire [4:0] _EVAL_155;
  wire [7:0] _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire [7:0] _EVAL_161;
  wire  _EVAL_162;
  wire [4:0] _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_171;
  wire  _EVAL_172;
  reg [3:0] _EVAL_173;
  reg [31:0] _RAND_6;
  reg [4:0] _EVAL_174;
  reg [31:0] _RAND_7;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  reg [3:0] _EVAL_178;
  reg [31:0] _RAND_8;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  reg [13:0] _EVAL_192;
  reg [31:0] _RAND_9;
  wire  _EVAL_193;
  wire [6:0] _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire [14:0] _EVAL_209;
  wire  _EVAL_210;
  wire [4:0] _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire [3:0] _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire [3:0] _EVAL_220;
  wire [6:0] _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  reg [2:0] _EVAL_224;
  reg [31:0] _RAND_10;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire [5:0] _EVAL_229;
  wire [5:0] _EVAL_230;
  wire [7:0] _EVAL_231;
  wire  _EVAL_232;
  wire [5:0] _EVAL_233;
  wire  _EVAL_234;
  reg [2:0] _EVAL_235;
  reg [31:0] _RAND_11;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire [1:0] _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire [3:0] _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire [7:0] _EVAL_256;
  wire  _EVAL_257;
  wire [7:0] _EVAL_258;
  wire  _EVAL_259;
  wire [4:0] _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_263;
  reg [5:0] _EVAL_264;
  reg [31:0] _RAND_12;
  wire  _EVAL_265;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_266;
  wire  _EVAL_267;
  reg [5:0] _EVAL_268;
  reg [31:0] _RAND_13;
  wire [4:0] _EVAL_269;
  wire  _EVAL_270;
  wire [4:0] _EVAL_271;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_41 = _EVAL_13 == _EVAL_224;
  assign _EVAL_67 = _EVAL_8 & _EVAL_40;
  assign _EVAL_201 = _EVAL_250 | _EVAL_0;
  assign _EVAL_162 = _EVAL_94 | _EVAL_254;
  assign _EVAL_185 = _EVAL_162 | _EVAL_0;
  assign _EVAL_216 = _EVAL_193 | _EVAL_0;
  assign _EVAL_57 = ~_EVAL_214;
  assign _EVAL_184 = _EVAL_193 | _EVAL_92;
  assign _EVAL_251 = _EVAL_119 & _EVAL_52;
  assign _EVAL_87 = _EVAL_253 == 4'h0;
  assign _EVAL_129 = _EVAL_46 + 32'h1;
  assign _EVAL_186 = _EVAL_11 <= 4'h2;
  assign _EVAL_207 = _EVAL_10[0];
  assign _EVAL_82 = _EVAL_8 & _EVAL_150;
  assign _EVAL_40 = ~_EVAL_126;
  assign _EVAL_33 = _EVAL_129[31:0];
  assign _EVAL_76 = _EVAL_10 & _EVAL_142;
  assign _EVAL_91 = _EVAL_6 >= 4'h2;
  assign _EVAL_36 = ~_EVAL_1;
  assign _EVAL_27 = _EVAL_183 | _EVAL_0;
  assign _EVAL_183 = _EVAL_105 | _EVAL_24;
  assign _EVAL_237 = _EVAL_43 == 6'h0;
  assign _EVAL_108 = {1'b0,$signed(_EVAL_31)};
  assign _EVAL_38 = _EVAL_121 & _EVAL_188;
  assign _EVAL_49 = _EVAL_87 | _EVAL_0;
  assign _EVAL_229 = _EVAL_221[5:0];
  assign _EVAL_29 = _EVAL == 3'h1;
  assign _EVAL_110 = _EVAL <= 3'h6;
  assign _EVAL_127 = $signed(_EVAL_108) & -15'sh1000;
  assign _EVAL_106 = ~_EVAL_165;
  assign _EVAL_124 = _EVAL_113 ? _EVAL_156 : 8'h0;
  assign _EVAL_37 = _EVAL == 3'h4;
  assign _EVAL_120 = _EVAL_119 & _EVAL_72;
  assign _EVAL_34 = _EVAL_91 | _EVAL_0;
  assign _EVAL_233 = _EVAL_146[5:0];
  assign _EVAL_23 = _EVAL_186 & _EVAL_234;
  assign _EVAL_64 = _EVAL_96 | _EVAL_97;
  assign _EVAL_68 = ~_EVAL_232;
  assign _EVAL_248 = ~_EVAL_141;
  assign _EVAL_95 = _EVAL_149 | _EVAL_0;
  assign _EVAL_249 = ~_EVAL_34;
  assign _EVAL_179 = _EVAL_15 == 3'h3;
  assign _EVAL_169 = ~_EVAL_49;
  assign _EVAL_154 = _EVAL_231[7:2];
  assign _EVAL_126 = _EVAL_268 == 6'h0;
  assign _EVAL_114 = ~_EVAL_95;
  assign _EVAL_107 = ~_EVAL_225;
  assign _EVAL_159 = _EVAL_151 | _EVAL_0;
  assign _EVAL_65 = _EVAL_11 == _EVAL_178;
  assign _EVAL_236 = ~_EVAL_182;
  assign _EVAL_19 = ~_EVAL_206;
  assign _EVAL_208 = _EVAL_269[0];
  assign _EVAL_150 = _EVAL_15 == 3'h2;
  assign _EVAL_194 = _EVAL_268 - 6'h1;
  assign _EVAL_205 = _EVAL_28 == 2'h1;
  assign _EVAL_56 = _EVAL_28 == 2'h0;
  assign _EVAL_92 = _EVAL_181 & _EVAL_191;
  assign _EVAL_28 = _EVAL_13[2:1];
  assign _EVAL_16 = _EVAL_174 >> _EVAL_2;
  assign _EVAL_175 = _EVAL_174 != 5'h0;
  assign _EVAL_104 = _EVAL_9 & _EVAL_157;
  assign _EVAL_155 = _EVAL_103 | _EVAL_174;
  assign _EVAL_180 = ~_EVAL_18;
  assign _EVAL_84 = _EVAL_64 | _EVAL_0;
  assign _EVAL_166 = _EVAL_14 != 3'h0;
  assign _EVAL_165 = _EVAL_147 | _EVAL_0;
  assign _EVAL_24 = _EVAL_2 == 3'h4;
  assign _EVAL_130 = _EVAL_21[7:0];
  assign _EVAL_244 = _EVAL_208 | _EVAL_0;
  assign _EVAL_231 = ~_EVAL_130;
  assign _EVAL_204 = ~_EVAL_84;
  assign _EVAL_225 = _EVAL_134 | _EVAL_0;
  assign _EVAL_118 = ~_EVAL_139;
  assign _EVAL_80 = _EVAL_132 | _EVAL_137;
  assign _EVAL_53 = _EVAL_6 == _EVAL_173;
  assign _EVAL_45 = _EVAL_11[0];
  assign _EVAL_111 = _EVAL_78 ? _EVAL_161 : 8'h0;
  assign _EVAL_112 = _EVAL_184 | _EVAL_267;
  assign _EVAL_221 = _EVAL_43 - 6'h1;
  assign _EVAL_17 = _EVAL_199 & _EVAL_176;
  assign _EVAL_240 = _EVAL_15 == 3'h7;
  assign _EVAL_160 = _EVAL_190 | _EVAL_0;
  assign _EVAL_22 = ~_EVAL_159;
  assign _EVAL_202 = ~_EVAL_270;
  assign _EVAL_252 = _EVAL_15 == _EVAL_48;
  assign _EVAL_78 = _EVAL_133 & _EVAL_195;
  assign _EVAL_102 = _EVAL_252 | _EVAL_0;
  assign _EVAL_218 = ~_EVAL_175;
  assign _EVAL_103 = _EVAL_111[4:0];
  assign _EVAL_197 = _EVAL_184 | _EVAL_120;
  assign _EVAL_133 = _EVAL_3 & _EVAL_8;
  assign _EVAL_222 = _EVAL_11 <= 4'h8;
  assign _EVAL_59 = _EVAL_47 - 6'h1;
  assign _EVAL_88 = _EVAL_9 & _EVAL_37;
  assign _EVAL_60 = ~_EVAL_201;
  assign _EVAL_132 = _EVAL_205 | _EVAL_56;
  assign _EVAL_227 = ~_EVAL_86;
  assign _EVAL_25 = _EVAL_9 & _EVAL_152;
  assign _EVAL_83 = _EVAL_133 & _EVAL_126;
  assign _EVAL_215 = _EVAL_246 == 2'h1;
  assign _EVAL_265 = _EVAL_222 & _EVAL_234;
  assign _EVAL_234 = $signed(_EVAL_209) == 15'sh0;
  assign _EVAL_270 = _EVAL_166 | _EVAL_0;
  assign _EVAL_55 = _EVAL_8 & _EVAL_117;
  assign _EVAL_116 = _EVAL_110 | _EVAL_0;
  assign _EVAL_152 = ~_EVAL_237;
  assign _EVAL_134 = _EVAL_14 <= 3'h2;
  assign _EVAL_200 = _EVAL_41 | _EVAL_0;
  assign _EVAL_211 = ~_EVAL_260;
  assign _EVAL_157 = _EVAL == 3'h2;
  assign _EVAL_195 = _EVAL_47 == 6'h0;
  assign _EVAL_113 = _EVAL_38 & _EVAL_54;
  assign _EVAL_32 = _EVAL_15 == 3'h6;
  assign _EVAL_54 = ~_EVAL_203;
  assign _EVAL_247 = _EVAL_181 & _EVAL_199;
  assign _EVAL_164 = ~_EVAL_219;
  assign _EVAL_90 = ~_EVAL_131;
  assign _EVAL_96 = _EVAL_103 != _EVAL_260;
  assign _EVAL_35 = _EVAL_194[5:0];
  assign _EVAL_243 = _EVAL_8 & _EVAL_74;
  assign _EVAL_196 = _EVAL == 3'h0;
  assign _EVAL_105 = _EVAL_215 | _EVAL_144;
  assign _EVAL_191 = _EVAL_10[1];
  assign _EVAL_131 = _EVAL_62 | _EVAL_0;
  assign _EVAL_100 = _EVAL_8 & _EVAL_179;
  assign _EVAL_259 = ~_EVAL_116;
  assign _EVAL_117 = _EVAL_15 == 3'h5;
  assign _EVAL_167 = _EVAL_1 | _EVAL_0;
  assign _EVAL_189 = ~_EVAL_200;
  assign _EVAL_119 = _EVAL_89[0];
  assign _EVAL_139 = _EVAL_53 | _EVAL_0;
  assign _EVAL_21 = 23'hff << _EVAL_6;
  assign _EVAL_52 = _EVAL_199 & _EVAL_207;
  assign _EVAL_153 = _EVAL_228 | _EVAL_251;
  assign _EVAL_145 = _EVAL == _EVAL_235;
  assign _EVAL_62 = _EVAL_14 <= 3'h3;
  assign _EVAL_140 = _EVAL_9 & _EVAL_203;
  assign _EVAL_193 = _EVAL_11 >= 4'h2;
  assign _EVAL_89 = _EVAL_123 | 2'h1;
  assign _EVAL_123 = 2'h1 << _EVAL_45;
  assign _EVAL_241 = _EVAL_119 & _EVAL_17;
  assign _EVAL_239 = _EVAL_9 & _EVAL_136;
  assign _EVAL_70 = _EVAL_9 & _EVAL_196;
  assign _EVAL_61 = _EVAL_258[7:2];
  assign _EVAL_51 = _EVAL_65 | _EVAL_0;
  assign _EVAL_161 = 8'h1 << _EVAL_2;
  assign _EVAL_198 = _EVAL_133 | _EVAL_121;
  assign _EVAL_42 = ~_EVAL_27;
  assign _EVAL_72 = _EVAL_191 & _EVAL_207;
  assign _EVAL_213 = _EVAL_14 <= 3'h1;
  assign _EVAL_94 = _EVAL_218 | _EVAL_217;
  assign _EVAL_203 = _EVAL == 3'h6;
  assign _EVAL_141 = _EVAL_80 | _EVAL_0;
  assign _EVAL_99 = 23'hff << _EVAL_11;
  assign _EVAL_77 = ~_EVAL_20;
  assign _EVAL_151 = ~_EVAL_73;
  assign _EVAL_257 = ~_EVAL_167;
  assign _EVAL_30 = _EVAL_9 & _EVAL_29;
  assign _EVAL_214 = {_EVAL_197,_EVAL_112,_EVAL_153,_EVAL_245};
  assign _EVAL_163 = _EVAL_174 | _EVAL_103;
  assign _EVAL_171 = _EVAL_220 == 4'h0;
  assign _EVAL_138 = _EVAL_10 == _EVAL_192;
  assign _EVAL_136 = _EVAL == 3'h5;
  assign _EVAL_190 = _EVAL_14 == 3'h0;
  assign _EVAL_226 = ~_EVAL_185;
  assign _EVAL_269 = _EVAL_155 >> _EVAL_13;
  assign _EVAL_206 = _EVAL_81 | _EVAL_0;
  assign _EVAL_122 = ~_EVAL_212;
  assign _EVAL_263 = _EVAL_36 | _EVAL_0;
  assign _EVAL_168 = ~_EVAL_160;
  assign _EVAL_128 = _EVAL_103 != 5'h0;
  assign _EVAL_31 = _EVAL_10 ^ 14'h3000;
  assign _EVAL_254 = _EVAL_46 < plusarg_reader_out;
  assign _EVAL_143 = _EVAL_15 == 3'h4;
  assign _EVAL_256 = _EVAL_99[7:0];
  assign _EVAL_209 = _EVAL_127;
  assign _EVAL_260 = _EVAL_124[4:0];
  assign _EVAL_253 = ~_EVAL_4;
  assign _EVAL_172 = _EVAL_15 == 3'h1;
  assign _EVAL_181 = _EVAL_89[1];
  assign _EVAL_97 = ~_EVAL_128;
  assign _EVAL_230 = _EVAL_59[5:0];
  assign _EVAL_39 = ~_EVAL_102;
  assign _EVAL_146 = _EVAL_264 - 6'h1;
  assign _EVAL_58 = _EVAL_8 & _EVAL_240;
  assign _EVAL_255 = ~_EVAL_148;
  assign _EVAL_144 = _EVAL_246 == 2'h0;
  assign _EVAL_245 = _EVAL_228 | _EVAL_241;
  assign _EVAL_142 = {{6'd0}, _EVAL_258};
  assign _EVAL_219 = _EVAL_145 | _EVAL_0;
  assign _EVAL_271 = _EVAL_163 & _EVAL_211;
  assign _EVAL_246 = _EVAL_2[2:1];
  assign _EVAL_266 = _EVAL_8 & _EVAL_143;
  assign _EVAL_20 = _EVAL_265 | _EVAL_0;
  assign _EVAL_121 = _EVAL_7 & _EVAL_9;
  assign _EVAL_156 = 8'h1 << _EVAL_13;
  assign _EVAL_177 = ~_EVAL_216;
  assign _EVAL_71 = _EVAL_171 | _EVAL_0;
  assign _EVAL_50 = ~_EVAL_51;
  assign _EVAL_44 = _EVAL_14 == _EVAL_26;
  assign _EVAL_135 = _EVAL_8 & _EVAL_32;
  assign _EVAL_73 = _EVAL_16[0];
  assign _EVAL_187 = ~_EVAL_0;
  assign _EVAL_86 = _EVAL_138 | _EVAL_0;
  assign _EVAL_220 = _EVAL_4 & _EVAL_57;
  assign _EVAL_267 = _EVAL_119 & _EVAL_101;
  assign _EVAL_210 = _EVAL_8 & _EVAL_172;
  assign _EVAL_147 = _EVAL_4 == _EVAL_214;
  assign _EVAL_176 = ~_EVAL_207;
  assign _EVAL_137 = _EVAL_13 == 3'h4;
  assign _EVAL_188 = _EVAL_264 == 6'h0;
  assign _EVAL_232 = _EVAL_44 | _EVAL_0;
  assign _EVAL_81 = ~_EVAL_5;
  assign _EVAL_115 = ~_EVAL_244;
  assign _EVAL_238 = ~_EVAL_71;
  assign _EVAL_250 = _EVAL_76 == 14'h0;
  assign _EVAL_158 = _EVAL_14 <= 3'h4;
  assign _EVAL_149 = _EVAL_2 == _EVAL_69;
  assign _EVAL_261 = ~_EVAL_263;
  assign _EVAL_212 = _EVAL_158 | _EVAL_0;
  assign _EVAL_182 = _EVAL_213 | _EVAL_0;
  assign _EVAL_148 = _EVAL_23 | _EVAL_0;
  assign _EVAL_18 = _EVAL_15[2];
  assign _EVAL_101 = _EVAL_191 & _EVAL_176;
  assign _EVAL_199 = ~_EVAL_191;
  assign _EVAL_258 = ~_EVAL_256;
  assign _EVAL_74 = _EVAL_15 == 3'h0;
  assign _EVAL_217 = plusarg_reader_out == 32'h0;
  assign _EVAL_66 = _EVAL[0];
  assign _EVAL_228 = _EVAL_193 | _EVAL_247;
  assign _EVAL_223 = _EVAL_121 & _EVAL_237;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_26 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_43 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_46 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_47 = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_48 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_69 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_173 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_174 = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_178 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_192 = _RAND_9[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_224 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_235 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_264 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_268 = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_12) begin
    if (_EVAL_83) begin
      _EVAL_26 <= _EVAL_14;
    end
    if (_EVAL_0) begin
      _EVAL_43 <= 6'h0;
    end else if (_EVAL_121) begin
      if (_EVAL_237) begin
        if (_EVAL_66) begin
          _EVAL_43 <= _EVAL_154;
        end else begin
          _EVAL_43 <= 6'h0;
        end
      end else begin
        _EVAL_43 <= _EVAL_229;
      end
    end
    if (_EVAL_0) begin
      _EVAL_46 <= 32'h0;
    end else if (_EVAL_198) begin
      _EVAL_46 <= 32'h0;
    end else begin
      _EVAL_46 <= _EVAL_33;
    end
    if (_EVAL_0) begin
      _EVAL_47 <= 6'h0;
    end else if (_EVAL_133) begin
      if (_EVAL_195) begin
        if (_EVAL_180) begin
          _EVAL_47 <= _EVAL_61;
        end else begin
          _EVAL_47 <= 6'h0;
        end
      end else begin
        _EVAL_47 <= _EVAL_230;
      end
    end
    if (_EVAL_83) begin
      _EVAL_48 <= _EVAL_15;
    end
    if (_EVAL_83) begin
      _EVAL_69 <= _EVAL_2;
    end
    if (_EVAL_223) begin
      _EVAL_173 <= _EVAL_6;
    end
    if (_EVAL_0) begin
      _EVAL_174 <= 5'h0;
    end else begin
      _EVAL_174 <= _EVAL_271;
    end
    if (_EVAL_83) begin
      _EVAL_178 <= _EVAL_11;
    end
    if (_EVAL_83) begin
      _EVAL_192 <= _EVAL_10;
    end
    if (_EVAL_223) begin
      _EVAL_224 <= _EVAL_13;
    end
    if (_EVAL_223) begin
      _EVAL_235 <= _EVAL;
    end
    if (_EVAL_0) begin
      _EVAL_264 <= 6'h0;
    end else if (_EVAL_121) begin
      if (_EVAL_188) begin
        if (_EVAL_66) begin
          _EVAL_264 <= _EVAL_154;
        end else begin
          _EVAL_264 <= 6'h0;
        end
      end else begin
        _EVAL_264 <= _EVAL_233;
      end
    end
    if (_EVAL_0) begin
      _EVAL_268 <= 6'h0;
    end else if (_EVAL_133) begin
      if (_EVAL_126) begin
        if (_EVAL_180) begin
          _EVAL_268 <= _EVAL_61;
        end else begin
          _EVAL_268 <= 6'h0;
        end
      end else begin
        _EVAL_268 <= _EVAL_35;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d225f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45c35af2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7aa6654e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(226e002f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aec7e71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a677ba72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88c928f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbe53af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_255) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(970ebbf6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8770f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(830ade40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2294554)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d24cff6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_255) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f770474)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb4b6d9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6f29885)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b33750a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95ab6f67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8a8911f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19e14fe3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3839f84c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d2d70eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(657b1c90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f622af41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6401a3ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3734d537)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b265870d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cd6c9a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b949dae8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7203560c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b27281c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(108733e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f35e0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77695318)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(386f8685)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a908e56e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfa44e54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ab36b77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e7541fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee6fd95c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_255) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(beaa0312)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edf815a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dd498a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c09398ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(912c3685)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbad827e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(408c9fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9bf77a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(222b3f4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5892ee75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfc595fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bac90f97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e749b36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a86f99a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d33ac015)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca2e0917)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34aa63d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24ee2409)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(241a5747)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22a750e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8f045e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32b2fe64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fcf9d2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4e73ef6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df398e44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0d6b0fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3628509)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d46ad006)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48cd8221)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(750e1987)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e75c1b38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88c7d2e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5bc9a4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_255) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c3cf9dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a27faab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20b93a20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d0030ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba8bf8d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e860a636)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7848492)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
