//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_154_assert(
  input         _EVAL,
  input  [1:0]  _EVAL_1,
  input  [1:0]  _EVAL_3,
  input         _EVAL_16,
  input         _EVAL_42,
  input         _EVAL_43,
  input         _EVAL_49,
  input         _EVAL_59,
  input         _EVAL_63,
  input         _EVAL_93,
  input  [2:0]  _EVAL_98,
  input  [11:0] _EVAL_101,
  input  [7:0]  _EVAL_108,
  input  [1:0]  _EVAL_116,
  input  [1:0]  _EVAL_129,
  input         _EVAL_218,
  input         _EVAL_337,
  input         _EVAL_368,
  input         _EVAL_425,
  input         _EVAL_446,
  input         _EVAL_525,
  input         _EVAL_550,
  input         _EVAL_555,
  input         _EVAL_596,
  input         _EVAL_659,
  input         _EVAL_700,
  input         _EVAL_758,
  input         _EVAL_789,
  input         _EVAL_841,
  input         _EVAL_889,
  input         _EVAL_985,
  input         _EVAL_1071,
  input         _EVAL_1095,
  input         _EVAL_1114,
  input         _EVAL_1117,
  input         _EVAL_1127,
  input         _EVAL_1146,
  input  [7:0]  _EVAL_1267,
  input         _EVAL_1274,
  input         _EVAL_1278,
  input         _EVAL_1294,
  input         _EVAL_1414,
  input         _EVAL_1464,
  input         _EVAL_1475,
  input         _EVAL_1610,
  input         _EVAL_1619,
  input         _EVAL_1659,
  input         _EVAL_1681,
  input         _EVAL_1700,
  input         _EVAL_1717,
  input         _EVAL_1740,
  input         _EVAL_1771,
  input         _EVAL_1807,
  input         _EVAL_1830,
  input         _EVAL_1842,
  input         _EVAL_1878,
  input         _EVAL_1898,
  input         _EVAL_1939,
  input         _EVAL_1966,
  input         _EVAL_2002,
  input         _EVAL_2081,
  input         _EVAL_2127,
  input  [1:0]  _EVAL_2147,
  input         _EVAL_2182,
  input         _EVAL_2193,
  input  [7:0]  _EVAL_2251,
  input         _EVAL_2305,
  input         _EVAL_2345,
  input         _EVAL_2380,
  input         _EVAL_2394,
  input         _EVAL_2421,
  input         _EVAL_2423,
  input         _EVAL_2443,
  input         _EVAL_2454,
  input         _EVAL_2501,
  input         _EVAL_2536,
  input         _EVAL_2538,
  input         _EVAL_2567,
  input         _EVAL_2659,
  input         _EVAL_2670,
  input         _EVAL_2680,
  input         _EVAL_2746,
  input         _EVAL_2778,
  input         _EVAL_2789,
  input         _EVAL_2920,
  input         _EVAL_3063,
  input         _EVAL_3088,
  input         _EVAL_3147,
  input         _EVAL_3148,
  input         _EVAL_3169,
  input         _EVAL_3207,
  input         _EVAL_3210,
  input  [31:0] _EVAL_3254
);
  wire  _EVAL_144;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_150;
  wire  _EVAL_154;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_185;
  wire  _EVAL_188;
  wire  _EVAL_195;
  wire  _EVAL_213;
  wire  _EVAL_216;
  wire  _EVAL_222;
  wire  _EVAL_225;
  wire  _EVAL_229;
  wire  _EVAL_231;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_246;
  wire  _EVAL_248;
  wire  _EVAL_255;
  wire  _EVAL_257;
  wire  _EVAL_268;
  wire  _EVAL_271;
  wire  _EVAL_289;
  wire  _EVAL_295;
  wire  _EVAL_300;
  wire  _EVAL_307;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_318;
  wire  _EVAL_321;
  wire  _EVAL_323;
  wire  _EVAL_324;
  wire  _EVAL_342;
  wire  _EVAL_343;
  wire  _EVAL_347;
  wire  _EVAL_348;
  wire  _EVAL_349;
  wire  _EVAL_352;
  wire  _EVAL_355;
  wire  _EVAL_359;
  wire  _EVAL_360;
  wire  _EVAL_371;
  wire  _EVAL_372;
  wire  _EVAL_378;
  wire  _EVAL_384;
  wire  _EVAL_389;
  wire  _EVAL_392;
  wire  _EVAL_393;
  wire  _EVAL_395;
  wire  _EVAL_396;
  wire  _EVAL_398;
  wire  _EVAL_400;
  wire  _EVAL_403;
  wire  _EVAL_416;
  wire  _EVAL_418;
  wire  _EVAL_426;
  wire  _EVAL_433;
  wire  _EVAL_434;
  wire  _EVAL_443;
  wire  _EVAL_450;
  wire  _EVAL_455;
  wire  _EVAL_458;
  wire  _EVAL_462;
  wire  _EVAL_464;
  wire  _EVAL_465;
  wire  _EVAL_488;
  wire  _EVAL_496;
  wire  _EVAL_511;
  wire  _EVAL_516;
  wire  _EVAL_517;
  wire  _EVAL_518;
  wire  _EVAL_527;
  wire  _EVAL_528;
  wire  _EVAL_529;
  wire  _EVAL_530;
  wire  _EVAL_533;
  wire  _EVAL_536;
  wire  _EVAL_538;
  wire  _EVAL_541;
  wire  _EVAL_545;
  wire  _EVAL_548;
  wire  _EVAL_549;
  wire  _EVAL_569;
  wire  _EVAL_574;
  wire  _EVAL_575;
  wire  _EVAL_577;
  wire  _EVAL_579;
  wire  _EVAL_580;
  wire  _EVAL_585;
  wire  _EVAL_587;
  wire  _EVAL_592;
  wire  _EVAL_593;
  wire  _EVAL_595;
  wire  _EVAL_603;
  wire  _EVAL_604;
  wire  _EVAL_614;
  wire  _EVAL_623;
  wire  _EVAL_633;
  wire  _EVAL_636;
  wire  _EVAL_638;
  wire  _EVAL_643;
  wire  _EVAL_647;
  wire  _EVAL_651;
  wire  _EVAL_652;
  wire  _EVAL_654;
  wire  _EVAL_658;
  wire  _EVAL_664;
  wire  _EVAL_665;
  wire  _EVAL_676;
  wire  _EVAL_678;
  wire  _EVAL_682;
  wire  _EVAL_687;
  wire  _EVAL_689;
  wire  _EVAL_695;
  wire  _EVAL_696;
  wire  _EVAL_697;
  wire  _EVAL_709;
  wire  _EVAL_723;
  wire [1:0] _EVAL_725;
  wire  _EVAL_735;
  wire  _EVAL_738;
  wire  _EVAL_744;
  wire  _EVAL_747;
  wire  _EVAL_750;
  wire  _EVAL_755;
  wire  _EVAL_756;
  wire  _EVAL_757;
  wire  _EVAL_760;
  wire  _EVAL_783;
  wire  _EVAL_792;
  wire  _EVAL_794;
  wire  _EVAL_796;
  wire  _EVAL_797;
  wire  _EVAL_803;
  wire  _EVAL_812;
  wire  _EVAL_816;
  wire  _EVAL_823;
  wire  _EVAL_827;
  wire  _EVAL_831;
  wire  _EVAL_837;
  wire  _EVAL_838;
  wire  _EVAL_839;
  wire  _EVAL_842;
  wire  _EVAL_844;
  wire  _EVAL_846;
  wire  _EVAL_847;
  wire  _EVAL_848;
  wire  _EVAL_858;
  wire  _EVAL_863;
  wire  _EVAL_867;
  wire  _EVAL_868;
  wire  _EVAL_869;
  wire  _EVAL_881;
  wire  _EVAL_888;
  wire  _EVAL_893;
  wire  _EVAL_894;
  wire  _EVAL_900;
  wire  _EVAL_921;
  wire  _EVAL_929;
  wire  _EVAL_930;
  wire  _EVAL_931;
  wire  _EVAL_939;
  wire  _EVAL_940;
  wire  _EVAL_942;
  wire  _EVAL_945;
  wire  _EVAL_949;
  wire  _EVAL_951;
  wire  _EVAL_955;
  wire  _EVAL_958;
  wire  _EVAL_965;
  wire  _EVAL_983;
  wire  _EVAL_984;
  wire  _EVAL_987;
  wire  _EVAL_988;
  wire  _EVAL_989;
  wire  _EVAL_990;
  wire  _EVAL_991;
  wire  _EVAL_992;
  wire  _EVAL_994;
  wire  _EVAL_998;
  wire  _EVAL_999;
  wire  _EVAL_1002;
  wire  _EVAL_1003;
  wire  _EVAL_1005;
  wire  _EVAL_1008;
  wire  _EVAL_1014;
  wire  _EVAL_1022;
  wire  _EVAL_1025;
  wire  _EVAL_1028;
  wire  _EVAL_1034;
  wire  _EVAL_1038;
  wire  _EVAL_1041;
  wire  _EVAL_1043;
  wire  _EVAL_1046;
  wire  _EVAL_1048;
  wire  _EVAL_1049;
  wire  _EVAL_1053;
  wire  _EVAL_1057;
  wire  _EVAL_1059;
  wire  _EVAL_1066;
  wire  _EVAL_1067;
  wire  _EVAL_1068;
  wire  _EVAL_1072;
  wire  _EVAL_1076;
  wire  _EVAL_1082;
  wire  _EVAL_1084;
  wire  _EVAL_1086;
  wire  _EVAL_1091;
  wire  _EVAL_1096;
  wire  _EVAL_1100;
  wire  _EVAL_1102;
  wire  _EVAL_1103;
  wire  _EVAL_1109;
  wire  _EVAL_1111;
  wire  _EVAL_1135;
  wire  _EVAL_1138;
  wire  _EVAL_1139;
  wire  _EVAL_1140;
  wire  _EVAL_1145;
  wire  _EVAL_1147;
  wire  _EVAL_1151;
  wire  _EVAL_1153;
  wire  _EVAL_1155;
  wire  _EVAL_1160;
  wire  _EVAL_1161;
  wire  _EVAL_1166;
  wire  _EVAL_1167;
  wire  _EVAL_1168;
  wire  _EVAL_1170;
  wire  _EVAL_1178;
  wire  _EVAL_1180;
  wire  _EVAL_1182;
  wire  _EVAL_1186;
  wire  _EVAL_1188;
  wire  _EVAL_1196;
  wire  _EVAL_1198;
  wire  _EVAL_1206;
  wire  _EVAL_1210;
  wire  _EVAL_1211;
  wire  _EVAL_1219;
  wire  _EVAL_1222;
  wire  _EVAL_1227;
  wire  _EVAL_1232;
  wire  _EVAL_1234;
  wire  _EVAL_1237;
  wire  _EVAL_1242;
  wire  _EVAL_1249;
  wire  _EVAL_1250;
  wire  _EVAL_1253;
  wire  _EVAL_1254;
  wire  _EVAL_1256;
  wire  _EVAL_1257;
  wire  _EVAL_1260;
  wire  _EVAL_1262;
  wire  _EVAL_1263;
  wire  _EVAL_1284;
  wire  _EVAL_1285;
  wire  _EVAL_1301;
  wire  _EVAL_1304;
  wire  _EVAL_1307;
  wire  _EVAL_1314;
  wire  _EVAL_1316;
  wire  _EVAL_1320;
  wire  _EVAL_1336;
  wire  _EVAL_1341;
  wire  _EVAL_1342;
  wire  _EVAL_1345;
  wire  _EVAL_1346;
  wire  _EVAL_1352;
  wire  _EVAL_1357;
  wire  _EVAL_1358;
  wire  _EVAL_1361;
  wire  _EVAL_1363;
  wire  _EVAL_1368;
  wire  _EVAL_1370;
  wire  _EVAL_1373;
  wire  _EVAL_1374;
  wire  _EVAL_1378;
  wire  _EVAL_1402;
  wire  _EVAL_1406;
  wire  _EVAL_1425;
  wire  _EVAL_1426;
  wire  _EVAL_1430;
  wire  _EVAL_1431;
  wire  _EVAL_1432;
  wire  _EVAL_1434;
  wire  _EVAL_1437;
  wire  _EVAL_1438;
  wire  _EVAL_1442;
  wire  _EVAL_1443;
  wire  _EVAL_1445;
  wire  _EVAL_1449;
  wire  _EVAL_1456;
  wire  _EVAL_1461;
  wire  _EVAL_1471;
  wire  _EVAL_1477;
  wire  _EVAL_1481;
  wire  _EVAL_1483;
  wire  _EVAL_1496;
  wire  _EVAL_1497;
  wire  _EVAL_1498;
  wire  _EVAL_1504;
  wire  _EVAL_1509;
  wire  _EVAL_1511;
  wire  _EVAL_1516;
  wire  _EVAL_1521;
  wire  _EVAL_1522;
  wire  _EVAL_1524;
  wire  _EVAL_1527;
  wire  _EVAL_1535;
  wire  _EVAL_1536;
  wire  _EVAL_1538;
  wire  _EVAL_1540;
  wire  _EVAL_1542;
  wire  _EVAL_1552;
  wire  _EVAL_1555;
  wire  _EVAL_1556;
  wire  _EVAL_1561;
  wire  _EVAL_1565;
  wire  _EVAL_1570;
  wire  _EVAL_1572;
  wire  _EVAL_1574;
  wire  _EVAL_1575;
  wire  _EVAL_1576;
  wire  _EVAL_1582;
  wire  _EVAL_1583;
  wire  _EVAL_1597;
  wire  _EVAL_1598;
  wire  _EVAL_1602;
  wire  _EVAL_1605;
  wire  _EVAL_1606;
  wire  _EVAL_1607;
  wire  _EVAL_1612;
  wire  _EVAL_1613;
  wire  _EVAL_1615;
  wire  _EVAL_1622;
  wire  _EVAL_1623;
  wire  _EVAL_1625;
  wire  _EVAL_1629;
  wire  _EVAL_1633;
  wire  _EVAL_1638;
  wire  _EVAL_1640;
  wire  _EVAL_1641;
  wire  _EVAL_1645;
  wire  _EVAL_1648;
  wire  _EVAL_1650;
  wire  _EVAL_1652;
  wire  _EVAL_1653;
  wire  _EVAL_1654;
  wire  _EVAL_1655;
  wire  _EVAL_1661;
  wire  _EVAL_1663;
  wire  _EVAL_1667;
  wire  _EVAL_1668;
  wire  _EVAL_1670;
  wire  _EVAL_1674;
  wire  _EVAL_1687;
  wire  _EVAL_1691;
  wire  _EVAL_1696;
  wire  _EVAL_1703;
  wire  _EVAL_1708;
  wire  _EVAL_1709;
  wire  _EVAL_1711;
  wire  _EVAL_1712;
  wire  _EVAL_1718;
  wire  _EVAL_1726;
  wire  _EVAL_1728;
  wire  _EVAL_1732;
  wire  _EVAL_1733;
  wire  _EVAL_1741;
  wire  _EVAL_1745;
  wire  _EVAL_1747;
  wire  _EVAL_1748;
  wire  _EVAL_1754;
  wire  _EVAL_1765;
  wire  _EVAL_1768;
  wire  _EVAL_1769;
  wire  _EVAL_1775;
  wire  _EVAL_1779;
  wire  _EVAL_1780;
  wire  _EVAL_1784;
  wire  _EVAL_1785;
  wire  _EVAL_1786;
  wire  _EVAL_1791;
  wire  _EVAL_1797;
  wire  _EVAL_1798;
  wire  _EVAL_1801;
  wire  _EVAL_1804;
  wire  _EVAL_1806;
  wire  _EVAL_1809;
  wire  _EVAL_1810;
  wire  _EVAL_1820;
  wire  _EVAL_1822;
  wire  _EVAL_1824;
  wire  _EVAL_1826;
  wire  _EVAL_1827;
  wire  _EVAL_1828;
  wire  _EVAL_1833;
  wire  _EVAL_1836;
  wire  _EVAL_1840;
  wire  _EVAL_1845;
  wire  _EVAL_1854;
  wire  _EVAL_1855;
  wire  _EVAL_1865;
  wire  _EVAL_1867;
  wire  _EVAL_1870;
  wire  _EVAL_1874;
  wire  _EVAL_1889;
  wire  _EVAL_1891;
  wire  _EVAL_1897;
  wire  _EVAL_1902;
  wire  _EVAL_1903;
  wire  _EVAL_1904;
  wire  _EVAL_1921;
  wire  _EVAL_1922;
  wire  _EVAL_1923;
  wire  _EVAL_1926;
  wire  _EVAL_1938;
  wire  _EVAL_1943;
  wire  _EVAL_1950;
  wire  _EVAL_1954;
  wire  _EVAL_1959;
  wire  _EVAL_1962;
  wire  _EVAL_1968;
  wire  _EVAL_1973;
  wire  _EVAL_1981;
  wire  _EVAL_1990;
  wire  _EVAL_1997;
  wire  _EVAL_2004;
  wire  _EVAL_2007;
  wire  _EVAL_2010;
  wire  _EVAL_2012;
  wire  _EVAL_2017;
  wire  _EVAL_2018;
  wire  _EVAL_2024;
  wire  _EVAL_2025;
  wire  _EVAL_2027;
  wire  _EVAL_2033;
  wire  _EVAL_2035;
  wire  _EVAL_2036;
  wire  _EVAL_2038;
  wire  _EVAL_2040;
  wire  _EVAL_2052;
  wire  _EVAL_2055;
  wire  _EVAL_2066;
  wire  _EVAL_2068;
  wire  _EVAL_2071;
  wire  _EVAL_2074;
  wire  _EVAL_2078;
  wire  _EVAL_2079;
  wire  _EVAL_2080;
  wire  _EVAL_2082;
  wire  _EVAL_2091;
  wire  _EVAL_2099;
  wire  _EVAL_2103;
  wire  _EVAL_2104;
  wire  _EVAL_2112;
  wire  _EVAL_2116;
  wire  _EVAL_2120;
  wire  _EVAL_2132;
  wire  _EVAL_2136;
  wire  _EVAL_2137;
  wire  _EVAL_2140;
  wire  _EVAL_2143;
  wire  _EVAL_2144;
  wire  _EVAL_2153;
  wire  _EVAL_2174;
  wire  _EVAL_2176;
  wire  _EVAL_2180;
  wire [1:0] _EVAL_2181;
  wire  _EVAL_2183;
  wire  _EVAL_2187;
  wire  _EVAL_2197;
  wire  _EVAL_2198;
  wire  _EVAL_2207;
  wire  _EVAL_2214;
  wire  _EVAL_2220;
  wire  _EVAL_2226;
  wire  _EVAL_2230;
  wire  _EVAL_2238;
  wire  _EVAL_2240;
  wire  _EVAL_2242;
  wire  _EVAL_2243;
  wire  _EVAL_2244;
  wire  _EVAL_2245;
  wire  _EVAL_2246;
  wire  _EVAL_2249;
  wire  _EVAL_2253;
  wire  _EVAL_2254;
  wire  _EVAL_2259;
  wire  _EVAL_2266;
  wire  _EVAL_2272;
  wire  _EVAL_2275;
  wire  _EVAL_2282;
  wire  _EVAL_2283;
  wire  _EVAL_2292;
  wire  _EVAL_2301;
  wire  _EVAL_2303;
  wire  _EVAL_2316;
  wire  _EVAL_2329;
  wire  _EVAL_2336;
  wire  _EVAL_2337;
  wire  _EVAL_2339;
  wire  _EVAL_2341;
  wire  _EVAL_2353;
  wire  _EVAL_2365;
  wire  _EVAL_2368;
  wire  _EVAL_2370;
  wire  _EVAL_2371;
  wire  _EVAL_2373;
  wire  _EVAL_2377;
  wire  _EVAL_2390;
  wire  _EVAL_2399;
  wire  _EVAL_2403;
  wire  _EVAL_2415;
  wire  _EVAL_2417;
  wire  _EVAL_2426;
  wire  _EVAL_2432;
  wire  _EVAL_2436;
  wire  _EVAL_2439;
  wire  _EVAL_2450;
  wire  _EVAL_2456;
  wire  _EVAL_2465;
  wire  _EVAL_2473;
  wire  _EVAL_2476;
  wire  _EVAL_2478;
  wire  _EVAL_2491;
  wire  _EVAL_2497;
  wire  _EVAL_2499;
  wire  _EVAL_2503;
  wire  _EVAL_2512;
  wire  _EVAL_2514;
  wire  _EVAL_2515;
  wire  _EVAL_2520;
  wire  _EVAL_2522;
  wire  _EVAL_2526;
  wire  _EVAL_2530;
  wire  _EVAL_2531;
  wire  _EVAL_2547;
  wire  _EVAL_2552;
  wire  _EVAL_2553;
  wire  _EVAL_2555;
  wire  _EVAL_2556;
  wire  _EVAL_2560;
  wire  _EVAL_2565;
  wire  _EVAL_2566;
  wire  _EVAL_2570;
  wire  _EVAL_2585;
  wire  _EVAL_2596;
  wire  _EVAL_2598;
  wire  _EVAL_2600;
  wire  _EVAL_2601;
  wire  _EVAL_2603;
  wire  _EVAL_2610;
  wire  _EVAL_2612;
  wire [2:0] _EVAL_2618;
  wire  _EVAL_2619;
  wire  _EVAL_2623;
  wire  _EVAL_2625;
  wire  _EVAL_2626;
  wire  _EVAL_2630;
  wire  _EVAL_2633;
  wire  _EVAL_2634;
  wire  _EVAL_2639;
  wire  _EVAL_2642;
  wire  _EVAL_2643;
  wire  _EVAL_2664;
  wire  _EVAL_2672;
  wire  _EVAL_2675;
  wire  _EVAL_2679;
  wire  _EVAL_2682;
  wire  _EVAL_2683;
  wire  _EVAL_2684;
  wire  _EVAL_2693;
  wire  _EVAL_2700;
  wire  _EVAL_2706;
  wire  _EVAL_2714;
  wire  _EVAL_2718;
  wire  _EVAL_2724;
  wire  _EVAL_2726;
  wire  _EVAL_2734;
  wire  _EVAL_2739;
  wire  _EVAL_2742;
  wire  _EVAL_2749;
  wire  _EVAL_2751;
  wire  _EVAL_2756;
  wire  _EVAL_2758;
  wire  _EVAL_2762;
  wire  _EVAL_2763;
  wire  _EVAL_2768;
  wire  _EVAL_2773;
  wire  _EVAL_2777;
  wire  _EVAL_2780;
  wire  _EVAL_2782;
  wire  _EVAL_2783;
  wire  _EVAL_2785;
  wire  _EVAL_2795;
  wire  _EVAL_2797;
  wire  _EVAL_2798;
  wire  _EVAL_2800;
  wire  _EVAL_2807;
  wire  _EVAL_2811;
  wire  _EVAL_2812;
  wire  _EVAL_2820;
  wire  _EVAL_2826;
  wire  _EVAL_2829;
  wire  _EVAL_2832;
  wire  _EVAL_2835;
  wire  _EVAL_2839;
  wire  _EVAL_2847;
  wire  _EVAL_2852;
  wire  _EVAL_2855;
  wire  _EVAL_2864;
  wire  _EVAL_2871;
  wire  _EVAL_2874;
  wire  _EVAL_2879;
  wire  _EVAL_2882;
  wire  _EVAL_2883;
  wire  _EVAL_2885;
  wire  _EVAL_2886;
  wire  _EVAL_2891;
  wire  _EVAL_2892;
  wire  _EVAL_2894;
  wire  _EVAL_2897;
  wire  _EVAL_2905;
  wire  _EVAL_2910;
  wire  _EVAL_2911;
  wire  _EVAL_2912;
  wire  _EVAL_2916;
  wire  _EVAL_2921;
  wire  _EVAL_2922;
  wire  _EVAL_2923;
  wire  _EVAL_2924;
  wire  _EVAL_2925;
  wire  _EVAL_2926;
  wire  _EVAL_2930;
  wire  _EVAL_2932;
  wire  _EVAL_2935;
  wire  _EVAL_2936;
  wire  _EVAL_2943;
  wire  _EVAL_2948;
  wire  _EVAL_2952;
  wire  _EVAL_2957;
  wire  _EVAL_2959;
  wire  _EVAL_2961;
  wire  _EVAL_2963;
  wire  _EVAL_2967;
  wire  _EVAL_2969;
  wire  _EVAL_2973;
  wire  _EVAL_2979;
  wire  _EVAL_2980;
  wire  _EVAL_2982;
  wire  _EVAL_2984;
  wire  _EVAL_2995;
  wire  _EVAL_2997;
  wire  _EVAL_3001;
  wire  _EVAL_3003;
  wire  _EVAL_3004;
  wire  _EVAL_3009;
  wire  _EVAL_3010;
  wire  _EVAL_3019;
  wire  _EVAL_3023;
  wire  _EVAL_3024;
  wire  _EVAL_3028;
  wire  _EVAL_3032;
  wire  _EVAL_3038;
  wire  _EVAL_3041;
  wire  _EVAL_3045;
  wire  _EVAL_3050;
  wire  _EVAL_3061;
  wire  _EVAL_3071;
  wire  _EVAL_3072;
  wire  _EVAL_3077;
  wire  _EVAL_3083;
  wire  _EVAL_3085;
  wire  _EVAL_3092;
  wire  _EVAL_3094;
  wire  _EVAL_3103;
  wire  _EVAL_3104;
  wire  _EVAL_3107;
  wire  _EVAL_3108;
  wire  _EVAL_3111;
  wire  _EVAL_3118;
  wire  _EVAL_3126;
  wire  _EVAL_3130;
  wire  _EVAL_3135;
  wire  _EVAL_3138;
  wire  _EVAL_3141;
  wire  _EVAL_3145;
  wire  _EVAL_3146;
  wire  _EVAL_3154;
  wire  _EVAL_3155;
  wire  _EVAL_3159;
  wire  _EVAL_3174;
  wire  _EVAL_3185;
  wire  _EVAL_3188;
  wire  _EVAL_3190;
  wire  _EVAL_3192;
  wire  _EVAL_3200;
  wire  _EVAL_3212;
  wire  _EVAL_3220;
  wire  _EVAL_3221;
  wire  _EVAL_3222;
  wire  _EVAL_3223;
  wire  _EVAL_3226;
  wire  _EVAL_3232;
  wire  _EVAL_3234;
  wire  _EVAL_3238;
  wire  _EVAL_3240;
  wire  _EVAL_3241;
  wire  _EVAL_3244;
  wire  _EVAL_3247;
  wire  _EVAL_3252;
  wire  _EVAL_3253;
  assign _EVAL_1779 = _EVAL_2930 & _EVAL_695;
  assign _EVAL_2684 = _EVAL_101 == 12'h337;
  assign _EVAL_2679 = _EVAL_101 == 12'h32d;
  assign _EVAL_1434 = _EVAL_2930 & _EVAL_3001;
  assign _EVAL_2074 = ~_EVAL_1842;
  assign _EVAL_2136 = _EVAL_848 | _EVAL_1661;
  assign _EVAL_545 = _EVAL_3254 == 32'h8000008b;
  assign _EVAL_1497 = _EVAL_101 == 12'hc9c;
  assign _EVAL_797 = _EVAL_2930 & _EVAL_2193;
  assign _EVAL_1810 = ~_EVAL_2025;
  assign _EVAL_2565 = _EVAL_101 == 12'hc12;
  assign _EVAL_3159 = _EVAL_1103 | _EVAL_1607;
  assign _EVAL_3083 = _EVAL_2930 & _EVAL_147;
  assign _EVAL_1100 = _EVAL_2930 & _EVAL_1155;
  assign _EVAL_2879 = _EVAL_101 == 12'hb9e;
  assign _EVAL_1345 = _EVAL_2930 & _EVAL_371;
  assign _EVAL_1357 = _EVAL_2443 | _EVAL_1304;
  assign _EVAL_1378 = _EVAL_1511 & _EVAL_213;
  assign _EVAL_987 = _EVAL_3254 == 32'h80000021;
  assign _EVAL_2763 = _EVAL_101 == 12'h3bd;
  assign _EVAL_403 = _EVAL_101 == 12'hc1c;
  assign _EVAL_1014 = _EVAL_2630 | _EVAL_2664;
  assign _EVAL_2244 = _EVAL_638 | _EVAL_1968;
  assign _EVAL_175 = _EVAL_3159 | _EVAL_1867;
  assign _EVAL_1346 = _EVAL_2930 & _EVAL_723;
  assign _EVAL_696 = _EVAL_3254 == 32'h8000002b;
  assign _EVAL_1938 = _EVAL_101 == 12'hb9b;
  assign _EVAL_2329 = _EVAL_3223 & _EVAL_2567;
  assign _EVAL_2995 = _EVAL_129 == _EVAL_116;
  assign _EVAL_2749 = _EVAL_2930 & _EVAL_2780;
  assign _EVAL_347 = _EVAL_2930 & _EVAL_1830;
  assign _EVAL_2116 = _EVAL_2930 & _EVAL_2682;
  assign _EVAL_2894 = _EVAL_101 == 12'hc08;
  assign _EVAL_735 = _EVAL_3254 == 32'h8000007c;
  assign _EVAL_1316 = _EVAL_101 == 12'h3b4;
  assign _EVAL_1654 = _EVAL_3254 == 32'h80000084;
  assign _EVAL_1570 = _EVAL_1613 & _EVAL_1464;
  assign _EVAL_3154 = _EVAL_2567 & _EVAL_1140;
  assign _EVAL_1691 = _EVAL_3254 == 32'h80000086;
  assign _EVAL_1445 = _EVAL_101 == 12'hc0d;
  assign _EVAL_518 = _EVAL_2930 & _EVAL_2980;
  assign _EVAL_2963 = _EVAL_3254 == 32'h80000036;
  assign _EVAL_2984 = _EVAL_395 | _EVAL_812;
  assign _EVAL_1997 = _EVAL_3254 == 32'h80000061;
  assign _EVAL_1432 = _EVAL_101 == 12'hc13;
  assign _EVAL_757 = _EVAL_2930 & _EVAL_1926;
  assign _EVAL_989 = _EVAL_101 == 12'hb93;
  assign _EVAL_2403 = _EVAL_1854 | _EVAL_939;
  assign _EVAL_2967 = _EVAL_2530 | _EVAL_2007;
  assign _EVAL_1504 = _EVAL_2930 & _EVAL_709;
  assign _EVAL_1768 = _EVAL_949 & _EVAL_659;
  assign _EVAL_676 = _EVAL_3254 == 32'h80000056;
  assign _EVAL_3071 = _EVAL_3254 == 32'h80000080;
  assign _EVAL_3185 = _EVAL_101 == 12'hb14;
  assign _EVAL_1084 = _EVAL_2930 & _EVAL_2789;
  assign _EVAL_462 = _EVAL_1461 | _EVAL_796;
  assign _EVAL_2456 = _EVAL_3254 == 32'h80000023;
  assign _EVAL_2370 = _EVAL_3254 == 32'h80000065;
  assign _EVAL_1135 = _EVAL_3254 == 32'h8000006c;
  assign _EVAL_3023 = _EVAL_318 & _EVAL_2882;
  assign _EVAL_2820 = _EVAL_1511 & _EVAL_633;
  assign _EVAL_1182 = _EVAL_1511 & _EVAL_2253;
  assign _EVAL_2036 = _EVAL_1511 & _EVAL_2417;
  assign _EVAL_2187 = _EVAL_516 & _EVAL_2567;
  assign _EVAL_847 = _EVAL_101 == 12'hb0b;
  assign _EVAL_839 = _EVAL_2930 & _EVAL_1845;
  assign _EVAL_2979 = _EVAL_3254 == 32'h80000070;
  assign _EVAL_2339 = _EVAL_43 & _EVAL_889;
  assign _EVAL_464 = _EVAL_2930 & _EVAL_841;
  assign _EVAL_2520 = _EVAL_3254 == 32'h8000008c;
  assign _EVAL_1598 = _EVAL_2930 & _EVAL_654;
  assign _EVAL_1687 = _EVAL_2336 | _EVAL_2811;
  assign _EVAL_1645 = _EVAL_2930 & _EVAL_1025;
  assign _EVAL_3028 = _EVAL_2930 & _EVAL_1703;
  assign _EVAL_1561 = _EVAL_3254 == 32'h7;
  assign _EVAL_1301 = _EVAL_101 == 12'hc10;
  assign _EVAL_2734 = _EVAL_3254 == 32'h80000052;
  assign _EVAL_1222 = _EVAL_1921 | _EVAL_1641;
  assign _EVAL_271 = _EVAL_1234 | _EVAL_1691;
  assign _EVAL_222 = _EVAL_101 == 12'hb99;
  assign _EVAL_1797 = _EVAL_101 == 12'h33a;
  assign _EVAL_1754 = _EVAL_2932 | _EVAL_1897;
  assign _EVAL_2724 = _EVAL_3254 == 32'h8000004b;
  assign _EVAL_1139 = _EVAL_2897 | _EVAL_2035;
  assign _EVAL_2491 = _EVAL_101 == 12'hc86;
  assign _EVAL_2839 = _EVAL_1602 | _EVAL_3190;
  assign _EVAL_1950 = _EVAL_1511 & _EVAL_2423;
  assign _EVAL_1865 = _EVAL_3254 == 32'h80000073;
  assign _EVAL_1667 = _EVAL_2567 & _EVAL_2948;
  assign _EVAL_392 = _EVAL_1511 & _EVAL_1497;
  assign _EVAL_1227 = _EVAL_2930 & _EVAL_1797;
  assign _EVAL_592 = _EVAL_129 != _EVAL_116;
  assign _EVAL_1509 = _EVAL_2567 & _EVAL_1368;
  assign _EVAL_324 = _EVAL_2930 & _EVAL_1747;
  assign _EVAL_575 = _EVAL_2930 & _EVAL_1153;
  assign _EVAL_1798 = _EVAL_1198 | _EVAL_2734;
  assign _EVAL_654 = _EVAL_101 == 12'h330;
  assign _EVAL_213 = _EVAL_101 == 12'hc17;
  assign _EVAL_2514 = _EVAL_101 == 12'hb09;
  assign _EVAL_1791 = _EVAL_3254 == 32'h80000060;
  assign _EVAL_1341 = _EVAL_318 & _EVAL_2874;
  assign _EVAL_1443 = _EVAL_2930 & _EVAL_2670;
  assign _EVAL_1425 = _EVAL_101 == 12'hb06;
  assign _EVAL_869 = ~_EVAL_93;
  assign _EVAL_3108 = _EVAL_3254 == 32'h8000004f;
  assign _EVAL_837 = _EVAL_2596 & _EVAL_1414;
  assign _EVAL_2826 = _EVAL_2905 | _EVAL_2207;
  assign _EVAL_1153 = _EVAL_101 == 12'hb0d;
  assign _EVAL_1822 = _EVAL_1048 | _EVAL_2714;
  assign _EVAL_1166 = _EVAL_101 == 12'h32a;
  assign _EVAL_1806 = _EVAL_3254 == 32'h80000075;
  assign _EVAL_652 = _EVAL_101 == 12'hb9c;
  assign _EVAL_2476 = _EVAL_1511 & _EVAL_239;
  assign _EVAL_2530 = _EVAL_195 | _EVAL_1806;
  assign _EVAL_2052 = _EVAL_101 == 12'hc9f;
  assign _EVAL_984 = _EVAL_101 == 12'hb1e;
  assign _EVAL_2959 = _EVAL_3254 == 32'h80000051;
  assign _EVAL_2365 = _EVAL_2930 & _EVAL_1425;
  assign _EVAL_1263 = _EVAL_2751 | _EVAL_1791;
  assign _EVAL_2071 = _EVAL_1284 | _EVAL_2439;
  assign _EVAL_3188 = _EVAL_101 == 12'hb1b;
  assign _EVAL_894 = _EVAL_1232 | _EVAL_3004;
  assign _EVAL_488 = _EVAL_2930 & _EVAL_1358;
  assign _EVAL_154 = _EVAL_3254 == 32'h80000007;
  assign _EVAL_1711 = _EVAL_3254 == 32'h80000019;
  assign _EVAL_1652 = _EVAL_3254 == 32'h8000003e;
  assign _EVAL_2798 = _EVAL_1068 | _EVAL_1552;
  assign _EVAL_2253 = _EVAL_101 == 12'hc8c;
  assign _EVAL_2948 = _EVAL_3254 == 32'hb;
  assign _EVAL_1943 = _EVAL_3254 == 32'h8000006b;
  assign _EVAL_1041 = _EVAL_101 == 12'hc0f;
  assign _EVAL_2811 = _EVAL_3254 == 32'h8000003d;
  assign _EVAL_433 = _EVAL_1 == _EVAL_129;
  assign _EVAL_1712 = _EVAL_2930 & _EVAL_1166;
  assign _EVAL_1498 = _EVAL_2930 & _EVAL_2718;
  assign _EVAL_2112 = _EVAL_3254 == 32'h2;
  assign _EVAL_2176 = _EVAL_400 & _EVAL_2567;
  assign _EVAL_2618 = _EVAL_2181 + _EVAL_725;
  assign _EVAL_2104 = _EVAL_3254 == 32'h8000007f;
  assign _EVAL_723 = _EVAL_101 == 12'hb8d;
  assign _EVAL_2892 = _EVAL_647 | _EVAL_831;
  assign _EVAL_2783 = _EVAL_3254 == 32'h80000035;
  assign _EVAL_2639 = _EVAL_101 == 12'hb0e;
  assign _EVAL_2503 = _EVAL_2930 & _EVAL_3061;
  assign _EVAL_2905 = _EVAL_1798 | _EVAL_2969;
  assign _EVAL_1091 = _EVAL_2930 & _EVAL_1114;
  assign _EVAL_3234 = _EVAL_3254 == 32'h80000011;
  assign _EVAL_528 = _EVAL_101 == 12'hb8e;
  assign _EVAL_2066 = _EVAL_2930 & _EVAL_2514;
  assign _EVAL_389 = _EVAL_2570 & _EVAL_3241;
  assign _EVAL_750 = _EVAL_2243 | _EVAL_1623;
  assign _EVAL_1552 = _EVAL_3254 == 32'h8000001e;
  assign _EVAL_1556 = _EVAL_1575 | _EVAL_1711;
  assign _EVAL_580 = _EVAL_101 == 12'h3b9;
  assign _EVAL_1607 = _EVAL_3254 == 32'h8000003a;
  assign _EVAL_1728 = _EVAL_2912 & _EVAL_827;
  assign _EVAL_1874 = _EVAL_2930 & _EVAL_3226;
  assign _EVAL_2782 = _EVAL_318 & _EVAL_1922;
  assign _EVAL_658 = _EVAL_3254 == 32'h8000000c;
  assign _EVAL_595 = _EVAL_2421 | _EVAL_218;
  assign _EVAL_931 = _EVAL_2930 & _EVAL_2879;
  assign _EVAL_2923 = _EVAL_1357 | _EVAL_63;
  assign _EVAL_1034 = _EVAL_3254 == 32'h80000029;
  assign _EVAL_2952 = _EVAL_2930 & _EVAL_1700;
  assign _EVAL_678 = _EVAL_101 == 12'hc1e;
  assign _EVAL_838 = _EVAL_1511 & _EVAL_2341;
  assign _EVAL_858 = _EVAL_1263 | _EVAL_1997;
  assign _EVAL_455 = _EVAL_2930 & _EVAL_396;
  assign _EVAL_1336 = _EVAL_1511 & _EVAL_596;
  assign _EVAL_323 = _EVAL_101 == 12'h327;
  assign _EVAL_816 = _EVAL_101 == 12'hb1c;
  assign _EVAL_2623 = _EVAL_1511 & _EVAL_2432;
  assign _EVAL_2642 = _EVAL_2531 | _EVAL_2104;
  assign _EVAL_1854 = _EVAL_2515 | _EVAL_225;
  assign _EVAL_2980 = _EVAL_101 == 12'hb0c;
  assign _EVAL_536 = _EVAL_2930 & _EVAL_1855;
  assign _EVAL_2040 = _EVAL_3254 == 32'h80000059;
  assign _EVAL_1922 = _EVAL_1842 & _EVAL_1274;
  assign _EVAL_842 = _EVAL_2283 & _EVAL_2380;
  assign _EVAL_2835 = _EVAL_3254 == 32'h4;
  assign _EVAL_372 = _EVAL_3254 == 32'h8000001c;
  assign _EVAL_1057 = _EVAL_3254 == 32'h8000004d;
  assign _EVAL_2718 = _EVAL_101 == 12'hb17;
  assign _EVAL_1582 = _EVAL_1511 & _EVAL_231;
  assign _EVAL_1576 = _EVAL_3254 == 32'h80000063;
  assign _EVAL_511 = _EVAL_101 == 12'hc8b;
  assign _EVAL_689 = _EVAL_2930 & _EVAL_1597;
  assign _EVAL_2272 = _EVAL_101 == 12'h336;
  assign _EVAL_2626 = _EVAL_101 == 12'h338;
  assign _EVAL_2426 = _EVAL_2930 & _EVAL_1801;
  assign _EVAL_2390 = _EVAL_101 == 12'hc11;
  assign _EVAL_343 = _EVAL_1511 & _EVAL_2182;
  assign _EVAL_988 = _EVAL_101 == 12'hc09;
  assign _EVAL_2068 = _EVAL_3254 == 32'h8000003c;
  assign _EVAL_516 = _EVAL_3138 | _EVAL_2497;
  assign _EVAL_2417 = _EVAL_101 == 12'hc1a;
  assign _EVAL_2091 = _EVAL_3254 == 32'h80000082;
  assign _EVAL_1072 = _EVAL_3254 == 32'h8000002d;
  assign _EVAL_393 = _EVAL_1718 | _EVAL_538;
  assign _EVAL_3045 = _EVAL_43 & _EVAL_2380;
  assign _EVAL_1511 = _EVAL_98 == 3'h2;
  assign _EVAL_1540 = _EVAL_101 == 12'hb11;
  assign _EVAL_1374 = _EVAL_2930 & _EVAL_1002;
  assign _EVAL_614 = _EVAL_1511 & _EVAL_1260;
  assign _EVAL_1352 = _EVAL_101 == 12'hc89;
  assign _EVAL_517 = _EVAL_2930 & _EVAL_580;
  assign _EVAL_1804 = _EVAL_101 == 12'hc19;
  assign _EVAL_1307 = _EVAL_3254 == 32'h80000062;
  assign _EVAL_533 = _EVAL_2672 | _EVAL_360;
  assign _EVAL_1897 = _EVAL_3254 == 32'h8000003f;
  assign _EVAL_747 = _EVAL_318 & _EVAL_1732;
  assign _EVAL_2526 = _EVAL_101 == 12'h33f;
  assign _EVAL_636 = _EVAL_101 == 12'h3b8;
  assign _EVAL_2925 = _EVAL_2930 & _EVAL_1406;
  assign _EVAL_1373 = _EVAL_49 & _EVAL_889;
  assign _EVAL_2922 = _EVAL_2618 <= 3'h1;
  assign _EVAL_574 = _EVAL_2930 & _EVAL_2935;
  assign _EVAL_1820 = _EVAL_2930 & _EVAL_2675;
  assign _EVAL_1973 = _EVAL_2642 | _EVAL_3071;
  assign _EVAL_755 = _EVAL_101 == 12'hb85;
  assign _EVAL_148 = _EVAL_3254 == 32'h80000085;
  assign _EVAL_2630 = _EVAL_1745 | _EVAL_1076;
  assign _EVAL_2598 = ~_EVAL_2923;
  assign _EVAL_1022 = _EVAL_2930 & _EVAL_994;
  assign _EVAL_1809 = _EVAL_1538 & _EVAL_1414;
  assign _EVAL_2596 = _EVAL_2659 & _EVAL_869;
  assign _EVAL_1981 = _EVAL_2567 & _EVAL_1561;
  assign _EVAL_1623 = _EVAL_3254 == 32'h80000028;
  assign _EVAL_2197 = _EVAL_2370 | _EVAL_1082;
  assign _EVAL_1048 = _EVAL_3220 | _EVAL_1576;
  assign _EVAL_1219 = _EVAL_2930 & _EVAL_238;
  assign _EVAL_3085 = _EVAL_101 == 12'hc06;
  assign _EVAL_1437 = _EVAL_1511 & _EVAL_3222;
  assign _EVAL_1260 = _EVAL_101 == 12'hc8d;
  assign _EVAL_1904 = _EVAL_2930 & _EVAL_1008;
  assign _EVAL_1076 = _EVAL_3254 == 32'h8000002e;
  assign _EVAL_2570 = _EVAL_1681 & _EVAL_3210;
  assign _EVAL_1827 = _EVAL_1511 & _EVAL_1432;
  assign _EVAL_2292 = ~_EVAL_63;
  assign _EVAL_1696 = _EVAL_1511 & _EVAL_426;
  assign _EVAL_496 = _EVAL_2930 & _EVAL_1717;
  assign _EVAL_2675 = _EVAL_101 == 12'h3b5;
  assign _EVAL_3010 = _EVAL_101 == 12'hc0e;
  assign _EVAL_1726 = _EVAL_1511 & _EVAL_3085;
  assign _EVAL_1038 = _EVAL_3254 == 32'h80000020;
  assign _EVAL_1257 = _EVAL_1511 & _EVAL_2565;
  assign _EVAL_2103 = _EVAL_101 == 12'hc1d;
  assign _EVAL_2882 = _EVAL_2074 & _EVAL_1274;
  assign _EVAL_744 = _EVAL_101 == 12'hc1f;
  assign _EVAL_2012 = _EVAL_2930 & _EVAL_1111;
  assign _EVAL_257 = _EVAL_3254 == 32'h80000010;
  assign _EVAL_604 = _EVAL_101 == 12'hc96;
  assign _EVAL_1028 = _EVAL_2930 & _EVAL_792;
  assign _EVAL_2700 = _EVAL_1511 & _EVAL_529;
  assign _EVAL_3004 = _EVAL_3254 == 32'h80000088;
  assign _EVAL_255 = _EVAL_2567 & _EVAL_2112;
  assign _EVAL_2181 = _EVAL_1117 + _EVAL_446;
  assign _EVAL_3192 = _EVAL_1057 | _EVAL_2259;
  assign _EVAL_2025 = _EVAL_2922 | _EVAL_63;
  assign _EVAL_3247 = _EVAL_3254 == 32'h80000040;
  assign _EVAL_990 = _EVAL_658 & _EVAL_2567;
  assign _EVAL_2795 = _EVAL_3254 == 32'h80000071;
  assign _EVAL_1524 = _EVAL_1556 | _EVAL_1826;
  assign _EVAL_2758 = _EVAL_101 == 12'hb91;
  assign _EVAL_2891 = _EVAL_3254 == 32'h80000079;
  assign _EVAL_2600 = _EVAL_101 == 12'h7c1;
  assign _EVAL_1962 = _EVAL_101 == 12'h3be;
  assign _EVAL_3032 = _EVAL_1650 | _EVAL_63;
  assign _EVAL_3003 = _EVAL_2567 & _EVAL_2835;
  assign _EVAL_1358 = _EVAL_101 == 12'hb98;
  assign _EVAL_1572 = _EVAL_3254 == 32'h80000012;
  assign _EVAL_195 = _EVAL_2921 | _EVAL_603;
  assign _EVAL_371 = _EVAL_101 == 12'h3bb;
  assign _EVAL_2855 = _EVAL_393 | _EVAL_3174;
  assign _EVAL_1210 = _EVAL_2930 & _EVAL_2368;
  assign _EVAL_3253 = _EVAL_1511 & _EVAL_3088;
  assign _EVAL_1889 = _EVAL_101 == 12'hc87;
  assign _EVAL_2634 = _EVAL_108 <= _EVAL_1267;
  assign _EVAL_1605 = _EVAL_1511 & _EVAL_1250;
  assign _EVAL_2143 = _EVAL_3146 | _EVAL_527;
  assign _EVAL_1674 = _EVAL_1891 | _EVAL_2612;
  assign _EVAL_1232 = _EVAL_271 | _EVAL_2800;
  assign _EVAL_1733 = _EVAL_3234 | _EVAL_1572;
  assign _EVAL_1262 = _EVAL_2930 & _EVAL_1146;
  assign _EVAL_2522 = _EVAL_101 == 12'hb86;
  assign _EVAL_443 = _EVAL_101 == 12'hc0c;
  assign _EVAL_1025 = _EVAL_101 == 12'h3ba;
  assign _EVAL_1521 = _EVAL_2930 & _EVAL_1059;
  assign _EVAL_2373 = _EVAL_999 | _EVAL_1342;
  assign _EVAL_2099 = _EVAL_1511 & _EVAL_2316;
  assign _EVAL_2266 = _EVAL_1511 & _EVAL_3103;
  assign _EVAL_1449 = _EVAL_2930 & _EVAL_2911;
  assign _EVAL_2957 = _EVAL_101 == 12'hc18;
  assign _EVAL_1363 = _EVAL_318 & _EVAL_2033;
  assign _EVAL_3241 = _EVAL_2634 & _EVAL_42;
  assign _EVAL_2007 = _EVAL_3254 == 32'h80000076;
  assign _EVAL_1046 = _EVAL_783 | _EVAL_1135;
  assign _EVAL_1780 = _EVAL_1511 & _EVAL_2081;
  assign _EVAL_664 = _EVAL_2930 & _EVAL_2758;
  assign _EVAL_529 = _EVAL_101 == 12'hc04;
  assign _EVAL_2785 = _EVAL_3254 == 32'h80000013;
  assign _EVAL_1555 = _EVAL_1511 & _EVAL_511;
  assign _EVAL_2800 = _EVAL_3254 == 32'h80000087;
  assign _EVAL_1237 = _EVAL_2930 & _EVAL_1370;
  assign _EVAL_2807 = _EVAL_1511 & _EVAL_2894;
  assign _EVAL_1431 = _EVAL_101 == 12'h3bc;
  assign _EVAL_638 = _EVAL_533 | _EVAL_1903;
  assign _EVAL_2682 = _EVAL_101 == 12'hb16;
  assign _EVAL_2585 = _EVAL_863 & _EVAL_2567;
  assign _EVAL_248 = _EVAL_2930 & _EVAL_2501;
  assign _EVAL_991 = _EVAL_2930 & _EVAL_579;
  assign _EVAL_2829 = _EVAL_2930 & _EVAL_222;
  assign _EVAL_1902 = _EVAL_2930 & _EVAL_2920;
  assign _EVAL_2997 = _EVAL_1511 & _EVAL_1041;
  assign _EVAL_1254 = _EVAL_2930 & _EVAL_1959;
  assign _EVAL_2560 = _EVAL_1511 & _EVAL_1939;
  assign _EVAL_384 = _EVAL_1222 | _EVAL_352;
  assign _EVAL_2301 = _EVAL_101 == 12'hc14;
  assign _EVAL_2762 = _EVAL_2930 & _EVAL_989;
  assign _EVAL_2961 = _EVAL_101 == 12'hb8f;
  assign _EVAL_643 = _EVAL_1511 & _EVAL_1889;
  assign _EVAL_1008 = _EVAL_101 == 12'hb9f;
  assign _EVAL_2230 = _EVAL_2930 & _EVAL_1619;
  assign _EVAL_3155 = _EVAL_2596 & _EVAL_1610;
  assign _EVAL_695 = _EVAL_101 == 12'hb04;
  assign _EVAL_1622 = _EVAL_101 == 12'h33e;
  assign _EVAL_2240 = _EVAL_2567 & _EVAL_378;
  assign _EVAL_378 = _EVAL_3254 == 32'h8;
  assign _EVAL_1668 = _EVAL_2079 | _EVAL_150;
  assign _EVAL_725 = _EVAL_1659 + _EVAL_93;
  assign _EVAL_225 = _EVAL_3254 == 32'h80000044;
  assign _EVAL_318 = _EVAL_2305 & _EVAL_2454;
  assign _EVAL_1082 = _EVAL_3254 == 32'h80000066;
  assign _EVAL_300 = _EVAL_101 == 12'hb13;
  assign _EVAL_2303 = _EVAL_2826 | _EVAL_1648;
  assign _EVAL_1066 = _EVAL_2570 & _EVAL_1824;
  assign _EVAL_796 = _EVAL_3254 == 32'h80000022;
  assign _EVAL_2683 = _EVAL_1511 & _EVAL_403;
  assign _EVAL_998 = _EVAL_3254 == 32'h8000000b;
  assign _EVAL_307 = _EVAL_2436 | _EVAL_1654;
  assign _EVAL_396 = _EVAL_101 == 12'h33c;
  assign _EVAL_1542 = _EVAL_1511 & _EVAL_604;
  assign _EVAL_246 = _EVAL_2570 & _EVAL_1653;
  assign _EVAL_2556 = _EVAL_2930 & _EVAL_229;
  assign _EVAL_1096 = _EVAL_1615 | _EVAL_2773;
  assign _EVAL_2478 = _EVAL_2930 & _EVAL_465;
  assign _EVAL_1663 = _EVAL_2930 & _EVAL_1431;
  assign _EVAL_1234 = _EVAL_307 | _EVAL_148;
  assign _EVAL_2921 = _EVAL_1836 | _EVAL_1865;
  assign _EVAL_2633 = _EVAL_3254 == 32'h3;
  assign _EVAL_2465 = _EVAL_2403 | _EVAL_3050;
  assign _EVAL_738 = _EVAL_101 == 12'hc1b;
  assign _EVAL_3038 = _EVAL_318 & _EVAL_2778;
  assign _EVAL_349 = _EVAL_1034 | _EVAL_1151;
  assign _EVAL_216 = _EVAL_2930 & _EVAL_2018;
  assign _EVAL_3222 = _EVAL_101 == 12'hc15;
  assign _EVAL_2911 = _EVAL_101 == 12'hb8b;
  assign _EVAL_1565 = _EVAL_3254 == 32'h8000006d;
  assign _EVAL_2930 = _EVAL_595 | _EVAL_2345;
  assign _EVAL_2916 = _EVAL_2930 & _EVAL_3148;
  assign _EVAL_682 = _EVAL_2930 & _EVAL_652;
  assign _EVAL_144 = _EVAL_2596 & _EVAL_889;
  assign _EVAL_3024 = _EVAL_1511 & _EVAL_1840;
  assign _EVAL_185 = _EVAL_1046 | _EVAL_1565;
  assign _EVAL_2214 = _EVAL_1511 & _EVAL_2017;
  assign _EVAL_2897 = _EVAL_1167 | _EVAL_3252;
  assign _EVAL_2132 = _EVAL_1511 & _EVAL_2680;
  assign _EVAL_2973 = _EVAL_2912 & _EVAL_3169;
  assign _EVAL_1342 = _EVAL_3254 == 32'h8000006a;
  assign _EVAL_2120 = _EVAL_750 & _EVAL_2567;
  assign _EVAL_1845 = _EVAL_101 == 12'h325;
  assign _EVAL_355 = _EVAL_2930 & _EVAL_1071;
  assign _EVAL_1538 = _EVAL_2659 & _EVAL_3207;
  assign _EVAL_3212 = _EVAL_101 == 12'h32b;
  assign _EVAL_2436 = _EVAL_687 | _EVAL_1086;
  assign _EVAL_2936 = _EVAL_2930 & _EVAL_3212;
  assign _EVAL_3001 = _EVAL_101 == 12'hb05;
  assign _EVAL_174 = _EVAL_2930 & _EVAL_3188;
  assign _EVAL_1612 = _EVAL_101 == 12'hc84;
  assign _EVAL_579 = _EVAL_101 == 12'hb07;
  assign _EVAL_1745 = _EVAL_2071 | _EVAL_1072;
  assign _EVAL_1145 = _EVAL_101 == 12'hb88;
  assign _EVAL_1461 = _EVAL_2619 | _EVAL_987;
  assign _EVAL_1661 = _EVAL_3254 == 32'h80000037;
  assign _EVAL_165 = _EVAL_1511 & _EVAL_700;
  assign _EVAL_3130 = _EVAL_2930 & _EVAL_555;
  assign _EVAL_2531 = _EVAL_1638 | _EVAL_940;
  assign _EVAL_1923 = _EVAL_2930 & _EVAL_636;
  assign _EVAL_2079 = _EVAL_2967 | _EVAL_2926;
  assign _EVAL_1053 = _EVAL_1822 & _EVAL_2567;
  assign _EVAL_342 = _EVAL_101 == 12'h329;
  assign _EVAL_1574 = _EVAL_1668 | _EVAL_2891;
  assign _EVAL_3244 = _EVAL_2930 & _EVAL_300;
  assign _EVAL_231 = _EVAL_101 == 12'hc8f;
  assign _EVAL_1068 = _EVAL_3254 == 32'h8000001d;
  assign _EVAL_868 = _EVAL_2040 | _EVAL_398;
  assign _EVAL_949 = _EVAL_2074 & _EVAL_2538;
  assign _EVAL_577 = _EVAL_2930 & _EVAL_1168;
  assign _EVAL_538 = _EVAL_3254 == 32'h80000016;
  assign _EVAL_3041 = _EVAL_257 & _EVAL_2567;
  assign _EVAL_3174 = _EVAL_3254 == 32'h80000017;
  assign _EVAL_2497 = _EVAL_3254 == 32'h8000008d;
  assign _EVAL_3107 = _EVAL_3254 == 32'h80000081;
  assign _EVAL_1002 = _EVAL_101 == 12'h339;
  assign _EVAL_2751 = _EVAL_3077 | _EVAL_1870;
  assign _EVAL_2249 = _EVAL_101 == 12'hc99;
  assign _EVAL_458 = _EVAL_541 & _EVAL_2567;
  assign _EVAL_1655 = _EVAL_2930 & _EVAL_2625;
  assign _EVAL_3111 = _EVAL_101 == 12'hc9d;
  assign _EVAL_1067 = _EVAL_2930 & _EVAL_1962;
  assign _EVAL_794 = _EVAL_2930 & _EVAL_3147;
  assign _EVAL_1826 = _EVAL_3254 == 32'h8000001a;
  assign _EVAL_1522 = _EVAL_3254 == 32'h80000047;
  assign _EVAL_1102 = _EVAL_43 & _EVAL_1464;
  assign _EVAL_3220 = _EVAL_858 | _EVAL_1307;
  assign _EVAL_1775 = _EVAL_2930 & _EVAL_1095;
  assign _EVAL_2871 = _EVAL_2930 & _EVAL_359;
  assign _EVAL_587 = _EVAL_2984 & _EVAL_2567;
  assign _EVAL_2499 = _EVAL_1511 & _EVAL_2693;
  assign _EVAL_2207 = _EVAL_3254 == 32'h80000054;
  assign _EVAL_1304 = ~_EVAL;
  assign _EVAL_2238 = _EVAL_1511 & _EVAL_2249;
  assign _EVAL_2601 = _EVAL_2930 & _EVAL_847;
  assign _EVAL_994 = _EVAL_101 == 12'h328;
  assign _EVAL_2726 = _EVAL_2930 & _EVAL_2679;
  assign _EVAL_3141 = _EVAL_2930 & _EVAL_3104;
  assign _EVAL_2935 = _EVAL_101 == 12'hb8c;
  assign _EVAL_2603 = _EVAL_1511 & _EVAL_2301;
  assign _EVAL_2038 = _EVAL_1524 | _EVAL_348;
  assign _EVAL_665 = _EVAL_2930 & _EVAL_1898;
  assign _EVAL_585 = _EVAL_2930 & _EVAL_1294;
  assign _EVAL_2246 = _EVAL_101 == 12'hc9e;
  assign _EVAL_812 = _EVAL_3254 == 32'h8000004c;
  assign _EVAL_1043 = _EVAL_2930 & _EVAL_1253;
  assign _EVAL_1442 = _EVAL_2353 & _EVAL_2567;
  assign _EVAL_1477 = _EVAL_43 & _EVAL_1414;
  assign _EVAL_647 = _EVAL_2197 | _EVAL_697;
  assign _EVAL_2847 = _EVAL_2074 & _EVAL_2706;
  assign _EVAL_2672 = _EVAL_1014 | _EVAL_2242;
  assign _EVAL_2512 = _EVAL_1511 & _EVAL_1804;
  assign _EVAL_888 = _EVAL_3254 == 32'h5;
  assign _EVAL_1855 = _EVAL_101 == 12'hb18;
  assign _EVAL_593 = _EVAL_3254 == 32'h80000069;
  assign _EVAL_2553 = _EVAL_1511 & _EVAL_549;
  assign _EVAL_3200 = _EVAL_3254 == 32'h80000018;
  assign _EVAL_359 = _EVAL_101 == 12'h331;
  assign _EVAL_697 = _EVAL_3254 == 32'h80000067;
  assign _EVAL_687 = _EVAL_1483 | _EVAL_2091;
  assign _EVAL_348 = _EVAL_3254 == 32'h8000001b;
  assign _EVAL_1602 = _EVAL_894 | _EVAL_2027;
  assign _EVAL_2714 = _EVAL_3254 == 32'h80000064;
  assign _EVAL_983 = ~_EVAL_3032;
  assign _EVAL_2439 = _EVAL_3254 == 32'h8000002c;
  assign _EVAL_1840 = _EVAL_101 == 12'hc0a;
  assign _EVAL_2243 = _EVAL_384 | _EVAL_2739;
  assign _EVAL_1648 = _EVAL_3254 == 32'h80000055;
  assign _EVAL_1249 = _EVAL_3254 == 32'h8000005e;
  assign _EVAL_1633 = _EVAL_101 == 12'h32e;
  assign _EVAL_150 = _EVAL_3254 == 32'h80000078;
  assign _EVAL_2183 = _EVAL_1511 & _EVAL_1206;
  assign _EVAL_2353 = _EVAL_1674 | _EVAL_735;
  assign _EVAL_239 = _EVAL_101 == 12'hffc;
  assign _EVAL_295 = _EVAL_1511 & _EVAL_1196;
  assign _EVAL_1921 = _EVAL_1833 | _EVAL_310;
  assign _EVAL_1870 = _EVAL_3254 == 32'h8000005f;
  assign _EVAL_2515 = _EVAL_965 | _EVAL_2883;
  assign _EVAL_1151 = _EVAL_3254 == 32'h8000002a;
  assign _EVAL_1103 = _EVAL_2275 | _EVAL_1160;
  assign _EVAL_2432 = _EVAL_101 == 12'hc97;
  assign _EVAL_921 = _EVAL_3254 == 32'h80000050;
  assign _EVAL_783 = _EVAL_2373 | _EVAL_1943;
  assign _EVAL_2415 = _EVAL_1511 & _EVAL_337;
  assign _EVAL_1496 = _EVAL_2930 & _EVAL_955;
  assign _EVAL_1833 = _EVAL_462 | _EVAL_2456;
  assign _EVAL_240 = _EVAL_2305 & _EVAL_2380;
  assign _EVAL_541 = _EVAL_3254 == 32'h8000008e;
  assign _EVAL_1168 = _EVAL_101 == 12'h3a2;
  assign _EVAL_1111 = _EVAL_101 == 12'hb1a;
  assign _EVAL_2943 = _EVAL_101 == 12'hc8e;
  assign _EVAL_1954 = _EVAL_2930 & _EVAL_1145;
  assign _EVAL_3240 = _EVAL_2839 | _EVAL_545;
  assign _EVAL_147 = _EVAL_101 == 12'h33d;
  assign _EVAL_395 = _EVAL_1139 | _EVAL_2724;
  assign _EVAL_1926 = _EVAL_101 == 12'hb92;
  assign _EVAL_352 = _EVAL_3254 == 32'h80000026;
  assign _EVAL_965 = _EVAL_3094 | _EVAL_2864;
  assign _EVAL_831 = _EVAL_3254 == 32'h80000068;
  assign _EVAL_951 = _EVAL_101 == 12'hb9d;
  assign _EVAL_3126 = _EVAL_2930 & _EVAL_1938;
  assign _EVAL_3146 = _EVAL_2303 | _EVAL_676;
  assign _EVAL_1138 = _EVAL_185 | _EVAL_1426;
  assign _EVAL_3226 = _EVAL_101 == 12'hb8a;
  assign _EVAL_1785 = _EVAL_2930 & _EVAL_2777;
  assign _EVAL_1824 = _EVAL_2634 & _EVAL_2394;
  assign _EVAL_416 = _EVAL_101 == 12'hb1d;
  assign _EVAL_2450 = _EVAL_2798 | _EVAL_1741;
  assign _EVAL_623 = _EVAL_1138 | _EVAL_1161;
  assign _EVAL_3072 = _EVAL_101 == 12'hc88;
  assign _EVAL_1836 = _EVAL_2795 | _EVAL_188;
  assign _EVAL_1903 = _EVAL_3254 == 32'h80000032;
  assign _EVAL_1155 = _EVAL_101 == 12'hb94;
  assign _EVAL_1167 = _EVAL_2337 | _EVAL_2832;
  assign _EVAL_229 = _EVAL_101 == 12'h335;
  assign _EVAL_3190 = _EVAL_3254 == 32'h8000008a;
  assign _EVAL_2033 = _EVAL_1740 & _EVAL_1670;
  assign _EVAL_418 = _EVAL_2930 & _EVAL_2140;
  assign _EVAL_548 = _EVAL_2567 & _EVAL_2633;
  assign _EVAL_1178 = _EVAL_2570 & _EVAL_1966;
  assign _EVAL_1186 = _EVAL_101 == 12'hc0b;
  assign _EVAL_2245 = _EVAL_2930 & _EVAL_3063;
  assign _EVAL_633 = _EVAL_101 == 12'hc91;
  assign _EVAL_3050 = _EVAL_3254 == 32'h80000046;
  assign _EVAL_289 = _EVAL_101 == 12'hb0f;
  assign _EVAL_3061 = _EVAL_101 == 12'h332;
  assign _EVAL_1613 = _EVAL_2659 & _EVAL_93;
  assign _EVAL_3138 = _EVAL_3240 | _EVAL_2520;
  assign _EVAL_1583 = _EVAL_2930 & _EVAL_2272;
  assign _EVAL_188 = _EVAL_3254 == 32'h80000072;
  assign _EVAL_2739 = _EVAL_3254 == 32'h80000027;
  assign _EVAL_2336 = _EVAL_175 | _EVAL_2068;
  assign _EVAL_848 = _EVAL_2783 | _EVAL_2963;
  assign _EVAL_846 = _EVAL_623 | _EVAL_2979;
  assign _EVAL_2812 = _EVAL_1511 & _EVAL_2103;
  assign _EVAL_2316 = _EVAL_101 == 12'hc90;
  assign _EVAL_2864 = _EVAL_3254 == 32'h80000042;
  assign _EVAL_2275 = _EVAL_2136 | _EVAL_2886;
  assign _EVAL_2226 = _EVAL_3254 == 32'h8000005b;
  assign _EVAL_1597 = _EVAL_101 == 12'hb87;
  assign _EVAL_1211 = _EVAL_1511 & _EVAL_1612;
  assign _EVAL_1256 = _EVAL_1511 & _EVAL_3072;
  assign _EVAL_651 = _EVAL_2198 | _EVAL_1828;
  assign _EVAL_1320 = _EVAL_43 & _EVAL_1610;
  assign _EVAL_1253 = _EVAL_101 == 12'h326;
  assign _EVAL_881 = _EVAL_1511 & _EVAL_443;
  assign _EVAL_2566 = _EVAL_1538 & _EVAL_1464;
  assign _EVAL_2018 = _EVAL_101 == 12'h333;
  assign _EVAL_2625 = _EVAL_101 == 12'hb12;
  assign _EVAL_2926 = _EVAL_3254 == 32'h80000077;
  assign _EVAL_1527 = _EVAL_1511 & _EVAL_678;
  assign _EVAL_1708 = _EVAL_846 & _EVAL_2567;
  assign _EVAL_3135 = _EVAL_1511 & _EVAL_1629;
  assign _EVAL_309 = _EVAL_1511 & _EVAL_2943;
  assign _EVAL_1361 = _EVAL_2930 & _EVAL_1540;
  assign _EVAL_434 = _EVAL_3254 == 32'h8000005d;
  assign _EVAL_2910 = _EVAL_1613 & _EVAL_1610;
  assign _EVAL_2055 = _EVAL_1511 & _EVAL_2390;
  assign _EVAL_2883 = _EVAL_3254 == 32'h80000043;
  assign _EVAL_2153 = _EVAL_1538 & _EVAL_889;
  assign _EVAL_1741 = _EVAL_3254 == 32'h8000001f;
  assign _EVAL_958 = _EVAL_2930 & _EVAL_2626;
  assign _EVAL_893 = _EVAL_2930 & _EVAL_985;
  assign _EVAL_3009 = _EVAL_2930 & _EVAL_368;
  assign _EVAL_2140 = _EVAL_101 == 12'hb84;
  assign _EVAL_940 = _EVAL_3254 == 32'h8000007e;
  assign _EVAL_803 = _EVAL_2930 & _EVAL_323;
  assign _EVAL_930 = _EVAL_2930 & _EVAL_2610;
  assign _EVAL_1990 = _EVAL_1511 & _EVAL_744;
  assign _EVAL_709 = _EVAL_101 == 12'hb96;
  assign _EVAL_400 = _EVAL_2038 | _EVAL_372;
  assign _EVAL_1438 = _EVAL_2930 & _EVAL_2684;
  assign _EVAL_1483 = _EVAL_1973 | _EVAL_3107;
  assign _EVAL_1891 = _EVAL_1574 | _EVAL_1285;
  assign _EVAL_1161 = _EVAL_3254 == 32'h8000006f;
  assign _EVAL_2643 = _EVAL_1511 & _EVAL_2957;
  assign _EVAL_2144 = _EVAL_2930 & _EVAL_2639;
  assign _EVAL_2282 = _EVAL_525 & _EVAL_530;
  assign _EVAL_2619 = _EVAL_2450 | _EVAL_1038;
  assign _EVAL_1801 = _EVAL_101 == 12'h334;
  assign _EVAL_1641 = _EVAL_3254 == 32'h80000025;
  assign _EVAL_1629 = _EVAL_101 == 12'hc9a;
  assign _EVAL_1732 = _EVAL_1842 & _EVAL_2706;
  assign _EVAL_1640 = _EVAL_318 & _EVAL_1768;
  assign _EVAL_2080 = _EVAL_1511 & _EVAL_2246;
  assign _EVAL_238 = _EVAL_101 == 12'hb1f;
  assign _EVAL_3252 = _EVAL_3254 == 32'h80000049;
  assign _EVAL_1968 = _EVAL_3254 == 32'h80000033;
  assign _EVAL_1368 = _EVAL_3254 == 32'h1;
  assign _EVAL_939 = _EVAL_3254 == 32'h80000045;
  assign _EVAL_1765 = _EVAL_2930 & _EVAL_1475;
  assign _EVAL_1575 = _EVAL_2855 | _EVAL_3200;
  assign _EVAL_1206 = _EVAL_101 == 12'hc07;
  assign _EVAL_1250 = _EVAL_101 == 12'hc16;
  assign _EVAL_2017 = _EVAL_101 == 12'hc95;
  assign _EVAL_2742 = _EVAL_2930 & _EVAL_2536;
  assign _EVAL_1709 = _EVAL_2930 & _EVAL_942;
  assign _EVAL_268 = _EVAL_2180 & _EVAL_2567;
  assign _EVAL_3094 = _EVAL_3254 == 32'h80000041;
  assign _EVAL_1314 = _EVAL_1625 & _EVAL_2567;
  assign _EVAL_1198 = _EVAL_2082 | _EVAL_2959;
  assign _EVAL_310 = _EVAL_3254 == 32'h80000024;
  assign _EVAL_2242 = _EVAL_3254 == 32'h80000030;
  assign _EVAL_945 = _EVAL_2930 & _EVAL_2763;
  assign _EVAL_1049 = _EVAL_2930 & _EVAL_1536;
  assign _EVAL_2912 = _EVAL_49 & _EVAL_1610;
  assign _EVAL_2886 = _EVAL_3254 == 32'h80000038;
  assign _EVAL_2082 = _EVAL_867 | _EVAL_921;
  assign _EVAL_2371 = _EVAL_3254 == 32'h80000034;
  assign _EVAL_1615 = _EVAL_868 | _EVAL_2226;
  assign _EVAL_2180 = _EVAL_2143 | _EVAL_844;
  assign _EVAL_2220 = _EVAL_1511 & _EVAL_1301;
  assign _EVAL_1535 = _EVAL_1613 & _EVAL_1414;
  assign _EVAL_2874 = _EVAL_949 & _EVAL_1670;
  assign _EVAL_2777 = _EVAL_101 == 12'h3b6;
  assign _EVAL_1670 = _EVAL_108 <= _EVAL_2251;
  assign _EVAL_1456 = _EVAL_2930 & _EVAL_1316;
  assign _EVAL_2885 = _EVAL_108 == 8'h0;
  assign _EVAL_3145 = _EVAL_2930 & _EVAL_951;
  assign _EVAL_2004 = _EVAL_2930 & _EVAL_550;
  assign _EVAL_756 = _EVAL_2930 & _EVAL_1127;
  assign _EVAL_2932 = _EVAL_1687 | _EVAL_1652;
  assign _EVAL_1828 = _EVAL_3254 == 32'h80000014;
  assign _EVAL_2035 = _EVAL_3254 == 32'h8000004a;
  assign _EVAL_942 = _EVAL_101 == 12'hb89;
  assign _EVAL_1406 = _EVAL_101 == 12'hb95;
  assign _EVAL_1285 = _EVAL_3254 == 32'h8000007a;
  assign _EVAL_569 = _EVAL_318 & _EVAL_2847;
  assign _EVAL_3019 = _EVAL_101 == 12'hb10;
  assign _EVAL_1516 = _EVAL_2930 & _EVAL_2526;
  assign _EVAL_1606 = _EVAL_2930 & _EVAL_1278;
  assign _EVAL_2982 = _EVAL_2930 & _EVAL_1633;
  assign _EVAL_2552 = _EVAL_2930 & _EVAL_2002;
  assign _EVAL_2341 = _EVAL_101 == 12'hc93;
  assign _EVAL_2337 = _EVAL_2465 | _EVAL_1522;
  assign _EVAL_2706 = _EVAL_3 < _EVAL_2147;
  assign _EVAL_1536 = _EVAL_101 == 12'hb19;
  assign _EVAL_2780 = _EVAL_101 == 12'hb97;
  assign _EVAL_2773 = _EVAL_3254 == 32'h8000005c;
  assign _EVAL_2924 = _EVAL_1511 & _EVAL_1352;
  assign _EVAL_1196 = _EVAL_101 == 12'hc9b;
  assign _EVAL_1625 = _EVAL_3254 == 32'h80000003;
  assign _EVAL_2010 = _EVAL_1538 & _EVAL_1610;
  assign _EVAL_1003 = _EVAL_2930 & _EVAL_1402;
  assign _EVAL_1370 = _EVAL_101 == 12'hb08;
  assign _EVAL_1005 = _EVAL_1511 & _EVAL_2491;
  assign _EVAL_2399 = _EVAL_2930 & _EVAL_1622;
  assign _EVAL_760 = _EVAL_2930 & _EVAL_416;
  assign _EVAL_527 = _EVAL_3254 == 32'h80000057;
  assign _EVAL_1147 = _EVAL_2930 & _EVAL_2555;
  assign _EVAL_3223 = _EVAL_2244 | _EVAL_2371;
  assign _EVAL_2664 = _EVAL_3254 == 32'h8000002f;
  assign _EVAL_1109 = _EVAL_3254 == 32'h80000015;
  assign _EVAL_1430 = _EVAL_2930 & _EVAL_1807;
  assign _EVAL_465 = _EVAL_101 == 12'hb0a;
  assign _EVAL_530 = ~_EVAL_59;
  assign _EVAL_1170 = _EVAL_1511 & _EVAL_738;
  assign _EVAL_321 = _EVAL_1511 & _EVAL_3010;
  assign _EVAL_2259 = _EVAL_3254 == 32'h8000004e;
  assign _EVAL_2612 = _EVAL_3254 == 32'h8000007b;
  assign _EVAL_1959 = _EVAL_101 == 12'hb90;
  assign _EVAL_1748 = _EVAL_998 & _EVAL_2567;
  assign _EVAL_426 = _EVAL_101 == 12'hc98;
  assign _EVAL_2174 = _EVAL_1511 & _EVAL_2052;
  assign _EVAL_3221 = _EVAL_1511 & _EVAL_1242;
  assign _EVAL_1481 = _EVAL_2930 & _EVAL_2600;
  assign _EVAL_1786 = _EVAL_1613 & _EVAL_889;
  assign _EVAL_1059 = _EVAL_101 == 12'h32f;
  assign _EVAL_1471 = _EVAL_2912 & _EVAL_433;
  assign _EVAL_603 = _EVAL_3254 == 32'h80000074;
  assign _EVAL_450 = _EVAL_2596 & _EVAL_1464;
  assign _EVAL_3232 = _EVAL_1511 & _EVAL_1186;
  assign _EVAL_2368 = _EVAL_101 == 12'hb9a;
  assign _EVAL_792 = _EVAL_101 == 12'h32c;
  assign _EVAL_2024 = _EVAL_2930 & _EVAL_289;
  assign _EVAL_1718 = _EVAL_651 | _EVAL_1109;
  assign _EVAL_2768 = _EVAL_1511 & _EVAL_988;
  assign _EVAL_955 = _EVAL_101 == 12'h3bf;
  assign _EVAL_2832 = _EVAL_3254 == 32'h80000048;
  assign _EVAL_1426 = _EVAL_3254 == 32'h8000006e;
  assign _EVAL_2377 = _EVAL_2930 & _EVAL_2961;
  assign _EVAL_1140 = _EVAL_3254 == 32'h6;
  assign _EVAL_3104 = _EVAL_101 == 12'h3a1;
  assign _EVAL_2078 = _EVAL_1096 | _EVAL_434;
  assign _EVAL_1867 = _EVAL_3254 == 32'h8000003b;
  assign _EVAL_2254 = _EVAL_1373 & _EVAL_433;
  assign _EVAL_3092 = _EVAL_1511 & _EVAL_2127;
  assign _EVAL_1650 = _EVAL_889 | _EVAL_1610;
  assign _EVAL_2610 = _EVAL_101 == 12'hb15;
  assign _EVAL_1160 = _EVAL_3254 == 32'h80000039;
  assign _EVAL_1180 = _EVAL_2930 & _EVAL_816;
  assign _EVAL_1188 = _EVAL_2930 & _EVAL_528;
  assign _EVAL_999 = _EVAL_2892 | _EVAL_593;
  assign _EVAL_1638 = _EVAL_3254 == 32'h8000007d;
  assign _EVAL_549 = _EVAL_101 == 12'hc92;
  assign _EVAL_398 = _EVAL_3254 == 32'h8000005a;
  assign _EVAL_3238 = _EVAL_1373 & _EVAL_827;
  assign _EVAL_929 = _EVAL_2930 & _EVAL_342;
  assign _EVAL_2555 = _EVAL_101 == 12'h3a3;
  assign _EVAL_823 = _EVAL_2930 & _EVAL_2522;
  assign _EVAL_360 = _EVAL_3254 == 32'h80000031;
  assign _EVAL_2027 = _EVAL_3254 == 32'h80000089;
  assign _EVAL_1653 = _EVAL_1771 & _EVAL_42;
  assign _EVAL_3103 = _EVAL_101 == 12'hc85;
  assign _EVAL_863 = _EVAL_1754 | _EVAL_3247;
  assign _EVAL_3118 = _EVAL_1511 & _EVAL_1445;
  assign _EVAL_1284 = _EVAL_349 | _EVAL_696;
  assign _EVAL_827 = _EVAL_1 > _EVAL_129;
  assign _EVAL_1703 = _EVAL_101 == 12'h324;
  assign _EVAL_2547 = _EVAL_2930 & _EVAL_3019;
  assign _EVAL_1784 = _EVAL_1511 & _EVAL_3111;
  assign _EVAL_1086 = _EVAL_3254 == 32'h80000083;
  assign _EVAL_2969 = _EVAL_3254 == 32'h80000053;
  assign _EVAL_1747 = _EVAL_101 == 12'h33b;
  assign _EVAL_2797 = _EVAL_2930 & _EVAL_1878;
  assign _EVAL_1402 = _EVAL_101 == 12'h3b7;
  assign _EVAL_900 = _EVAL_1511 & _EVAL_2852;
  assign _EVAL_2756 = _EVAL_2567 & _EVAL_888;
  assign _EVAL_2137 = _EVAL_154 & _EVAL_2567;
  assign _EVAL_844 = _EVAL_3254 == 32'h80000058;
  assign _EVAL_1769 = _EVAL_2930 & _EVAL_789;
  assign _EVAL_3077 = _EVAL_2078 | _EVAL_1249;
  assign _EVAL_2198 = _EVAL_1733 | _EVAL_2785;
  assign _EVAL_867 = _EVAL_3192 | _EVAL_3108;
  assign _EVAL_992 = _EVAL_2930 & _EVAL_3185;
  assign _EVAL_2283 = _EVAL_2746 & _EVAL_3207;
  assign _EVAL_1242 = _EVAL_101 == 12'hc8a;
  assign _EVAL_2852 = _EVAL_101 == 12'hc05;
  assign _EVAL_2473 = _EVAL_2930 & _EVAL_755;
  assign _EVAL_166 = _EVAL_2930 & _EVAL_984;
  assign _EVAL_2693 = _EVAL_101 == 12'hc94;
  always @(posedge _EVAL_16) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1606 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4cd9f6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eeb48d1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1188 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(123e07fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6636f64b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3155 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fa1c5ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1227 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91a3e215)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1516 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca1357ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1028 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f8d4168)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2560 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(933f12b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_418 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9523bf50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2952 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50612f69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1663 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2aa9df26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2596 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a5ec829)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1923 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68125add)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_425 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da687d45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3130 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c971200)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2245 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87c722b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2036 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fb4fee7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2556 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fce93f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1003 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a627c871)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1066 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0dff74a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3003 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34d2532c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3024 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3bcdc2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2137 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ee5da53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1605 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(348d4b99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2552 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50cd5526)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1257 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3316d92f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3118 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33a29cdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_324 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0486f05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2797 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5dc95029)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2820 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f867649)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1053 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7febae35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2238 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(771adde5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1542 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dba4669)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_343 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d125dfc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2982 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c174c2ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2742 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9a90e14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_837 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc30d2f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1443 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4042c04f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1481 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf46c47a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_664 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8686f2e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3154 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8717df8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_758 & _EVAL_983) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1655 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(239e619e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1254 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d06c80ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_517 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6261ed33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc0b075f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2329 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d442a89d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2066 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53210bc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3009 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2bbe0af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2598) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(480d6a97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2871 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32527930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1521 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eae57084)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_575 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f89d2a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_945 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2866821d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2339 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e46b4577)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_574 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec53bc1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1582 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be134a74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2230 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6d545fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1430 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a15c067)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2473 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(205c4601)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1067 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94cebba6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2603 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df9a07f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3250e9a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1712 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14283b37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2220 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(889e5216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_760 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72e665c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1373 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4590f2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3041 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88e4c30d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_577 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc62b4d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1180 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(652f1905)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1785 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d40d584b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1640 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba64184f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1696 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be52dc0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_931 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9422ade)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1256 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9eee867)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1437 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b80a060)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1210 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b7acb19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2726 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(966899da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1728 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d3c132)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2153 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99223b74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1314 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(516a611b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3221 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1501690b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_842 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(680dcb53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a8b0c92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2601 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f688333)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3023 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dcab60ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2643 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2acb4f82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1147 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7980aae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3145 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aee62e81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1496 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e288faa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1341 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fda8a525)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1874 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fa10550)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1414 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d121a1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2916 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24d4c095)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6875099)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3038 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bbcbc6bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_389 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86b520eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1346 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c125135)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_518 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e0029ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2080 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec73625e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_757 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(611e8ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2503 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1144761)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_990 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebb19096)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2266 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37e781d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1022 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e13824b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_803 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef9b8dfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_585 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b563ff31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3092 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7733a25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2116 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28028cbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2997 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f819c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2240 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d94a6930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1438 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76762689)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1784 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b86c5cd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_794 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab48b48c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1504 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2773dda8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2768 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(689b4796)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1363 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99949532)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1610 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66a94c24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1748 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e33e2c9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3028 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cfa1616)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2214 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c6cc9df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1765 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ca37106)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_747 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13b4d1a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1527 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7160774a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_893 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28268785)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1102 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fea4893f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2476 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e066bd0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1498 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2adf84f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1442 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3185e846)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1786 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(499e0990)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcbe0471)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2377 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f92e7192)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1726 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa9bbade)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2512 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff39447c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2399 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(428dde92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3244 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62ff2d3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebcc0269)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5dd10f3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2700 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(404081ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1361 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c69da2f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_900 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12f73d80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1456 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48271ce3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_758 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f76cc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_355 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91e0f00f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1211 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(914c5ed1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3126 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(805e67bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1477 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74b4225c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_930 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1854f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2282 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad84efec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38d40446)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1809 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5405c5a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1820 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0e0c498)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1810) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_889 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a07770c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1170 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75dc2b16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2055 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb0f1e3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2829 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d8829b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1827 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(473caf73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1084 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c09c75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3232 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5056e45b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cabd20fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2995 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35bb4588)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_665 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57ac47a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1449 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a271e21b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2120 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a18b0a77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_392 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43080b53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3141 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e588dc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1509 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b8eadaa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2547 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72730911)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3253 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7dbc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2924 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acb76751)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1708 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bb4e77b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2024 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50427b79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2910 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16da371)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1219 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94e0cdf5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_496 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2e16d69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_592 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(168a09d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2973 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40fc3f8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1981 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(946c1804)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1990 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d636f2c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2756 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7eb56a1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_881 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ede100b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3238 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(966de3e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3135 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30d03e1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2183 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(380f976d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2623 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17c8da49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2499 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20f1a19c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bf4459)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1810) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62ee322c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2305 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f02dfc14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2762 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ddd45f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3045 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(969ab45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1345 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3eda91c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1613 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7609c8a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1237 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3da94af7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2885 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc05f140)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1779 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27656e24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1471 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4ba153c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2365 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(427ca843)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1374 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a5ed0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_455 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf95be2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1100 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93cd9711)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1904 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dcaca933)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1043 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5bcd95d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2132 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bff4187)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_929 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b780bdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1598 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad8964e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2566 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7202a9e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3083 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a109477)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_992 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b98d3f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1178 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2914560f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1775 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3e716fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2187 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ee40578)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_548 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9919068)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_958 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23f92c57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_838 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38ee122e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1769 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22f3fe61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_569 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92e17e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2099 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fd6d5ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_682 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa71585b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1954 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83633c86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2925 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26e8f639)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2415 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(656aa95b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1320 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8152ae18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2254 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16dc5ee2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2553 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2be6a072)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_756 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a3b43f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_614 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51d26df4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2782 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(380449ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1378 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4defe9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2426 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f0ef4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1583 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d18a0558)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_839 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff6bf50f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2176 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(568b6a9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2812 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6edf7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2012 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d72a34e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1780 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bee83ca8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1049 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(883e332a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1570 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c423c69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2004 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44bb12fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1902 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d94c490c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2683 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f7793e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1645 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(775b45e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1535 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdf00a42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2598) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2478 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31a8d0e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2749 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff991fba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9302185f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1709 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(464283a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_758 & _EVAL_983) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7130518c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1434 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(437ddcb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2144 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55f9b75d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1262 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(699425d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_689 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33c5dab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2585 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7394006f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1950 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55678743)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1464 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(770ebdf1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_488 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a68e0660)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1555 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ce99ec7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_991 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e517579)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbda3825)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1005 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dde968ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2807 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a091fdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2936 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59be3cce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2174 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e24ac76a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7029b88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_450 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a10dd0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_823 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea3c78ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_536 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49489d97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1b61b71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1182 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3b7256d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_797 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32ca6995)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1336 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4468c086)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1667 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87c587df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_458 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc8a629c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1091 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb2e0539)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_464 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbdf0478)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2010 & _EVAL_2292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae700054)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
