//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_80_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [1:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [11:0] _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input  [3:0]  _EVAL_12,
  input  [1:0]  _EVAL_13,
  input         _EVAL_14
);
  wire [1:0] _EVAL_15;
  wire [4:0] _EVAL_16;
  wire [4:0] _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire [1:0] _EVAL_24;
  reg [4:0] _EVAL_25;
  reg [31:0] _RAND_0;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire [4:0] _EVAL_28;
  reg  _EVAL_30;
  reg [31:0] _RAND_1;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire [1:0] _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire [7:0] _EVAL_44;
  reg [2:0] _EVAL_45;
  reg [31:0] _RAND_2;
  wire [4:0] _EVAL_46;
  wire [1:0] _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire [1:0] _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire [3:0] _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire [1:0] _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire [4:0] _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire [1:0] _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire [31:0] _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire [12:0] _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire [4:0] _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_107;
  wire [11:0] _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire [4:0] _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  reg [1:0] _EVAL_123;
  reg [31:0] _RAND_3;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire [1:0] _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  reg [1:0] _EVAL_136;
  reg [31:0] _RAND_4;
  wire [4:0] _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  reg [2:0] _EVAL_141;
  reg [31:0] _RAND_5;
  wire  _EVAL_142;
  wire  _EVAL_143;
  reg  _EVAL_144;
  reg [31:0] _RAND_6;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  reg [2:0] _EVAL_151;
  reg [31:0] _RAND_7;
  wire  _EVAL_152;
  reg [31:0] _EVAL_153;
  reg [31:0] _RAND_8;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire [1:0] _EVAL_160;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire [12:0] _EVAL_165;
  wire [1:0] _EVAL_166;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire [3:0] _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [32:0] _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire [7:0] _EVAL_184;
  wire [7:0] _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  reg [11:0] _EVAL_190;
  reg [31:0] _RAND_9;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire [7:0] _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  reg [2:0] _EVAL_209;
  reg [31:0] _RAND_10;
  wire [4:0] _EVAL_210;
  wire  _EVAL_211;
  reg  _EVAL_212;
  reg [31:0] _RAND_11;
  wire  _EVAL_213;
  wire [12:0] _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire [3:0] _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire [3:0] _EVAL_229;
  wire [11:0] _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  reg  _EVAL_234;
  reg [31:0] _RAND_12;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  reg [2:0] _EVAL_238;
  reg [31:0] _RAND_13;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_80 = _EVAL_8 & _EVAL_158;
  assign _EVAL_55 = _EVAL_10 == 3'h4;
  assign _EVAL_21 = ~_EVAL_130;
  assign _EVAL_178 = ~_EVAL_7;
  assign _EVAL_146 = _EVAL_2 & _EVAL_67;
  assign _EVAL_166 = _EVAL_0[2:1];
  assign _EVAL_47 = _EVAL_30 - 1'h1;
  assign _EVAL_51 = _EVAL_191 | _EVAL_1;
  assign _EVAL_237 = _EVAL_8 & _EVAL_82;
  assign _EVAL_244 = _EVAL_10 == _EVAL_45;
  assign _EVAL_213 = ~_EVAL_50;
  assign _EVAL_217 = _EVAL_27 | _EVAL_97;
  assign _EVAL_99 = _EVAL_47[0];
  assign _EVAL_69 = _EVAL_10[2:1];
  assign _EVAL_66 = _EVAL_145 | _EVAL_1;
  assign _EVAL_182 = _EVAL_162 | _EVAL_122;
  assign _EVAL_220 = _EVAL_6 == 3'h2;
  assign _EVAL_82 = _EVAL_6 == 3'h4;
  assign _EVAL_137 = 5'h3 << _EVAL_13;
  assign _EVAL_208 = _EVAL_13[0];
  assign _EVAL_132 = ~_EVAL_207;
  assign _EVAL_112 = _EVAL_110 | _EVAL_1;
  assign _EVAL_154 = _EVAL_6 == 3'h0;
  assign _EVAL_197 = _EVAL_2 & _EVAL_114;
  assign _EVAL_147 = _EVAL & _EVAL_2;
  assign _EVAL_119 = _EVAL_13 >= 2'h2;
  assign _EVAL_111 = _EVAL_5 == _EVAL_141;
  assign _EVAL_131 = _EVAL_41[0];
  assign _EVAL_172 = _EVAL_8 & _EVAL_117;
  assign _EVAL_164 = _EVAL_229 == 4'h0;
  assign _EVAL_184 = _EVAL_58 ? _EVAL_205 : 8'h0;
  assign _EVAL_189 = _EVAL_155 & _EVAL_140;
  assign _EVAL_149 = ~_EVAL_170;
  assign _EVAL_165 = _EVAL_214;
  assign _EVAL_188 = _EVAL_204 & _EVAL_140;
  assign _EVAL_58 = _EVAL_240 & _EVAL_77;
  assign _EVAL_54 = _EVAL_5 <= 3'h1;
  assign _EVAL_59 = ~_EVAL_88;
  assign _EVAL_155 = _EVAL_9[1];
  assign _EVAL_94 = _EVAL_175 | _EVAL_169;
  assign _EVAL_191 = _EVAL_40 & _EVAL_36;
  assign _EVAL_70 = _EVAL_224 == 4'h0;
  assign _EVAL_230 = _EVAL_9 & _EVAL_108;
  assign _EVAL_138 = _EVAL_3 == _EVAL_151;
  assign _EVAL_125 = _EVAL_4 >= 2'h2;
  assign _EVAL_120 = _EVAL_204 & _EVAL_95;
  assign _EVAL_193 = _EVAL_201 | _EVAL_1;
  assign _EVAL_240 = _EVAL_14 & _EVAL_8;
  assign _EVAL_86 = _EVAL_73 | _EVAL_1;
  assign _EVAL_196 = _EVAL_41[1];
  assign _EVAL_104 = _EVAL_76 | _EVAL_25;
  assign _EVAL_113 = _EVAL_5 != 3'h0;
  assign _EVAL_207 = _EVAL_63 | _EVAL_1;
  assign _EVAL_133 = _EVAL_54 | _EVAL_1;
  assign _EVAL_20 = _EVAL_3 == 3'h2;
  assign _EVAL_176 = ~_EVAL_53;
  assign _EVAL_96 = _EVAL_119 | _EVAL_232;
  assign _EVAL_68 = ~_EVAL_102;
  assign _EVAL_148 = _EVAL_131 & _EVAL_242;
  assign _EVAL_22 = ~_EVAL_37;
  assign _EVAL_241 = ~_EVAL_212;
  assign _EVAL_79 = _EVAL_121 | _EVAL_1;
  assign _EVAL_171 = ~_EVAL_65;
  assign _EVAL_187 = _EVAL_8 & _EVAL_154;
  assign _EVAL_17 = _EVAL_25 | _EVAL_76;
  assign _EVAL_152 = ~_EVAL_56;
  assign _EVAL_173 = _EVAL_4 == _EVAL_123;
  assign _EVAL_215 = ~_EVAL_129;
  assign _EVAL_62 = _EVAL_131 & _EVAL_189;
  assign _EVAL_60 = ~_EVAL_32;
  assign _EVAL_126 = _EVAL_2 & _EVAL_26;
  assign _EVAL_49 = ~_EVAL_198;
  assign _EVAL_211 = _EVAL_96 | _EVAL_148;
  assign _EVAL_35 = _EVAL_5 <= 3'h4;
  assign _EVAL_53 = _EVAL_202 | _EVAL_1;
  assign _EVAL_200 = _EVAL_164 | _EVAL_1;
  assign _EVAL_124 = ~_EVAL_79;
  assign _EVAL_194 = ~_EVAL_86;
  assign _EVAL_169 = _EVAL_69 == 2'h0;
  assign _EVAL_31 = ~_EVAL_133;
  assign _EVAL_150 = _EVAL_96 | _EVAL_62;
  assign _EVAL_231 = _EVAL_35 | _EVAL_1;
  assign _EVAL_109 = _EVAL_138 | _EVAL_1;
  assign _EVAL_33 = _EVAL_240 & _EVAL_241;
  assign _EVAL_203 = _EVAL_25 != 5'h0;
  assign _EVAL_40 = _EVAL_13 <= 2'h2;
  assign _EVAL_206 = _EVAL_8 & _EVAL_181;
  assign _EVAL_163 = ~_EVAL_219;
  assign _EVAL_236 = _EVAL_244 | _EVAL_1;
  assign _EVAL_36 = $signed(_EVAL_165) == 13'sh0;
  assign _EVAL_227 = ~_EVAL_1;
  assign _EVAL_76 = _EVAL_184[4:0];
  assign _EVAL_46 = _EVAL_17 & _EVAL_28;
  assign _EVAL_201 = _EVAL_5 <= 3'h2;
  assign _EVAL_183 = _EVAL_0 == _EVAL_238;
  assign _EVAL_221 = _EVAL_15[0];
  assign _EVAL_140 = ~_EVAL_95;
  assign _EVAL_48 = _EVAL_3 <= 3'h6;
  assign _EVAL_175 = _EVAL_69 == 2'h1;
  assign _EVAL_170 = _EVAL_49 | _EVAL_1;
  assign _EVAL_110 = _EVAL_94 | _EVAL_55;
  assign _EVAL_139 = ~_EVAL_231;
  assign _EVAL_219 = _EVAL_103 | _EVAL_1;
  assign _EVAL_101 = _EVAL_8 & _EVAL_177;
  assign _EVAL_199 = _EVAL_8 & _EVAL_220;
  assign _EVAL_179 = _EVAL_70 | _EVAL_1;
  assign _EVAL_23 = _EVAL_2 & _EVAL_243;
  assign _EVAL_214 = $signed(_EVAL_100) & -13'sh1000;
  assign _EVAL_103 = _EVAL_182 | _EVAL_135;
  assign _EVAL_115 = _EVAL_44[4:0];
  assign _EVAL_162 = _EVAL_166 == 2'h1;
  assign _EVAL_105 = ~_EVAL_51;
  assign _EVAL_229 = ~_EVAL_12;
  assign _EVAL_180 = _EVAL_3 == 3'h1;
  assign _EVAL_160 = 2'h1 << _EVAL_208;
  assign _EVAL_157 = ~_EVAL_114;
  assign _EVAL_243 = _EVAL_3 == 3'h0;
  assign _EVAL_98 = _EVAL_217 | _EVAL_18;
  assign _EVAL_142 = _EVAL_64 | _EVAL_1;
  assign _EVAL_42 = ~_EVAL_179;
  assign _EVAL_121 = _EVAL_12 == _EVAL_65;
  assign _EVAL_37 = _EVAL_239 | _EVAL_1;
  assign _EVAL_73 = _EVAL_9 == _EVAL_190;
  assign _EVAL_83 = _EVAL_131 & _EVAL_120;
  assign _EVAL_87 = ~_EVAL_144;
  assign _EVAL_242 = _EVAL_155 & _EVAL_95;
  assign _EVAL_74 = _EVAL_240 | _EVAL_147;
  assign _EVAL_168 = _EVAL_2 & _EVAL_159;
  assign _EVAL_181 = _EVAL_6 == 3'h1;
  assign _EVAL_28 = ~_EVAL_115;
  assign _EVAL_92 = _EVAL_196 & _EVAL_204;
  assign _EVAL_156 = ~_EVAL_193;
  assign _EVAL_210 = _EVAL_104 >> _EVAL_10;
  assign _EVAL_91 = ~_EVAL_142;
  assign _EVAL_93 = _EVAL_174[31:0];
  assign _EVAL_177 = _EVAL_6 == 3'h7;
  assign _EVAL_85 = _EVAL_98 | _EVAL_1;
  assign _EVAL_134 = ~_EVAL_241;
  assign _EVAL_185 = 8'h1 << _EVAL_10;
  assign _EVAL_27 = ~_EVAL_203;
  assign _EVAL_116 = ~_EVAL_112;
  assign _EVAL_41 = _EVAL_160 | 2'h1;
  assign _EVAL_130 = _EVAL_125 | _EVAL_1;
  assign _EVAL_88 = _EVAL_137[1:0];
  assign _EVAL_233 = ~_EVAL_234;
  assign _EVAL_75 = _EVAL_173 | _EVAL_1;
  assign _EVAL_84 = _EVAL_178 | _EVAL_1;
  assign _EVAL_159 = ~_EVAL_233;
  assign _EVAL_117 = _EVAL_6 == 3'h5;
  assign _EVAL_64 = _EVAL_6 == _EVAL_209;
  assign _EVAL_222 = ~_EVAL_200;
  assign _EVAL_34 = _EVAL_6 == 3'h3;
  assign _EVAL_129 = _EVAL_119 | _EVAL_1;
  assign _EVAL_135 = _EVAL_0 == 3'h4;
  assign _EVAL_145 = _EVAL_5 == 3'h0;
  assign _EVAL_122 = _EVAL_166 == 2'h0;
  assign _EVAL_15 = _EVAL_144 - 1'h1;
  assign _EVAL_106 = _EVAL_48 | _EVAL_1;
  assign _EVAL_228 = _EVAL_147 & _EVAL_233;
  assign _EVAL_26 = _EVAL_3 == 3'h5;
  assign _EVAL_97 = plusarg_reader_out == 32'h0;
  assign _EVAL_107 = _EVAL_13 == _EVAL_136;
  assign _EVAL_95 = _EVAL_9[0];
  assign _EVAL_224 = _EVAL_12 & _EVAL_171;
  assign _EVAL_24 = _EVAL_234 - 1'h1;
  assign _EVAL_114 = _EVAL_3 == 3'h6;
  assign _EVAL_71 = _EVAL_128 | _EVAL_216;
  assign _EVAL_50 = _EVAL_183 | _EVAL_1;
  assign _EVAL_143 = _EVAL_57 & _EVAL_157;
  assign _EVAL_202 = _EVAL_5 <= 3'h3;
  assign _EVAL_52 = _EVAL_128 | _EVAL_83;
  assign _EVAL_43 = _EVAL_2 & _EVAL_180;
  assign _EVAL_77 = ~_EVAL_30;
  assign _EVAL_57 = _EVAL_147 & _EVAL_87;
  assign _EVAL_235 = _EVAL_8 & _EVAL_34;
  assign _EVAL_174 = _EVAL_153 + 32'h1;
  assign _EVAL_63 = _EVAL_230 == 12'h0;
  assign _EVAL_158 = _EVAL_6 == 3'h6;
  assign _EVAL_118 = ~_EVAL_75;
  assign _EVAL_216 = _EVAL_131 & _EVAL_188;
  assign _EVAL_198 = _EVAL_16[0];
  assign _EVAL_225 = _EVAL_24[0];
  assign _EVAL_108 = {{10'd0}, _EVAL_59};
  assign _EVAL_232 = _EVAL_196 & _EVAL_155;
  assign _EVAL_65 = {_EVAL_211,_EVAL_150,_EVAL_52,_EVAL_71};
  assign _EVAL_192 = ~_EVAL_109;
  assign _EVAL_100 = {1'b0,$signed(_EVAL_9)};
  assign _EVAL_89 = _EVAL_2 & _EVAL_20;
  assign _EVAL_19 = ~_EVAL_85;
  assign _EVAL_67 = _EVAL_3 == 3'h4;
  assign _EVAL_195 = ~_EVAL_84;
  assign _EVAL_102 = _EVAL_111 | _EVAL_1;
  assign _EVAL_32 = _EVAL_107 | _EVAL_1;
  assign _EVAL_223 = ~_EVAL_106;
  assign _EVAL_56 = _EVAL_113 | _EVAL_1;
  assign _EVAL_44 = _EVAL_143 ? _EVAL_185 : 8'h0;
  assign _EVAL_226 = _EVAL_8 & _EVAL_134;
  assign _EVAL_128 = _EVAL_119 | _EVAL_92;
  assign _EVAL_204 = ~_EVAL_155;
  assign _EVAL_205 = 8'h1 << _EVAL_0;
  assign _EVAL_218 = _EVAL_127[0];
  assign _EVAL_127 = _EVAL_212 - 1'h1;
  assign _EVAL_18 = _EVAL_153 < plusarg_reader_out;
  assign _EVAL_186 = ~_EVAL_66;
  assign _EVAL_39 = ~_EVAL_236;
  assign _EVAL_239 = _EVAL_210[0];
  assign _EVAL_16 = _EVAL_25 >> _EVAL_0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_25 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_30 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_45 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_123 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_136 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_141 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_144 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_151 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_153 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_190 = _RAND_9[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_209 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_212 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_234 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_238 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_11) begin
    if (_EVAL_1) begin
      _EVAL_25 <= 5'h0;
    end else begin
      _EVAL_25 <= _EVAL_46;
    end
    if (_EVAL_1) begin
      _EVAL_30 <= 1'h0;
    end else if (_EVAL_240) begin
      if (_EVAL_77) begin
        _EVAL_30 <= 1'h0;
      end else begin
        _EVAL_30 <= _EVAL_99;
      end
    end
    if (_EVAL_228) begin
      _EVAL_45 <= _EVAL_10;
    end
    if (_EVAL_228) begin
      _EVAL_123 <= _EVAL_4;
    end
    if (_EVAL_33) begin
      _EVAL_136 <= _EVAL_13;
    end
    if (_EVAL_33) begin
      _EVAL_141 <= _EVAL_5;
    end
    if (_EVAL_1) begin
      _EVAL_144 <= 1'h0;
    end else if (_EVAL_147) begin
      if (_EVAL_87) begin
        _EVAL_144 <= 1'h0;
      end else begin
        _EVAL_144 <= _EVAL_221;
      end
    end
    if (_EVAL_228) begin
      _EVAL_151 <= _EVAL_3;
    end
    if (_EVAL_1) begin
      _EVAL_153 <= 32'h0;
    end else if (_EVAL_74) begin
      _EVAL_153 <= 32'h0;
    end else begin
      _EVAL_153 <= _EVAL_93;
    end
    if (_EVAL_33) begin
      _EVAL_190 <= _EVAL_9;
    end
    if (_EVAL_33) begin
      _EVAL_209 <= _EVAL_6;
    end
    if (_EVAL_1) begin
      _EVAL_212 <= 1'h0;
    end else if (_EVAL_240) begin
      if (_EVAL_241) begin
        _EVAL_212 <= 1'h0;
      end else begin
        _EVAL_212 <= _EVAL_218;
      end
    end
    if (_EVAL_1) begin
      _EVAL_234 <= 1'h0;
    end else if (_EVAL_147) begin
      if (_EVAL_233) begin
        _EVAL_234 <= 1'h0;
      end else begin
        _EVAL_234 <= _EVAL_225;
      end
    end
    if (_EVAL_33) begin
      _EVAL_238 <= _EVAL_0;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87e8197d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ba8f164)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_31) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2b609d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5dbcf504)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fdb73eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85ba0774)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2aa40293)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4304c3d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7f130b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac32d959)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab477b73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b336102)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8186b77f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(315a9271)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(345da65b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24d31e43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23a4b902)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33b8daee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87f165b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(758788b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9fffef8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21691188)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ab8c23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6854a34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_31) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6db65ac3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d5ecbae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67a0fa0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb218809)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83afe4f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(838b80c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14d093b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e3bb302)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1c87887)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aca1aa18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aab4e071)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(242b7670)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77bd5b57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63e0385f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51fddbd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ab440c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fb75324)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d72d997)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e056997a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f0dbb67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f7f0c8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e938e52d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37f2582e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e6d67b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec903ad9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef2eb349)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3fff6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c8c0cbe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec33a0ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d25796a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4341c6eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f574cde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b561d557)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fab0bdfd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ed8a9bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(659e3aff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87fc8607)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ee3279d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77293d95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb0ee467)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(756e7d97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3afb4e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7edfa8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(299a6283)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(287bbdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2d59905)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bfcd8e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5d67933)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
