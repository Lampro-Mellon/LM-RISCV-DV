//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_2_assert(
  input  [3:0]  _EVAL,
  input  [3:0]  _EVAL_0,
  input  [31:0] _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [3:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [1:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16,
  input  [2:0]  _EVAL_17,
  input         _EVAL_18
);
  wire  _EVAL_19;
  wire [6:0] _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire [32:0] _EVAL_30;
  reg [5:0] _EVAL_31;
  reg [31:0] _RAND_0;
  wire  _EVAL_32;
  reg [1:0] _EVAL_33;
  reg [31:0] _RAND_1;
  wire [32:0] _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire [32:0] _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire [3:0] _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire [7:0] _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire [32:0] _EVAL_55;
  wire  _EVAL_56;
  wire [7:0] _EVAL_57;
  wire  _EVAL_58;
  wire [3:0] _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire [31:0] _EVAL_63;
  wire [31:0] _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire [32:0] _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire [1:0] _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire [1:0] _EVAL_88;
  wire [7:0] _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  reg [5:0] _EVAL_92;
  reg [31:0] _RAND_2;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  reg  _EVAL_96;
  reg [31:0] _RAND_3;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_106;
  wire [32:0] _EVAL_107;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire [1:0] _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  reg [1:0] _EVAL_134;
  reg [31:0] _RAND_4;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire [22:0] _EVAL_137;
  wire [6:0] _EVAL_138;
  reg [3:0] _EVAL_139;
  reg [31:0] _RAND_5;
  reg  _EVAL_140;
  reg [31:0] _RAND_6;
  wire  _EVAL_141;
  wire [32:0] _EVAL_142;
  wire [1:0] _EVAL_143;
  wire [31:0] _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire [1:0] _EVAL_147;
  wire  _EVAL_148;
  wire [7:0] _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire [31:0] _EVAL_152;
  wire [32:0] _EVAL_154;
  wire [5:0] _EVAL_155;
  wire [3:0] _EVAL_156;
  wire [1:0] _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire [5:0] _EVAL_162;
  wire  _EVAL_163;
  reg [31:0] _EVAL_164;
  reg [31:0] _RAND_7;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire [32:0] _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire [6:0] _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire [32:0] _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_196;
  wire [31:0] _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire [32:0] _EVAL_200;
  wire [1:0] _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire [31:0] _EVAL_204;
  wire  _EVAL_205;
  wire [32:0] _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  reg [5:0] _EVAL_215;
  reg [31:0] _RAND_8;
  wire  _EVAL_216;
  wire  _EVAL_217;
  reg [2:0] _EVAL_218;
  reg [31:0] _RAND_9;
  wire [1:0] _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire [3:0] _EVAL_227;
  wire  _EVAL_228;
  wire [32:0] _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  reg  _EVAL_234;
  reg [31:0] _RAND_10;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire [5:0] _EVAL_237;
  wire [22:0] _EVAL_238;
  wire  _EVAL_239;
  reg [2:0] _EVAL_240;
  reg [31:0] _RAND_11;
  wire [1:0] _EVAL_241;
  wire  _EVAL_242;
  wire [1:0] _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire [5:0] _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire [1:0] _EVAL_258;
  wire [5:0] _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire [32:0] _EVAL_263;
  wire [32:0] _EVAL_264;
  wire  _EVAL_265;
  wire [31:0] _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire [1:0] _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_272;
  reg [5:0] _EVAL_273;
  reg [31:0] _RAND_12;
  wire [5:0] _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  reg [2:0] _EVAL_278;
  reg [31:0] _RAND_13;
  wire  _EVAL_279;
  wire [6:0] _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire [32:0] _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  reg [31:0] _EVAL_293;
  reg [31:0] _RAND_14;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  reg [3:0] _EVAL_298;
  reg [31:0] _RAND_15;
  wire  _EVAL_299;
  wire [32:0] _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire [31:0] _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire [32:0] _EVAL_321;
  reg  _EVAL_322;
  reg [31:0] _RAND_16;
  wire  _EVAL_323;
  wire  _EVAL_324;
  wire [32:0] _EVAL_325;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_50 = $signed(_EVAL_69) == 33'sh0;
  assign _EVAL_245 = ~_EVAL_310;
  assign _EVAL_228 = _EVAL_214 | _EVAL_16;
  assign _EVAL_264 = $signed(_EVAL_178) & -33'sh1000;
  assign _EVAL_171 = ~_EVAL_71;
  assign _EVAL_198 = _EVAL_3 == 3'h5;
  assign _EVAL_104 = _EVAL_4 == _EVAL_96;
  assign _EVAL_295 = ~_EVAL_210;
  assign _EVAL_256 = ~_EVAL_252;
  assign _EVAL_166 = _EVAL_15 == 3'h3;
  assign _EVAL_306 = _EVAL_15 == 3'h1;
  assign _EVAL_266 = _EVAL_263[31:0];
  assign _EVAL_121 = ~_EVAL_160;
  assign _EVAL_209 = _EVAL_11 & _EVAL_166;
  assign _EVAL_60 = _EVAL_3 == 3'h4;
  assign _EVAL_145 = ~_EVAL_175;
  assign _EVAL_192 = _EVAL_205 | _EVAL_16;
  assign _EVAL_248 = _EVAL_290 | _EVAL_16;
  assign _EVAL_288 = $signed(_EVAL_39) & -33'sh5000;
  assign _EVAL_276 = ~_EVAL_23;
  assign _EVAL_216 = _EVAL_181 | _EVAL_16;
  assign _EVAL_323 = _EVAL_8 == _EVAL_322;
  assign _EVAL_208 = _EVAL_211 | _EVAL_203;
  assign _EVAL_312 = _EVAL_123 | _EVAL_265;
  assign _EVAL_110 = _EVAL_15 == 3'h0;
  assign _EVAL_99 = ~_EVAL_318;
  assign _EVAL_55 = _EVAL_167;
  assign _EVAL_78 = ~_EVAL_314;
  assign _EVAL_265 = _EVAL_113 & _EVAL_267;
  assign _EVAL_202 = _EVAL_122 & _EVAL_211;
  assign _EVAL_48 = _EVAL_297 | _EVAL_165;
  assign _EVAL_113 = _EVAL_7 <= 4'h6;
  assign _EVAL_309 = ~_EVAL_193;
  assign _EVAL_117 = ~_EVAL_307;
  assign _EVAL_120 = $signed(_EVAL_206) == 33'sh0;
  assign _EVAL_207 = _EVAL_17 <= 3'h4;
  assign _EVAL_196 = _EVAL_15 == 3'h6;
  assign _EVAL_210 = _EVAL_35 | _EVAL_16;
  assign _EVAL_165 = _EVAL_130 & _EVAL_103;
  assign _EVAL_226 = _EVAL_12 != 2'h2;
  assign _EVAL_73 = $signed(_EVAL_229) == 33'sh0;
  assign _EVAL_125 = _EVAL_164 < plusarg_reader_out;
  assign _EVAL_87 = _EVAL_12 <= 2'h2;
  assign _EVAL_324 = _EVAL_73 | _EVAL_235;
  assign _EVAL_243 = 2'h1 << _EVAL_4;
  assign _EVAL_237 = _EVAL_20[5:0];
  assign _EVAL_128 = _EVAL_25 | _EVAL_16;
  assign _EVAL_74 = 2'h1 << _EVAL_151;
  assign _EVAL_263 = _EVAL_164 + 32'h1;
  assign _EVAL_27 = _EVAL_157[0];
  assign _EVAL_64 = _EVAL_1 ^ 32'h40000000;
  assign _EVAL_270 = _EVAL_252 & _EVAL_65;
  assign _EVAL_95 = _EVAL_312 | _EVAL_225;
  assign _EVAL_155 = _EVAL_172[5:0];
  assign _EVAL_291 = _EVAL_3 == 3'h2;
  assign _EVAL_181 = _EVAL_2 == _EVAL_234;
  assign _EVAL_45 = _EVAL_148 | _EVAL_184;
  assign _EVAL_77 = _EVAL_315 | _EVAL_102;
  assign _EVAL_86 = _EVAL_316 | _EVAL_16;
  assign _EVAL_172 = _EVAL_273 - 6'h1;
  assign _EVAL_124 = _EVAL_226 | _EVAL_16;
  assign _EVAL_51 = ~_EVAL_212;
  assign _EVAL_287 = _EVAL_11 & _EVAL_182;
  assign _EVAL_244 = _EVAL_122 & _EVAL_203;
  assign _EVAL_136 = _EVAL_15 == 3'h4;
  assign _EVAL_183 = _EVAL_301 & _EVAL_29;
  assign _EVAL_313 = _EVAL_50 | _EVAL_235;
  assign _EVAL_131 = _EVAL_104 | _EVAL_16;
  assign _EVAL_44 = _EVAL_43 | _EVAL_203;
  assign _EVAL_269 = _EVAL_241 & _EVAL_147;
  assign _EVAL_177 = _EVAL_255 | _EVAL_16;
  assign _EVAL_320 = _EVAL_130 & _EVAL_270;
  assign _EVAL_231 = _EVAL_18 & _EVAL_60;
  assign _EVAL_197 = _EVAL_1 ^ 32'h80000000;
  assign _EVAL_285 = ~_EVAL_28;
  assign _EVAL_290 = ~_EVAL_61;
  assign _EVAL_301 = _EVAL_102 & _EVAL_111;
  assign _EVAL_123 = _EVAL_122 & _EVAL_208;
  assign _EVAL_261 = _EVAL_18 & _EVAL_37;
  assign _EVAL_61 = _EVAL_258[0];
  assign _EVAL_62 = _EVAL_282 | _EVAL_125;
  assign _EVAL_144 = _EVAL_1 ^ 32'h3000;
  assign _EVAL_151 = _EVAL_7[0];
  assign _EVAL_112 = _EVAL_256 & _EVAL_180;
  assign _EVAL_25 = _EVAL_122 & _EVAL_44;
  assign _EVAL_180 = ~_EVAL_65;
  assign _EVAL_325 = {1'b0,$signed(_EVAL_64)};
  assign _EVAL_53 = ~_EVAL_67;
  assign _EVAL_149 = ~_EVAL_89;
  assign _EVAL_94 = _EVAL_17 == _EVAL_218;
  assign _EVAL_138 = _EVAL_215 - 6'h1;
  assign _EVAL_119 = _EVAL_62 | _EVAL_16;
  assign _EVAL_65 = _EVAL_1[0];
  assign _EVAL_242 = ~_EVAL_16;
  assign _EVAL_36 = ~_EVAL_233;
  assign _EVAL_294 = _EVAL_11 & _EVAL_110;
  assign _EVAL_84 = ~_EVAL_279;
  assign _EVAL_106 = ~_EVAL_192;
  assign _EVAL_255 = ~_EVAL_13;
  assign _EVAL_251 = _EVAL_152 == 32'h0;
  assign _EVAL_170 = ~_EVAL_221;
  assign _EVAL_129 = _EVAL_74 | 2'h1;
  assign _EVAL_259 = _EVAL_149[7:2];
  assign _EVAL_223 = _EVAL_12 == _EVAL_134;
  assign _EVAL_319 = _EVAL_102 & _EVAL_160;
  assign _EVAL_111 = _EVAL_273 == 6'h0;
  assign _EVAL_107 = $signed(_EVAL_34) & -33'sh1000000;
  assign _EVAL_148 = _EVAL_214 | _EVAL_217;
  assign _EVAL_66 = _EVAL_11 & _EVAL_136;
  assign _EVAL_163 = ~_EVAL_146;
  assign _EVAL_97 = _EVAL_11 & _EVAL_232;
  assign _EVAL_29 = ~_EVAL_222;
  assign _EVAL_58 = ~_EVAL_169;
  assign _EVAL_47 = _EVAL_0 & _EVAL_59;
  assign _EVAL_56 = ~_EVAL_38;
  assign _EVAL_220 = _EVAL_183 ? _EVAL_243 : 2'h0;
  assign _EVAL_277 = _EVAL_3 <= 3'h6;
  assign _EVAL_24 = _EVAL_11 & _EVAL_196;
  assign _EVAL_227 = {_EVAL_100,_EVAL_48,_EVAL_194,_EVAL_45};
  assign _EVAL_316 = _EVAL_10 == _EVAL_140;
  assign _EVAL_23 = _EVAL_289 | _EVAL_16;
  assign _EVAL_205 = _EVAL_17 == 3'h0;
  assign _EVAL_186 = _EVAL_3 == 3'h1;
  assign _EVAL_311 = ~_EVAL_228;
  assign _EVAL_238 = 23'hff << _EVAL_7;
  assign _EVAL_321 = {1'b0,$signed(_EVAL_197)};
  assign _EVAL_59 = ~_EVAL_227;
  assign _EVAL_39 = {1'b0,$signed(_EVAL_1)};
  assign _EVAL_178 = {1'b0,$signed(_EVAL_144)};
  assign _EVAL_75 = _EVAL_15[2];
  assign _EVAL_146 = _EVAL_141 | _EVAL_16;
  assign _EVAL_67 = _EVAL_292 | _EVAL_16;
  assign _EVAL_310 = _EVAL_286 | _EVAL_16;
  assign _EVAL_80 = ~_EVAL_119;
  assign _EVAL_156 = ~_EVAL_0;
  assign _EVAL_289 = _EVAL_15 == _EVAL_240;
  assign _EVAL_76 = ~_EVAL_131;
  assign _EVAL_307 = _EVAL_87 | _EVAL_16;
  assign _EVAL_152 = _EVAL_1 & _EVAL_63;
  assign _EVAL_90 = ~_EVAL_216;
  assign _EVAL_194 = _EVAL_148 | _EVAL_49;
  assign _EVAL_249 = ~_EVAL_257;
  assign _EVAL_203 = $signed(_EVAL_30) == 33'sh0;
  assign _EVAL_40 = ~_EVAL_81;
  assign _EVAL_57 = _EVAL_238[7:0];
  assign _EVAL_30 = _EVAL_200;
  assign _EVAL_85 = _EVAL_3 == _EVAL_278;
  assign _EVAL_303 = _EVAL_15 == 3'h2;
  assign _EVAL_82 = _EVAL_15 == 3'h5;
  assign _EVAL_100 = _EVAL_297 | _EVAL_320;
  assign _EVAL_20 = _EVAL_92 - 6'h1;
  assign _EVAL_189 = _EVAL_17 != 3'h0;
  assign _EVAL_115 = _EVAL_215 == 6'h0;
  assign _EVAL_89 = _EVAL_137[7:0];
  assign _EVAL_28 = _EVAL_132 | _EVAL_16;
  assign _EVAL_193 = _EVAL_95 | _EVAL_16;
  assign _EVAL_239 = _EVAL_11 & _EVAL_303;
  assign _EVAL_169 = _EVAL_173 | _EVAL_16;
  assign _EVAL_257 = _EVAL_27 | _EVAL_16;
  assign _EVAL_162 = _EVAL_138[5:0];
  assign _EVAL_130 = _EVAL_129[0];
  assign _EVAL_254 = _EVAL_47 == 4'h0;
  assign _EVAL_102 = _EVAL_9 & _EVAL_18;
  assign _EVAL_185 = _EVAL_275 | _EVAL_16;
  assign _EVAL_83 = _EVAL_11 & _EVAL_306;
  assign _EVAL_315 = _EVAL_6 & _EVAL_11;
  assign _EVAL_274 = _EVAL_280[5:0];
  assign _EVAL_141 = _EVAL_17 <= 3'h3;
  assign _EVAL_35 = ~_EVAL_14;
  assign _EVAL_211 = _EVAL_324 | _EVAL_120;
  assign _EVAL_292 = _EVAL_12 == 2'h0;
  assign _EVAL_213 = _EVAL >= 4'h2;
  assign _EVAL_173 = _EVAL_7 == _EVAL_298;
  assign _EVAL_93 = ~_EVAL_101;
  assign _EVAL_236 = ~_EVAL_126;
  assign _EVAL_147 = ~_EVAL_220;
  assign _EVAL_158 = ~_EVAL_177;
  assign _EVAL_167 = $signed(_EVAL_325) & -33'sh2000;
  assign _EVAL_135 = _EVAL_129[1];
  assign _EVAL_272 = _EVAL_156 == 4'h0;
  assign _EVAL_199 = _EVAL_315 & _EVAL_262;
  assign _EVAL_63 = {{24'd0}, _EVAL_52};
  assign _EVAL_81 = _EVAL_189 | _EVAL_16;
  assign _EVAL_200 = $signed(_EVAL_142) & -33'sh2000;
  assign _EVAL_70 = plusarg_reader_out == 32'h0;
  assign _EVAL_300 = _EVAL_107;
  assign _EVAL_79 = ~_EVAL_179;
  assign _EVAL_150 = ~_EVAL_72;
  assign _EVAL_317 = ~_EVAL_26;
  assign _EVAL_38 = _EVAL_213 | _EVAL_16;
  assign _EVAL_297 = _EVAL_214 | _EVAL_46;
  assign _EVAL_225 = _EVAL_308 & _EVAL_50;
  assign _EVAL_280 = _EVAL_31 - 6'h1;
  assign _EVAL_318 = _EVAL_19 | _EVAL_16;
  assign _EVAL_253 = _EVAL_52[7:2];
  assign _EVAL_222 = _EVAL_3 == 3'h6;
  assign _EVAL_42 = _EVAL_202 | _EVAL_225;
  assign _EVAL_262 = _EVAL_31 == 6'h0;
  assign _EVAL_176 = _EVAL_265 | _EVAL_225;
  assign _EVAL_302 = _EVAL_315 & _EVAL_115;
  assign _EVAL_284 = ~_EVAL_161;
  assign _EVAL_26 = _EVAL_33 != 2'h0;
  assign _EVAL_126 = _EVAL_109 | _EVAL_16;
  assign _EVAL_224 = _EVAL_207 | _EVAL_16;
  assign _EVAL_260 = ~_EVAL_248;
  assign _EVAL_157 = _EVAL_201 >> _EVAL_4;
  assign _EVAL_37 = _EVAL_3 == 3'h0;
  assign _EVAL_43 = _EVAL_313 | _EVAL_120;
  assign _EVAL_283 = _EVAL_88 != 2'h0;
  assign _EVAL_214 = _EVAL_7 >= 4'h2;
  assign _EVAL_142 = {1'b0,$signed(_EVAL_305)};
  assign _EVAL_32 = ~_EVAL_124;
  assign _EVAL_206 = _EVAL_288;
  assign _EVAL_101 = _EVAL_22 | _EVAL_16;
  assign _EVAL_34 = {1'b0,$signed(_EVAL_204)};
  assign _EVAL_160 = _EVAL_92 == 6'h0;
  assign _EVAL_98 = ~_EVAL_246;
  assign _EVAL_188 = ~_EVAL_185;
  assign _EVAL_133 = _EVAL_54 | _EVAL_68;
  assign _EVAL_282 = _EVAL_317 | _EVAL_70;
  assign _EVAL_184 = _EVAL_130 & _EVAL_112;
  assign _EVAL_72 = _EVAL_254 | _EVAL_16;
  assign _EVAL_258 = _EVAL_33 >> _EVAL_2;
  assign _EVAL_279 = _EVAL_223 | _EVAL_16;
  assign _EVAL_122 = _EVAL_7 <= 4'h2;
  assign _EVAL_46 = _EVAL_135 & _EVAL_252;
  assign _EVAL_305 = _EVAL_1 ^ 32'h20000000;
  assign _EVAL_49 = _EVAL_130 & _EVAL_168;
  assign _EVAL_247 = _EVAL_18 & _EVAL_222;
  assign _EVAL_296 = _EVAL_18 & _EVAL_186;
  assign _EVAL_233 = _EVAL_230 | _EVAL_16;
  assign _EVAL_179 = _EVAL_133 | _EVAL_16;
  assign _EVAL_159 = _EVAL_3[0];
  assign _EVAL_88 = _EVAL_199 ? _EVAL_143 : 2'h0;
  assign _EVAL_281 = _EVAL_18 & _EVAL_291;
  assign _EVAL_91 = ~_EVAL_128;
  assign _EVAL_154 = $signed(_EVAL_321) & -33'shc000;
  assign _EVAL_116 = _EVAL_272 | _EVAL_16;
  assign _EVAL_241 = _EVAL_33 | _EVAL_88;
  assign _EVAL_246 = _EVAL_42 | _EVAL_16;
  assign _EVAL_212 = _EVAL_251 | _EVAL_16;
  assign _EVAL_187 = ~_EVAL_224;
  assign _EVAL_52 = ~_EVAL_57;
  assign _EVAL_299 = _EVAL_11 & _EVAL_82;
  assign _EVAL_168 = _EVAL_256 & _EVAL_65;
  assign _EVAL_54 = _EVAL_88 != _EVAL_220;
  assign _EVAL_71 = _EVAL_21 | _EVAL_16;
  assign _EVAL_22 = _EVAL_17 <= 3'h2;
  assign _EVAL_217 = _EVAL_135 & _EVAL_256;
  assign _EVAL_268 = ~_EVAL_116;
  assign _EVAL_68 = ~_EVAL_283;
  assign _EVAL_19 = _EVAL_132 | _EVAL_14;
  assign _EVAL_175 = _EVAL_94 | _EVAL_16;
  assign _EVAL_314 = _EVAL_323 | _EVAL_16;
  assign _EVAL_230 = _EVAL_0 == _EVAL_227;
  assign _EVAL_69 = _EVAL_264;
  assign _EVAL_232 = ~_EVAL_115;
  assign _EVAL_182 = _EVAL_15 == 3'h7;
  assign _EVAL_275 = _EVAL == _EVAL_139;
  assign _EVAL_161 = _EVAL_85 | _EVAL_16;
  assign _EVAL_132 = ~_EVAL_8;
  assign _EVAL_204 = _EVAL_1 ^ 32'h2000000;
  assign _EVAL_267 = $signed(_EVAL_55) == 33'sh0;
  assign _EVAL_103 = _EVAL_252 & _EVAL_180;
  assign _EVAL_235 = $signed(_EVAL_300) == 33'sh0;
  assign _EVAL_109 = _EVAL_1 == _EVAL_293;
  assign _EVAL_250 = ~_EVAL_86;
  assign _EVAL_229 = _EVAL_154;
  assign _EVAL_118 = _EVAL_18 & _EVAL_121;
  assign _EVAL_127 = _EVAL_18 & _EVAL_198;
  assign _EVAL_252 = _EVAL_1[1];
  assign _EVAL_21 = _EVAL_17 <= 3'h1;
  assign _EVAL_137 = 23'hff << _EVAL;
  assign _EVAL_174 = ~_EVAL_75;
  assign _EVAL_286 = _EVAL_176 | _EVAL_244;
  assign _EVAL_201 = _EVAL_88 | _EVAL_33;
  assign _EVAL_308 = _EVAL_7 <= 4'h8;
  assign _EVAL_143 = 2'h1 << _EVAL_2;
  assign _EVAL_221 = _EVAL_277 | _EVAL_16;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_31 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_33 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_92 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_96 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_134 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_139 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_140 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_164 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_215 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_218 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_234 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_240 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_273 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_278 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_293 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_298 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_322 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_5) begin
    if (_EVAL_16) begin
      _EVAL_31 <= 6'h0;
    end else if (_EVAL_315) begin
      if (_EVAL_262) begin
        if (_EVAL_174) begin
          _EVAL_31 <= _EVAL_253;
        end else begin
          _EVAL_31 <= 6'h0;
        end
      end else begin
        _EVAL_31 <= _EVAL_274;
      end
    end
    if (_EVAL_16) begin
      _EVAL_33 <= 2'h0;
    end else begin
      _EVAL_33 <= _EVAL_269;
    end
    if (_EVAL_16) begin
      _EVAL_92 <= 6'h0;
    end else if (_EVAL_102) begin
      if (_EVAL_160) begin
        if (_EVAL_159) begin
          _EVAL_92 <= _EVAL_259;
        end else begin
          _EVAL_92 <= 6'h0;
        end
      end else begin
        _EVAL_92 <= _EVAL_237;
      end
    end
    if (_EVAL_319) begin
      _EVAL_96 <= _EVAL_4;
    end
    if (_EVAL_319) begin
      _EVAL_134 <= _EVAL_12;
    end
    if (_EVAL_319) begin
      _EVAL_139 <= _EVAL;
    end
    if (_EVAL_319) begin
      _EVAL_140 <= _EVAL_10;
    end
    if (_EVAL_16) begin
      _EVAL_164 <= 32'h0;
    end else if (_EVAL_77) begin
      _EVAL_164 <= 32'h0;
    end else begin
      _EVAL_164 <= _EVAL_266;
    end
    if (_EVAL_16) begin
      _EVAL_215 <= 6'h0;
    end else if (_EVAL_315) begin
      if (_EVAL_115) begin
        if (_EVAL_174) begin
          _EVAL_215 <= _EVAL_253;
        end else begin
          _EVAL_215 <= 6'h0;
        end
      end else begin
        _EVAL_215 <= _EVAL_162;
      end
    end
    if (_EVAL_302) begin
      _EVAL_218 <= _EVAL_17;
    end
    if (_EVAL_302) begin
      _EVAL_234 <= _EVAL_2;
    end
    if (_EVAL_302) begin
      _EVAL_240 <= _EVAL_15;
    end
    if (_EVAL_16) begin
      _EVAL_273 <= 6'h0;
    end else if (_EVAL_102) begin
      if (_EVAL_111) begin
        if (_EVAL_159) begin
          _EVAL_273 <= _EVAL_259;
        end else begin
          _EVAL_273 <= 6'h0;
        end
      end else begin
        _EVAL_273 <= _EVAL_155;
      end
    end
    if (_EVAL_319) begin
      _EVAL_278 <= _EVAL_3;
    end
    if (_EVAL_302) begin
      _EVAL_293 <= _EVAL_1;
    end
    if (_EVAL_302) begin
      _EVAL_298 <= _EVAL_7;
    end
    if (_EVAL_319) begin
      _EVAL_322 <= _EVAL_8;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fbec639)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24b53c84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6b601d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2311623)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c7edd79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_311) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(580a3bae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81e6e8c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f70a2cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8bc1f39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12b6cfb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd45e65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41ea3de8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c59db345)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59138e4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3afc8c94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(600bfe77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(972d6dae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fee5e2cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86704b9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ad2e16c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12571839)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8713448b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_311) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4257c170)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e69f04a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0b0bfc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac58bd0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bcd3e4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bf21e11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_284) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31d4dc58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c971df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d0934cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb841113)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(141cb4b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b296215)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f5c37fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a05834e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70cb1ddb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dfd0ff3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8153f534)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(413ddb52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8413df02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8b236a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f02288de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(494bbd2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(656f9ae0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b22621f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b03ad3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b65778bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_311) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(149fafb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d87329dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95221b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fd6ffa9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(249d0a44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7a0d144)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8e2b3f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bb05d5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7d9019b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6045112d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40ca7ad4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b91bdb48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(beb1bf11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53713af4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32cce197)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28c50f4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce783a54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(768a4027)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a263aab5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b2a5c98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffe2bbed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2409232)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48c6e2d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ce0c38a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cf2b741)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(530ce1d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_284) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_311) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd291055)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(472f913c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87b8f0af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
