//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_156_assert(
  input        _EVAL,
  input  [1:0] _EVAL_2,
  input        _EVAL_3,
  input        _EVAL_5,
  input        _EVAL_6,
  input        _EVAL_7,
  input        _EVAL_8,
  input        _EVAL_9,
  input  [1:0] _EVAL_11,
  input        _EVAL_13,
  input        _EVAL_15,
  input        _EVAL_16,
  input        _EVAL_18,
  input  [1:0] _EVAL_20,
  input        _EVAL_21,
  input        _EVAL_22,
  input        _EVAL_27,
  input        _EVAL_28,
  input        _EVAL_29,
  input  [1:0] _EVAL_30,
  input        _EVAL_31,
  input        _EVAL_33,
  input        _EVAL_44,
  input        _EVAL_54,
  input        _EVAL_57,
  input        _EVAL_78,
  input        _EVAL_94,
  input        _EVAL_118,
  input        _EVAL_167,
  input        _EVAL_169
);
  wire  _EVAL_36;
  wire  _EVAL_38;
  wire  _EVAL_40;
  wire  _EVAL_42;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire [2:0] _EVAL_53;
  wire  _EVAL_56;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_68;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_79;
  wire  _EVAL_82;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_90;
  wire  _EVAL_92;
  wire  _EVAL_95;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_117;
  wire  _EVAL_119;
  wire  _EVAL_122;
  wire  _EVAL_124;
  wire [2:0] _EVAL_126;
  wire [2:0] _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_144;
  wire  _EVAL_149;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_158;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire [2:0] _EVAL_166;
  wire  _EVAL_168;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_177;
  wire  _EVAL_180;
  wire  _EVAL_183;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_194;
  wire  _EVAL_197;
  assign _EVAL_68 = _EVAL_36 & _EVAL_185;
  assign _EVAL_48 = _EVAL_20 == 2'h3;
  assign _EVAL_87 = _EVAL_180 & _EVAL_112;
  assign _EVAL_153 = _EVAL_126 == 3'h1;
  assign _EVAL_151 = _EVAL_53 == 3'h3;
  assign _EVAL_109 = _EVAL_136 & _EVAL_48;
  assign _EVAL_185 = _EVAL_2 == 2'h1;
  assign _EVAL_70 = _EVAL_127 == 3'h3;
  assign _EVAL_47 = _EVAL_166 == 3'h3;
  assign _EVAL_190 = _EVAL_36 & _EVAL_112;
  assign _EVAL_71 = _EVAL_38 & _EVAL_149;
  assign _EVAL_127 = {_EVAL_18,_EVAL_6,_EVAL_9};
  assign _EVAL_166 = {_EVAL_31,_EVAL_7,_EVAL_16};
  assign _EVAL_168 = _EVAL_126 == 3'h7;
  assign _EVAL_136 = _EVAL_8 & _EVAL_78;
  assign _EVAL_154 = _EVAL_100 & _EVAL_122;
  assign _EVAL_165 = _EVAL_53 == 3'h7;
  assign _EVAL_79 = _EVAL_33 & _EVAL_167;
  assign _EVAL_194 = _EVAL_20 == 2'h2;
  assign _EVAL_117 = _EVAL_38 & _EVAL_122;
  assign _EVAL_90 = _EVAL_38 & _EVAL_107;
  assign _EVAL_149 = _EVAL_11 == 2'h1;
  assign _EVAL_171 = _EVAL_2 == 2'h3;
  assign _EVAL_119 = _EVAL_126 == 3'h5;
  assign _EVAL_133 = _EVAL_53 == 3'h0;
  assign _EVAL_50 = _EVAL_100 & _EVAL_107;
  assign _EVAL_92 = _EVAL_136 & _EVAL_194;
  assign _EVAL_65 = _EVAL_166 == 3'h0;
  assign _EVAL_64 = _EVAL_100 & _EVAL_149;
  assign _EVAL_36 = _EVAL_158 & _EVAL_44;
  assign _EVAL_40 = _EVAL_30 == 2'h2;
  assign _EVAL_122 = _EVAL_11 == 2'h3;
  assign _EVAL_86 = _EVAL_79 & _EVAL_189;
  assign _EVAL_180 = _EVAL_22 & _EVAL_44;
  assign _EVAL_46 = _EVAL_127 == 3'h4;
  assign _EVAL_104 = _EVAL_60 & _EVAL_74;
  assign _EVAL_53 = {_EVAL_21,_EVAL_29,_EVAL_27};
  assign _EVAL_188 = _EVAL_20 == 2'h0;
  assign _EVAL_60 = _EVAL_172 & _EVAL_78;
  assign _EVAL_52 = _EVAL_2 == 2'h0;
  assign _EVAL_114 = _EVAL_53 == 3'h4;
  assign _EVAL_99 = _EVAL_126 == 3'h4;
  assign _EVAL_155 = _EVAL_166 == 3'h7;
  assign _EVAL_164 = _EVAL_177 & _EVAL_103;
  assign _EVAL_186 = ~_EVAL_118;
  assign _EVAL_189 = _EVAL_30 == 2'h1;
  assign _EVAL_73 = _EVAL_127 == 3'h0;
  assign _EVAL_38 = _EVAL_186 & _EVAL_57;
  assign _EVAL_95 = _EVAL_53 == 3'h5;
  assign _EVAL_107 = _EVAL_11 == 2'h2;
  assign _EVAL_163 = _EVAL_180 & _EVAL_185;
  assign _EVAL_197 = ~_EVAL_94;
  assign _EVAL_111 = _EVAL_177 & _EVAL_40;
  assign _EVAL_158 = ~_EVAL_54;
  assign _EVAL_126 = {_EVAL_15,_EVAL_13,_EVAL_5};
  assign _EVAL_135 = _EVAL_79 & _EVAL_103;
  assign _EVAL_103 = _EVAL_30 == 2'h3;
  assign _EVAL_108 = _EVAL_127 == 3'h7;
  assign _EVAL_112 = _EVAL_2 == 2'h2;
  assign _EVAL_192 = _EVAL_127 == 3'h5;
  assign _EVAL_177 = _EVAL_197 & _EVAL_167;
  assign _EVAL_152 = _EVAL_60 & _EVAL_48;
  assign _EVAL_128 = _EVAL_79 & _EVAL_40;
  assign _EVAL_110 = _EVAL_166 == 3'h1;
  assign _EVAL_134 = _EVAL_166 == 3'h5;
  assign _EVAL_51 = _EVAL_136 & _EVAL_74;
  assign _EVAL_162 = _EVAL_166 == 3'h4;
  assign _EVAL_74 = _EVAL_20 == 2'h1;
  assign _EVAL_172 = ~_EVAL_169;
  assign _EVAL_115 = _EVAL_30 == 2'h0;
  assign _EVAL_56 = _EVAL_36 & _EVAL_171;
  assign _EVAL_59 = _EVAL_126 == 3'h3;
  assign _EVAL_42 = _EVAL_53 == 3'h1;
  assign _EVAL_124 = ~_EVAL_28;
  assign _EVAL_129 = _EVAL_127 == 3'h1;
  assign _EVAL_82 = _EVAL_60 & _EVAL_194;
  assign _EVAL_144 = _EVAL_180 & _EVAL_171;
  assign _EVAL_100 = _EVAL_3 & _EVAL_57;
  assign _EVAL_45 = _EVAL_177 & _EVAL_189;
  assign _EVAL_191 = _EVAL_11 == 2'h0;
  assign _EVAL_183 = _EVAL_126 == 3'h0;
  always @(posedge _EVAL) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(139b2fc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(394146e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56901a8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83b2d90a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc7fe073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a044c85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7237de2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3634d084)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7237de2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e7c1114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(139b2fc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e7c1114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80c29208)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab4a2067)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc9c4008)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7237de2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80c29208)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2b7c8bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2b7c8bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a362ac83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a044c85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fbd717)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a362ac83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(394146e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fbd717)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80c29208)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59d0eac9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e7c1114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a362ac83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a044c85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0e2c90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a044c85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83b2d90a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7237de2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(139b2fc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e7c1114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc9c4008)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56901a8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(139b2fc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59d0eac9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc9c4008)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80c29208)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59d0eac9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc7fe073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3634d084)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc9c4008)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc7fe073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83b2d90a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3634d084)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0e2c90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83b2d90a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(394146e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0e2c90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a362ac83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59d0eac9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab4a2067)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_8 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab4a2067)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56901a8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc7fe073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3634d084)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fbd717)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab4a2067)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fbd717)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2b7c8bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0e2c90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(394146e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56901a8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2b7c8bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
