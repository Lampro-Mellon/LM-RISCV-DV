//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_107(
  input  [31:0] _EVAL,
  input         _EVAL_0,
  output [3:0]  _EVAL_1,
  output [2:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [31:0] _EVAL_7,
  output [31:0] _EVAL_8,
  input  [1:0]  _EVAL_9,
  input  [31:0] _EVAL_10,
  output        _EVAL_11,
  input         _EVAL_12,
  output [29:0] _EVAL_13,
  input  [2:0]  _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16,
  input  [1:0]  _EVAL_17,
  output        _EVAL_18,
  input  [2:0]  _EVAL_19,
  output [3:0]  _EVAL_20,
  output [2:0]  _EVAL_21,
  output [11:0] _EVAL_22,
  input         _EVAL_23,
  output        _EVAL_24,
  output [31:0] _EVAL_25,
  output [1:0]  _EVAL_26,
  output [1:0]  _EVAL_27,
  output        _EVAL_28,
  output [2:0]  _EVAL_29,
  output [1:0]  _EVAL_30,
  output        _EVAL_31,
  output [31:0] _EVAL_32,
  input  [1:0]  _EVAL_34,
  input         _EVAL_35,
  output        _EVAL_36,
  output [2:0]  _EVAL_37,
  input         _EVAL_38,
  output        _EVAL_39,
  input         _EVAL_40,
  input  [31:0] _EVAL_41,
  input         _EVAL_42,
  input         _EVAL_43,
  output [25:0] _EVAL_44,
  output [3:0]  _EVAL_45,
  output [2:0]  _EVAL_46,
  output [2:0]  _EVAL_47,
  input  [2:0]  _EVAL_48,
  input  [3:0]  _EVAL_49,
  input  [2:0]  _EVAL_50,
  output [3:0]  _EVAL_51,
  output        _EVAL_52,
  input  [2:0]  _EVAL_54,
  output [31:0] _EVAL_55,
  output        _EVAL_56,
  input         _EVAL_57,
  output [31:0] _EVAL_58,
  input         _EVAL_59,
  output        _EVAL_60,
  input  [31:0] _EVAL_61,
  input  [3:0]  _EVAL_62,
  input         _EVAL_63,
  output [14:0] _EVAL_64,
  output [2:0]  _EVAL_65,
  input  [29:0] _EVAL_66,
  input         _EVAL_67,
  output [1:0]  _EVAL_68,
  input  [2:0]  _EVAL_69,
  output        _EVAL_70,
  output        _EVAL_71,
  output [2:0]  _EVAL_72,
  output        _EVAL_73,
  input  [2:0]  _EVAL_74,
  input         _EVAL_75,
  output [2:0]  _EVAL_76,
  output        _EVAL_77,
  output        _EVAL_78,
  output [3:0]  _EVAL_79,
  input         _EVAL_80,
  output [2:0]  _EVAL_81,
  output [2:0]  _EVAL_82,
  input         _EVAL_83,
  input         _EVAL_84,
  output [1:0]  _EVAL_85,
  output        _EVAL_86,
  output [2:0]  _EVAL_87,
  input         _EVAL_88,
  input  [2:0]  _EVAL_89,
  output        _EVAL_90
);
  wire [2:0] coupler_to_testIndicator__EVAL;
  wire  coupler_to_testIndicator__EVAL_0;
  wire  coupler_to_testIndicator__EVAL_1;
  wire  coupler_to_testIndicator__EVAL_2;
  wire [1:0] coupler_to_testIndicator__EVAL_3;
  wire [1:0] coupler_to_testIndicator__EVAL_4;
  wire [31:0] coupler_to_testIndicator__EVAL_5;
  wire  coupler_to_testIndicator__EVAL_6;
  wire  coupler_to_testIndicator__EVAL_7;
  wire  coupler_to_testIndicator__EVAL_8;
  wire [3:0] coupler_to_testIndicator__EVAL_9;
  wire  coupler_to_testIndicator__EVAL_10;
  wire  coupler_to_testIndicator__EVAL_11;
  wire [31:0] coupler_to_testIndicator__EVAL_12;
  wire [14:0] coupler_to_testIndicator__EVAL_13;
  wire [1:0] coupler_to_testIndicator__EVAL_14;
  wire [2:0] coupler_to_testIndicator__EVAL_15;
  wire [2:0] coupler_to_testIndicator__EVAL_16;
  wire  coupler_to_testIndicator__EVAL_17;
  wire [1:0] coupler_to_testIndicator__EVAL_18;
  wire [3:0] coupler_to_testIndicator__EVAL_19;
  wire [2:0] coupler_to_testIndicator__EVAL_20;
  wire [2:0] coupler_to_testIndicator__EVAL_21;
  wire [2:0] coupler_to_testIndicator__EVAL_22;
  wire [31:0] coupler_to_testIndicator__EVAL_23;
  wire  coupler_to_testIndicator__EVAL_24;
  wire [2:0] coupler_to_testIndicator__EVAL_25;
  wire [31:0] coupler_to_testIndicator__EVAL_26;
  wire [14:0] coupler_to_testIndicator__EVAL_27;
  wire  coupler_to_testIndicator__EVAL_28;
  wire [2:0] coupler_to_testIndicator__EVAL_29;
  wire [2:0] coupler_to_testIndicator__EVAL_30;
  wire  coupler_to_testIndicator__EVAL_31;
  wire [2:0] coupler_to_testIndicator__EVAL_32;
  wire  buffer__EVAL;
  wire [1:0] buffer__EVAL_0;
  wire  buffer__EVAL_1;
  wire  buffer__EVAL_2;
  wire  buffer__EVAL_3;
  wire  buffer__EVAL_4;
  wire [2:0] buffer__EVAL_5;
  wire  buffer__EVAL_6;
  wire [2:0] buffer__EVAL_7;
  wire  buffer__EVAL_8;
  wire  buffer__EVAL_9;
  wire [3:0] buffer__EVAL_10;
  wire  buffer__EVAL_11;
  wire  buffer__EVAL_12;
  wire  buffer__EVAL_13;
  wire  buffer__EVAL_14;
  wire [31:0] buffer__EVAL_15;
  wire  buffer__EVAL_16;
  wire [2:0] buffer__EVAL_17;
  wire  buffer__EVAL_18;
  wire  buffer__EVAL_19;
  wire  buffer__EVAL_20;
  wire [3:0] buffer__EVAL_21;
  wire  buffer__EVAL_22;
  wire [3:0] buffer__EVAL_23;
  wire [2:0] buffer__EVAL_24;
  wire  buffer__EVAL_25;
  wire  buffer__EVAL_26;
  wire [2:0] buffer__EVAL_27;
  wire  buffer__EVAL_28;
  wire [3:0] buffer__EVAL_29;
  wire  buffer__EVAL_30;
  wire  buffer__EVAL_31;
  wire  buffer__EVAL_32;
  wire [3:0] buffer__EVAL_33;
  wire [1:0] buffer__EVAL_34;
  wire [2:0] buffer__EVAL_35;
  wire [29:0] buffer__EVAL_36;
  wire [3:0] buffer__EVAL_37;
  wire  buffer__EVAL_38;
  wire [31:0] buffer__EVAL_39;
  wire [29:0] buffer__EVAL_40;
  wire [2:0] buffer__EVAL_41;
  wire [2:0] buffer__EVAL_42;
  wire  buffer__EVAL_43;
  wire [31:0] buffer__EVAL_44;
  wire  buffer__EVAL_45;
  wire [2:0] buffer__EVAL_46;
  wire [2:0] buffer__EVAL_47;
  wire [31:0] buffer__EVAL_48;
  wire  wrapped_error_device__EVAL;
  wire [3:0] wrapped_error_device__EVAL_0;
  wire [1:0] wrapped_error_device__EVAL_1;
  wire  wrapped_error_device__EVAL_2;
  wire [2:0] wrapped_error_device__EVAL_3;
  wire  wrapped_error_device__EVAL_4;
  wire [2:0] wrapped_error_device__EVAL_5;
  wire [2:0] wrapped_error_device__EVAL_6;
  wire  wrapped_error_device__EVAL_7;
  wire  wrapped_error_device__EVAL_8;
  wire [13:0] wrapped_error_device__EVAL_9;
  wire [2:0] wrapped_error_device__EVAL_10;
  wire [3:0] wrapped_error_device__EVAL_11;
  wire [2:0] wrapped_error_device__EVAL_12;
  wire  wrapped_error_device__EVAL_13;
  wire  wrapped_error_device__EVAL_14;
  wire [3:0] wrapped_error_device__EVAL_15;
  wire [31:0] wrapped_error_device__EVAL_16;
  wire  wrapped_error_device__EVAL_17;
  wire  wrapped_error_device__EVAL_18;
  wire  wrapped_error_device__EVAL_19;
  wire [25:0] coupler_to_clic__EVAL;
  wire [2:0] coupler_to_clic__EVAL_0;
  wire  coupler_to_clic__EVAL_1;
  wire  coupler_to_clic__EVAL_2;
  wire [2:0] coupler_to_clic__EVAL_3;
  wire  coupler_to_clic__EVAL_4;
  wire [3:0] coupler_to_clic__EVAL_5;
  wire [3:0] coupler_to_clic__EVAL_6;
  wire  coupler_to_clic__EVAL_7;
  wire  coupler_to_clic__EVAL_8;
  wire [1:0] coupler_to_clic__EVAL_9;
  wire [2:0] coupler_to_clic__EVAL_10;
  wire  coupler_to_clic__EVAL_11;
  wire  coupler_to_clic__EVAL_12;
  wire [1:0] coupler_to_clic__EVAL_13;
  wire  coupler_to_clic__EVAL_14;
  wire  coupler_to_clic__EVAL_15;
  wire [2:0] coupler_to_clic__EVAL_16;
  wire  coupler_to_clic__EVAL_17;
  wire [2:0] coupler_to_clic__EVAL_18;
  wire  coupler_to_clic__EVAL_19;
  wire [25:0] coupler_to_clic__EVAL_20;
  wire [31:0] coupler_to_clic__EVAL_21;
  wire [2:0] coupler_to_clic__EVAL_22;
  wire [2:0] coupler_to_clic__EVAL_23;
  wire [1:0] coupler_to_clic__EVAL_24;
  wire [31:0] coupler_to_clic__EVAL_25;
  wire [31:0] coupler_to_clic__EVAL_26;
  wire [2:0] coupler_to_clic__EVAL_27;
  wire [2:0] coupler_to_clic__EVAL_28;
  wire [31:0] coupler_to_clic__EVAL_29;
  wire [1:0] coupler_to_clic__EVAL_30;
  wire  coupler_to_clic__EVAL_31;
  wire [2:0] coupler_to_clic__EVAL_32;
  wire [1:0] coupler_to_port_named_ahb_periph_port__EVAL;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_0;
  wire [29:0] coupler_to_port_named_ahb_periph_port__EVAL_1;
  wire [1:0] coupler_to_port_named_ahb_periph_port__EVAL_2;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_3;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_4;
  wire [31:0] coupler_to_port_named_ahb_periph_port__EVAL_5;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_6;
  wire [1:0] coupler_to_port_named_ahb_periph_port__EVAL_7;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_8;
  wire [2:0] coupler_to_port_named_ahb_periph_port__EVAL_9;
  wire [1:0] coupler_to_port_named_ahb_periph_port__EVAL_10;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_11;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_12;
  wire [29:0] coupler_to_port_named_ahb_periph_port__EVAL_13;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_14;
  wire [31:0] coupler_to_port_named_ahb_periph_port__EVAL_15;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_16;
  wire [2:0] coupler_to_port_named_ahb_periph_port__EVAL_17;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_18;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_19;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_20;
  wire [2:0] coupler_to_port_named_ahb_periph_port__EVAL_21;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_22;
  wire [2:0] coupler_to_port_named_ahb_periph_port__EVAL_23;
  wire [2:0] coupler_to_port_named_ahb_periph_port__EVAL_24;
  wire [31:0] coupler_to_port_named_ahb_periph_port__EVAL_25;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_26;
  wire [3:0] coupler_to_port_named_ahb_periph_port__EVAL_27;
  wire [31:0] coupler_to_port_named_ahb_periph_port__EVAL_28;
  wire [2:0] coupler_to_port_named_ahb_periph_port__EVAL_29;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_30;
  wire [3:0] coupler_to_port_named_ahb_periph_port__EVAL_31;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_32;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_33;
  wire [2:0] out_xbar__EVAL;
  wire  out_xbar__EVAL_0;
  wire [31:0] out_xbar__EVAL_1;
  wire [2:0] out_xbar__EVAL_2;
  wire [1:0] out_xbar__EVAL_3;
  wire [25:0] out_xbar__EVAL_4;
  wire  out_xbar__EVAL_5;
  wire [31:0] out_xbar__EVAL_6;
  wire  out_xbar__EVAL_7;
  wire [2:0] out_xbar__EVAL_8;
  wire [3:0] out_xbar__EVAL_9;
  wire  out_xbar__EVAL_10;
  wire [1:0] out_xbar__EVAL_11;
  wire [3:0] out_xbar__EVAL_12;
  wire  out_xbar__EVAL_13;
  wire [2:0] out_xbar__EVAL_14;
  wire [13:0] out_xbar__EVAL_15;
  wire [2:0] out_xbar__EVAL_16;
  wire  out_xbar__EVAL_17;
  wire  out_xbar__EVAL_18;
  wire [2:0] out_xbar__EVAL_19;
  wire  out_xbar__EVAL_20;
  wire [2:0] out_xbar__EVAL_21;
  wire  out_xbar__EVAL_22;
  wire [31:0] out_xbar__EVAL_23;
  wire  out_xbar__EVAL_24;
  wire [2:0] out_xbar__EVAL_25;
  wire [31:0] out_xbar__EVAL_26;
  wire  out_xbar__EVAL_27;
  wire [2:0] out_xbar__EVAL_28;
  wire  out_xbar__EVAL_29;
  wire  out_xbar__EVAL_30;
  wire  out_xbar__EVAL_31;
  wire [1:0] out_xbar__EVAL_32;
  wire  out_xbar__EVAL_33;
  wire [1:0] out_xbar__EVAL_34;
  wire  out_xbar__EVAL_35;
  wire  out_xbar__EVAL_36;
  wire [3:0] out_xbar__EVAL_37;
  wire [3:0] out_xbar__EVAL_38;
  wire [2:0] out_xbar__EVAL_39;
  wire  out_xbar__EVAL_40;
  wire [29:0] out_xbar__EVAL_41;
  wire [3:0] out_xbar__EVAL_42;
  wire [14:0] out_xbar__EVAL_43;
  wire [2:0] out_xbar__EVAL_44;
  wire [2:0] out_xbar__EVAL_45;
  wire [1:0] out_xbar__EVAL_46;
  wire [2:0] out_xbar__EVAL_47;
  wire  out_xbar__EVAL_48;
  wire [31:0] out_xbar__EVAL_49;
  wire [1:0] out_xbar__EVAL_50;
  wire  out_xbar__EVAL_51;
  wire [1:0] out_xbar__EVAL_52;
  wire  out_xbar__EVAL_53;
  wire [3:0] out_xbar__EVAL_54;
  wire [31:0] out_xbar__EVAL_55;
  wire [2:0] out_xbar__EVAL_56;
  wire  out_xbar__EVAL_57;
  wire  out_xbar__EVAL_58;
  wire [3:0] out_xbar__EVAL_59;
  wire [29:0] out_xbar__EVAL_60;
  wire  out_xbar__EVAL_61;
  wire [31:0] out_xbar__EVAL_62;
  wire  out_xbar__EVAL_63;
  wire  out_xbar__EVAL_64;
  wire  out_xbar__EVAL_65;
  wire  out_xbar__EVAL_66;
  wire [11:0] out_xbar__EVAL_67;
  wire [2:0] out_xbar__EVAL_68;
  wire  out_xbar__EVAL_69;
  wire [2:0] out_xbar__EVAL_70;
  wire  out_xbar__EVAL_71;
  wire  out_xbar__EVAL_72;
  wire [2:0] out_xbar__EVAL_73;
  wire  out_xbar__EVAL_74;
  wire [2:0] out_xbar__EVAL_75;
  wire [2:0] out_xbar__EVAL_76;
  wire [1:0] out_xbar__EVAL_77;
  wire [2:0] out_xbar__EVAL_78;
  wire  out_xbar__EVAL_79;
  wire  out_xbar__EVAL_80;
  wire  out_xbar__EVAL_81;
  wire  out_xbar__EVAL_82;
  wire [3:0] out_xbar__EVAL_83;
  wire  out_xbar__EVAL_84;
  wire [2:0] out_xbar__EVAL_85;
  wire  out_xbar__EVAL_86;
  wire  out_xbar__EVAL_87;
  wire [1:0] out_xbar__EVAL_88;
  wire [3:0] out_xbar__EVAL_89;
  wire [3:0] out_xbar__EVAL_90;
  wire  out_xbar__EVAL_91;
  wire [2:0] out_xbar__EVAL_92;
  wire [2:0] out_xbar__EVAL_93;
  wire [1:0] out_xbar__EVAL_94;
  wire [31:0] out_xbar__EVAL_95;
  wire  out_xbar__EVAL_96;
  wire [31:0] out_xbar__EVAL_97;
  wire [2:0] out_xbar__EVAL_98;
  wire [1:0] out_xbar__EVAL_99;
  wire [2:0] out_xbar__EVAL_100;
  wire  out_xbar__EVAL_101;
  wire  out_xbar__EVAL_102;
  wire [2:0] out_xbar__EVAL_103;
  wire [31:0] out_xbar__EVAL_104;
  wire  out_xbar__EVAL_105;
  wire  out_xbar__EVAL_106;
  wire  out_xbar__EVAL_107;
  wire  out_xbar__EVAL_108;
  wire [2:0] out_xbar__EVAL_109;
  wire [2:0] out_xbar__EVAL_110;
  wire  out_xbar__EVAL_111;
  wire [2:0] out_xbar__EVAL_112;
  wire [2:0] out_xbar__EVAL_113;
  wire [31:0] out_xbar__EVAL_114;
  wire  out_xbar__EVAL_115;
  wire  coupler_to_debug__EVAL;
  wire [3:0] coupler_to_debug__EVAL_0;
  wire [2:0] coupler_to_debug__EVAL_1;
  wire [31:0] coupler_to_debug__EVAL_2;
  wire [31:0] coupler_to_debug__EVAL_3;
  wire [2:0] coupler_to_debug__EVAL_4;
  wire  coupler_to_debug__EVAL_5;
  wire [11:0] coupler_to_debug__EVAL_6;
  wire  coupler_to_debug__EVAL_7;
  wire  coupler_to_debug__EVAL_8;
  wire [2:0] coupler_to_debug__EVAL_9;
  wire  coupler_to_debug__EVAL_10;
  wire  coupler_to_debug__EVAL_11;
  wire [2:0] coupler_to_debug__EVAL_12;
  wire [1:0] coupler_to_debug__EVAL_13;
  wire [1:0] coupler_to_debug__EVAL_14;
  wire [2:0] coupler_to_debug__EVAL_15;
  wire [3:0] coupler_to_debug__EVAL_16;
  wire [1:0] coupler_to_debug__EVAL_17;
  wire [2:0] coupler_to_debug__EVAL_18;
  wire  coupler_to_debug__EVAL_19;
  wire [2:0] coupler_to_debug__EVAL_20;
  wire [2:0] coupler_to_debug__EVAL_21;
  wire  coupler_to_debug__EVAL_22;
  wire  coupler_to_debug__EVAL_23;
  wire  coupler_to_debug__EVAL_24;
  wire [2:0] coupler_to_debug__EVAL_25;
  wire [31:0] coupler_to_debug__EVAL_26;
  wire [11:0] coupler_to_debug__EVAL_27;
  wire [31:0] coupler_to_debug__EVAL_28;
  wire  coupler_to_debug__EVAL_29;
  wire [1:0] coupler_to_debug__EVAL_30;
  wire [2:0] coupler_to_debug__EVAL_31;
  wire  coupler_to_debug__EVAL_32;
  wire  subsystem_cbus_clock_groups__EVAL_0;
  wire  subsystem_cbus_clock_groups__EVAL_4;
  wire  subsystem_cbus_clock_groups__EVAL_5;
  wire  subsystem_cbus_clock_groups__EVAL_6;
  wire  buffer_1__EVAL;
  wire  buffer_1__EVAL_0;
  wire [29:0] buffer_1__EVAL_1;
  wire  buffer_1__EVAL_2;
  wire  buffer_1__EVAL_3;
  wire  buffer_1__EVAL_4;
  wire  buffer_1__EVAL_5;
  wire  buffer_1__EVAL_6;
  wire [31:0] buffer_1__EVAL_7;
  wire [2:0] buffer_1__EVAL_8;
  wire [1:0] buffer_1__EVAL_9;
  wire  buffer_1__EVAL_10;
  wire [31:0] buffer_1__EVAL_11;
  wire  buffer_1__EVAL_12;
  wire [2:0] buffer_1__EVAL_13;
  wire [1:0] buffer_1__EVAL_14;
  wire [2:0] buffer_1__EVAL_15;
  wire [2:0] buffer_1__EVAL_16;
  wire [2:0] buffer_1__EVAL_17;
  wire  buffer_1__EVAL_18;
  wire [3:0] buffer_1__EVAL_19;
  wire  buffer_1__EVAL_20;
  wire [3:0] buffer_1__EVAL_21;
  wire  buffer_1__EVAL_22;
  wire [2:0] buffer_1__EVAL_23;
  wire [2:0] buffer_1__EVAL_24;
  wire [3:0] buffer_1__EVAL_25;
  wire [31:0] buffer_1__EVAL_26;
  wire  buffer_1__EVAL_27;
  wire  buffer_1__EVAL_28;
  wire [2:0] buffer_1__EVAL_29;
  wire  buffer_1__EVAL_30;
  wire  buffer_1__EVAL_31;
  wire [2:0] buffer_1__EVAL_32;
  wire  buffer_1__EVAL_33;
  wire [3:0] buffer_1__EVAL_34;
  wire  buffer_1__EVAL_35;
  wire [3:0] buffer_1__EVAL_36;
  wire  buffer_1__EVAL_37;
  wire [31:0] buffer_1__EVAL_38;
  wire  buffer_1__EVAL_39;
  wire [2:0] buffer_1__EVAL_40;
  wire  buffer_1__EVAL_41;
  wire  buffer_1__EVAL_42;
  wire [29:0] buffer_1__EVAL_43;
  wire  buffer_1__EVAL_44;
  wire  buffer_1__EVAL_45;
  wire  buffer_1__EVAL_46;
  wire  buffer_1__EVAL_47;
  wire  buffer_1__EVAL_48;
  wire  buffer_1__EVAL_49;
  wire  buffer_1__EVAL_50;
  wire  buffer_1__EVAL_51;
  wire [3:0] buffer_1__EVAL_52;
  wire  buffer_1__EVAL_53;
  wire  buffer_1__EVAL_54;
  wire [2:0] in_xbar__EVAL;
  wire  in_xbar__EVAL_0;
  wire  in_xbar__EVAL_1;
  wire [31:0] in_xbar__EVAL_2;
  wire  in_xbar__EVAL_3;
  wire [31:0] in_xbar__EVAL_4;
  wire [31:0] in_xbar__EVAL_5;
  wire [29:0] in_xbar__EVAL_6;
  wire [3:0] in_xbar__EVAL_7;
  wire  in_xbar__EVAL_8;
  wire  in_xbar__EVAL_9;
  wire  in_xbar__EVAL_10;
  wire  in_xbar__EVAL_11;
  wire  in_xbar__EVAL_12;
  wire  in_xbar__EVAL_13;
  wire  in_xbar__EVAL_14;
  wire [2:0] in_xbar__EVAL_15;
  wire  in_xbar__EVAL_16;
  wire [2:0] in_xbar__EVAL_17;
  wire [1:0] in_xbar__EVAL_18;
  wire  in_xbar__EVAL_19;
  wire  in_xbar__EVAL_20;
  wire  in_xbar__EVAL_21;
  wire [2:0] in_xbar__EVAL_22;
  wire [3:0] in_xbar__EVAL_23;
  wire  in_xbar__EVAL_24;
  wire  in_xbar__EVAL_25;
  wire  in_xbar__EVAL_26;
  wire  in_xbar__EVAL_27;
  wire  in_xbar__EVAL_28;
  wire  in_xbar__EVAL_29;
  wire [2:0] in_xbar__EVAL_30;
  wire [29:0] in_xbar__EVAL_31;
  wire [2:0] in_xbar__EVAL_32;
  wire [2:0] in_xbar__EVAL_33;
  wire  in_xbar__EVAL_34;
  wire  in_xbar__EVAL_35;
  wire  in_xbar__EVAL_36;
  wire  in_xbar__EVAL_37;
  wire [3:0] in_xbar__EVAL_38;
  wire  in_xbar__EVAL_39;
  wire  in_xbar__EVAL_40;
  wire [3:0] in_xbar__EVAL_41;
  wire [3:0] in_xbar__EVAL_42;
  wire  in_xbar__EVAL_43;
  wire [3:0] in_xbar__EVAL_44;
  wire [2:0] in_xbar__EVAL_45;
  wire  in_xbar__EVAL_46;
  wire [2:0] in_xbar__EVAL_47;
  wire [2:0] in_xbar__EVAL_48;
  wire [31:0] in_xbar__EVAL_49;
  wire  in_xbar__EVAL_50;
  wire  in_xbar__EVAL_51;
  wire  in_xbar__EVAL_52;
  wire  in_xbar__EVAL_53;
  wire [1:0] in_xbar__EVAL_54;
  wire  clockGroup__EVAL;
  wire  clockGroup__EVAL_0;
  wire  clockGroup__EVAL_1;
  wire  clockGroup__EVAL_2;
  wire  fixedClockNode__EVAL;
  wire  fixedClockNode__EVAL_0;
  wire  fixedClockNode__EVAL_1;
  wire  fixedClockNode__EVAL_2;
  wire  atomics__EVAL;
  wire [31:0] atomics__EVAL_0;
  wire  atomics__EVAL_1;
  wire  atomics__EVAL_2;
  wire [2:0] atomics__EVAL_3;
  wire  atomics__EVAL_4;
  wire [2:0] atomics__EVAL_5;
  wire [2:0] atomics__EVAL_6;
  wire [2:0] atomics__EVAL_7;
  wire [1:0] atomics__EVAL_8;
  wire  atomics__EVAL_9;
  wire  atomics__EVAL_10;
  wire [31:0] atomics__EVAL_11;
  wire [31:0] atomics__EVAL_12;
  wire  atomics__EVAL_13;
  wire  atomics__EVAL_14;
  wire  atomics__EVAL_15;
  wire  atomics__EVAL_16;
  wire  atomics__EVAL_17;
  wire [29:0] atomics__EVAL_18;
  wire  atomics__EVAL_19;
  wire  atomics__EVAL_20;
  wire  atomics__EVAL_21;
  wire  atomics__EVAL_22;
  wire [1:0] atomics__EVAL_23;
  wire [2:0] atomics__EVAL_24;
  wire [3:0] atomics__EVAL_25;
  wire [3:0] atomics__EVAL_26;
  wire  atomics__EVAL_27;
  wire [3:0] atomics__EVAL_28;
  wire  atomics__EVAL_29;
  wire [2:0] atomics__EVAL_30;
  wire  atomics__EVAL_31;
  wire  atomics__EVAL_32;
  wire [2:0] atomics__EVAL_33;
  wire  atomics__EVAL_34;
  wire [2:0] atomics__EVAL_35;
  wire [2:0] atomics__EVAL_36;
  wire [3:0] atomics__EVAL_37;
  wire  atomics__EVAL_38;
  wire  atomics__EVAL_39;
  wire [3:0] atomics__EVAL_40;
  wire [31:0] atomics__EVAL_41;
  wire  atomics__EVAL_42;
  wire  atomics__EVAL_43;
  wire  atomics__EVAL_44;
  wire [2:0] atomics__EVAL_45;
  wire  atomics__EVAL_46;
  wire  atomics__EVAL_47;
  wire  atomics__EVAL_48;
  wire  atomics__EVAL_49;
  wire [29:0] atomics__EVAL_50;
  wire [3:0] atomics__EVAL_51;
  wire [31:0] fixer__EVAL;
  wire  fixer__EVAL_0;
  wire  fixer__EVAL_1;
  wire  fixer__EVAL_2;
  wire [2:0] fixer__EVAL_3;
  wire  fixer__EVAL_4;
  wire  fixer__EVAL_5;
  wire [31:0] fixer__EVAL_6;
  wire [29:0] fixer__EVAL_7;
  wire [2:0] fixer__EVAL_8;
  wire  fixer__EVAL_9;
  wire  fixer__EVAL_10;
  wire [31:0] fixer__EVAL_11;
  wire  fixer__EVAL_12;
  wire [3:0] fixer__EVAL_13;
  wire  fixer__EVAL_14;
  wire  fixer__EVAL_15;
  wire [29:0] fixer__EVAL_16;
  wire [3:0] fixer__EVAL_17;
  wire  fixer__EVAL_18;
  wire [3:0] fixer__EVAL_19;
  wire [2:0] fixer__EVAL_20;
  wire [3:0] fixer__EVAL_21;
  wire [2:0] fixer__EVAL_22;
  wire  fixer__EVAL_23;
  wire [2:0] fixer__EVAL_24;
  wire [1:0] fixer__EVAL_25;
  wire  fixer__EVAL_26;
  wire [2:0] fixer__EVAL_27;
  wire [31:0] fixer__EVAL_28;
  wire  fixer__EVAL_29;
  wire  fixer__EVAL_30;
  wire  fixer__EVAL_31;
  wire  fixer__EVAL_32;
  wire [1:0] fixer__EVAL_33;
  wire  fixer__EVAL_34;
  wire [3:0] fixer__EVAL_35;
  wire  fixer__EVAL_36;
  wire  fixer__EVAL_37;
  wire [3:0] fixer__EVAL_38;
  wire [2:0] fixer__EVAL_39;
  wire  fixer__EVAL_40;
  wire  fixer__EVAL_41;
  wire  fixer__EVAL_42;
  wire  fixer__EVAL_43;
  wire [2:0] fixer__EVAL_44;
  wire [2:0] fixer__EVAL_45;
  wire  fixer__EVAL_46;
  wire  fixer__EVAL_47;
  wire [2:0] fixer__EVAL_48;
  _EVAL_102 coupler_to_testIndicator (
    ._EVAL(coupler_to_testIndicator__EVAL),
    ._EVAL_0(coupler_to_testIndicator__EVAL_0),
    ._EVAL_1(coupler_to_testIndicator__EVAL_1),
    ._EVAL_2(coupler_to_testIndicator__EVAL_2),
    ._EVAL_3(coupler_to_testIndicator__EVAL_3),
    ._EVAL_4(coupler_to_testIndicator__EVAL_4),
    ._EVAL_5(coupler_to_testIndicator__EVAL_5),
    ._EVAL_6(coupler_to_testIndicator__EVAL_6),
    ._EVAL_7(coupler_to_testIndicator__EVAL_7),
    ._EVAL_8(coupler_to_testIndicator__EVAL_8),
    ._EVAL_9(coupler_to_testIndicator__EVAL_9),
    ._EVAL_10(coupler_to_testIndicator__EVAL_10),
    ._EVAL_11(coupler_to_testIndicator__EVAL_11),
    ._EVAL_12(coupler_to_testIndicator__EVAL_12),
    ._EVAL_13(coupler_to_testIndicator__EVAL_13),
    ._EVAL_14(coupler_to_testIndicator__EVAL_14),
    ._EVAL_15(coupler_to_testIndicator__EVAL_15),
    ._EVAL_16(coupler_to_testIndicator__EVAL_16),
    ._EVAL_17(coupler_to_testIndicator__EVAL_17),
    ._EVAL_18(coupler_to_testIndicator__EVAL_18),
    ._EVAL_19(coupler_to_testIndicator__EVAL_19),
    ._EVAL_20(coupler_to_testIndicator__EVAL_20),
    ._EVAL_21(coupler_to_testIndicator__EVAL_21),
    ._EVAL_22(coupler_to_testIndicator__EVAL_22),
    ._EVAL_23(coupler_to_testIndicator__EVAL_23),
    ._EVAL_24(coupler_to_testIndicator__EVAL_24),
    ._EVAL_25(coupler_to_testIndicator__EVAL_25),
    ._EVAL_26(coupler_to_testIndicator__EVAL_26),
    ._EVAL_27(coupler_to_testIndicator__EVAL_27),
    ._EVAL_28(coupler_to_testIndicator__EVAL_28),
    ._EVAL_29(coupler_to_testIndicator__EVAL_29),
    ._EVAL_30(coupler_to_testIndicator__EVAL_30),
    ._EVAL_31(coupler_to_testIndicator__EVAL_31),
    ._EVAL_32(coupler_to_testIndicator__EVAL_32)
  );
  _EVAL_67 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32),
    ._EVAL_33(buffer__EVAL_33),
    ._EVAL_34(buffer__EVAL_34),
    ._EVAL_35(buffer__EVAL_35),
    ._EVAL_36(buffer__EVAL_36),
    ._EVAL_37(buffer__EVAL_37),
    ._EVAL_38(buffer__EVAL_38),
    ._EVAL_39(buffer__EVAL_39),
    ._EVAL_40(buffer__EVAL_40),
    ._EVAL_41(buffer__EVAL_41),
    ._EVAL_42(buffer__EVAL_42),
    ._EVAL_43(buffer__EVAL_43),
    ._EVAL_44(buffer__EVAL_44),
    ._EVAL_45(buffer__EVAL_45),
    ._EVAL_46(buffer__EVAL_46),
    ._EVAL_47(buffer__EVAL_47),
    ._EVAL_48(buffer__EVAL_48)
  );
  _EVAL_76 wrapped_error_device (
    ._EVAL(wrapped_error_device__EVAL),
    ._EVAL_0(wrapped_error_device__EVAL_0),
    ._EVAL_1(wrapped_error_device__EVAL_1),
    ._EVAL_2(wrapped_error_device__EVAL_2),
    ._EVAL_3(wrapped_error_device__EVAL_3),
    ._EVAL_4(wrapped_error_device__EVAL_4),
    ._EVAL_5(wrapped_error_device__EVAL_5),
    ._EVAL_6(wrapped_error_device__EVAL_6),
    ._EVAL_7(wrapped_error_device__EVAL_7),
    ._EVAL_8(wrapped_error_device__EVAL_8),
    ._EVAL_9(wrapped_error_device__EVAL_9),
    ._EVAL_10(wrapped_error_device__EVAL_10),
    ._EVAL_11(wrapped_error_device__EVAL_11),
    ._EVAL_12(wrapped_error_device__EVAL_12),
    ._EVAL_13(wrapped_error_device__EVAL_13),
    ._EVAL_14(wrapped_error_device__EVAL_14),
    ._EVAL_15(wrapped_error_device__EVAL_15),
    ._EVAL_16(wrapped_error_device__EVAL_16),
    ._EVAL_17(wrapped_error_device__EVAL_17),
    ._EVAL_18(wrapped_error_device__EVAL_18),
    ._EVAL_19(wrapped_error_device__EVAL_19)
  );
  _EVAL_79 coupler_to_clic (
    ._EVAL(coupler_to_clic__EVAL),
    ._EVAL_0(coupler_to_clic__EVAL_0),
    ._EVAL_1(coupler_to_clic__EVAL_1),
    ._EVAL_2(coupler_to_clic__EVAL_2),
    ._EVAL_3(coupler_to_clic__EVAL_3),
    ._EVAL_4(coupler_to_clic__EVAL_4),
    ._EVAL_5(coupler_to_clic__EVAL_5),
    ._EVAL_6(coupler_to_clic__EVAL_6),
    ._EVAL_7(coupler_to_clic__EVAL_7),
    ._EVAL_8(coupler_to_clic__EVAL_8),
    ._EVAL_9(coupler_to_clic__EVAL_9),
    ._EVAL_10(coupler_to_clic__EVAL_10),
    ._EVAL_11(coupler_to_clic__EVAL_11),
    ._EVAL_12(coupler_to_clic__EVAL_12),
    ._EVAL_13(coupler_to_clic__EVAL_13),
    ._EVAL_14(coupler_to_clic__EVAL_14),
    ._EVAL_15(coupler_to_clic__EVAL_15),
    ._EVAL_16(coupler_to_clic__EVAL_16),
    ._EVAL_17(coupler_to_clic__EVAL_17),
    ._EVAL_18(coupler_to_clic__EVAL_18),
    ._EVAL_19(coupler_to_clic__EVAL_19),
    ._EVAL_20(coupler_to_clic__EVAL_20),
    ._EVAL_21(coupler_to_clic__EVAL_21),
    ._EVAL_22(coupler_to_clic__EVAL_22),
    ._EVAL_23(coupler_to_clic__EVAL_23),
    ._EVAL_24(coupler_to_clic__EVAL_24),
    ._EVAL_25(coupler_to_clic__EVAL_25),
    ._EVAL_26(coupler_to_clic__EVAL_26),
    ._EVAL_27(coupler_to_clic__EVAL_27),
    ._EVAL_28(coupler_to_clic__EVAL_28),
    ._EVAL_29(coupler_to_clic__EVAL_29),
    ._EVAL_30(coupler_to_clic__EVAL_30),
    ._EVAL_31(coupler_to_clic__EVAL_31),
    ._EVAL_32(coupler_to_clic__EVAL_32)
  );
  _EVAL_97 coupler_to_port_named_ahb_periph_port (
    ._EVAL(coupler_to_port_named_ahb_periph_port__EVAL),
    ._EVAL_0(coupler_to_port_named_ahb_periph_port__EVAL_0),
    ._EVAL_1(coupler_to_port_named_ahb_periph_port__EVAL_1),
    ._EVAL_2(coupler_to_port_named_ahb_periph_port__EVAL_2),
    ._EVAL_3(coupler_to_port_named_ahb_periph_port__EVAL_3),
    ._EVAL_4(coupler_to_port_named_ahb_periph_port__EVAL_4),
    ._EVAL_5(coupler_to_port_named_ahb_periph_port__EVAL_5),
    ._EVAL_6(coupler_to_port_named_ahb_periph_port__EVAL_6),
    ._EVAL_7(coupler_to_port_named_ahb_periph_port__EVAL_7),
    ._EVAL_8(coupler_to_port_named_ahb_periph_port__EVAL_8),
    ._EVAL_9(coupler_to_port_named_ahb_periph_port__EVAL_9),
    ._EVAL_10(coupler_to_port_named_ahb_periph_port__EVAL_10),
    ._EVAL_11(coupler_to_port_named_ahb_periph_port__EVAL_11),
    ._EVAL_12(coupler_to_port_named_ahb_periph_port__EVAL_12),
    ._EVAL_13(coupler_to_port_named_ahb_periph_port__EVAL_13),
    ._EVAL_14(coupler_to_port_named_ahb_periph_port__EVAL_14),
    ._EVAL_15(coupler_to_port_named_ahb_periph_port__EVAL_15),
    ._EVAL_16(coupler_to_port_named_ahb_periph_port__EVAL_16),
    ._EVAL_17(coupler_to_port_named_ahb_periph_port__EVAL_17),
    ._EVAL_18(coupler_to_port_named_ahb_periph_port__EVAL_18),
    ._EVAL_19(coupler_to_port_named_ahb_periph_port__EVAL_19),
    ._EVAL_20(coupler_to_port_named_ahb_periph_port__EVAL_20),
    ._EVAL_21(coupler_to_port_named_ahb_periph_port__EVAL_21),
    ._EVAL_22(coupler_to_port_named_ahb_periph_port__EVAL_22),
    ._EVAL_23(coupler_to_port_named_ahb_periph_port__EVAL_23),
    ._EVAL_24(coupler_to_port_named_ahb_periph_port__EVAL_24),
    ._EVAL_25(coupler_to_port_named_ahb_periph_port__EVAL_25),
    ._EVAL_26(coupler_to_port_named_ahb_periph_port__EVAL_26),
    ._EVAL_27(coupler_to_port_named_ahb_periph_port__EVAL_27),
    ._EVAL_28(coupler_to_port_named_ahb_periph_port__EVAL_28),
    ._EVAL_29(coupler_to_port_named_ahb_periph_port__EVAL_29),
    ._EVAL_30(coupler_to_port_named_ahb_periph_port__EVAL_30),
    ._EVAL_31(coupler_to_port_named_ahb_periph_port__EVAL_31),
    ._EVAL_32(coupler_to_port_named_ahb_periph_port__EVAL_32),
    ._EVAL_33(coupler_to_port_named_ahb_periph_port__EVAL_33)
  );
  _EVAL_63 out_xbar (
    ._EVAL(out_xbar__EVAL),
    ._EVAL_0(out_xbar__EVAL_0),
    ._EVAL_1(out_xbar__EVAL_1),
    ._EVAL_2(out_xbar__EVAL_2),
    ._EVAL_3(out_xbar__EVAL_3),
    ._EVAL_4(out_xbar__EVAL_4),
    ._EVAL_5(out_xbar__EVAL_5),
    ._EVAL_6(out_xbar__EVAL_6),
    ._EVAL_7(out_xbar__EVAL_7),
    ._EVAL_8(out_xbar__EVAL_8),
    ._EVAL_9(out_xbar__EVAL_9),
    ._EVAL_10(out_xbar__EVAL_10),
    ._EVAL_11(out_xbar__EVAL_11),
    ._EVAL_12(out_xbar__EVAL_12),
    ._EVAL_13(out_xbar__EVAL_13),
    ._EVAL_14(out_xbar__EVAL_14),
    ._EVAL_15(out_xbar__EVAL_15),
    ._EVAL_16(out_xbar__EVAL_16),
    ._EVAL_17(out_xbar__EVAL_17),
    ._EVAL_18(out_xbar__EVAL_18),
    ._EVAL_19(out_xbar__EVAL_19),
    ._EVAL_20(out_xbar__EVAL_20),
    ._EVAL_21(out_xbar__EVAL_21),
    ._EVAL_22(out_xbar__EVAL_22),
    ._EVAL_23(out_xbar__EVAL_23),
    ._EVAL_24(out_xbar__EVAL_24),
    ._EVAL_25(out_xbar__EVAL_25),
    ._EVAL_26(out_xbar__EVAL_26),
    ._EVAL_27(out_xbar__EVAL_27),
    ._EVAL_28(out_xbar__EVAL_28),
    ._EVAL_29(out_xbar__EVAL_29),
    ._EVAL_30(out_xbar__EVAL_30),
    ._EVAL_31(out_xbar__EVAL_31),
    ._EVAL_32(out_xbar__EVAL_32),
    ._EVAL_33(out_xbar__EVAL_33),
    ._EVAL_34(out_xbar__EVAL_34),
    ._EVAL_35(out_xbar__EVAL_35),
    ._EVAL_36(out_xbar__EVAL_36),
    ._EVAL_37(out_xbar__EVAL_37),
    ._EVAL_38(out_xbar__EVAL_38),
    ._EVAL_39(out_xbar__EVAL_39),
    ._EVAL_40(out_xbar__EVAL_40),
    ._EVAL_41(out_xbar__EVAL_41),
    ._EVAL_42(out_xbar__EVAL_42),
    ._EVAL_43(out_xbar__EVAL_43),
    ._EVAL_44(out_xbar__EVAL_44),
    ._EVAL_45(out_xbar__EVAL_45),
    ._EVAL_46(out_xbar__EVAL_46),
    ._EVAL_47(out_xbar__EVAL_47),
    ._EVAL_48(out_xbar__EVAL_48),
    ._EVAL_49(out_xbar__EVAL_49),
    ._EVAL_50(out_xbar__EVAL_50),
    ._EVAL_51(out_xbar__EVAL_51),
    ._EVAL_52(out_xbar__EVAL_52),
    ._EVAL_53(out_xbar__EVAL_53),
    ._EVAL_54(out_xbar__EVAL_54),
    ._EVAL_55(out_xbar__EVAL_55),
    ._EVAL_56(out_xbar__EVAL_56),
    ._EVAL_57(out_xbar__EVAL_57),
    ._EVAL_58(out_xbar__EVAL_58),
    ._EVAL_59(out_xbar__EVAL_59),
    ._EVAL_60(out_xbar__EVAL_60),
    ._EVAL_61(out_xbar__EVAL_61),
    ._EVAL_62(out_xbar__EVAL_62),
    ._EVAL_63(out_xbar__EVAL_63),
    ._EVAL_64(out_xbar__EVAL_64),
    ._EVAL_65(out_xbar__EVAL_65),
    ._EVAL_66(out_xbar__EVAL_66),
    ._EVAL_67(out_xbar__EVAL_67),
    ._EVAL_68(out_xbar__EVAL_68),
    ._EVAL_69(out_xbar__EVAL_69),
    ._EVAL_70(out_xbar__EVAL_70),
    ._EVAL_71(out_xbar__EVAL_71),
    ._EVAL_72(out_xbar__EVAL_72),
    ._EVAL_73(out_xbar__EVAL_73),
    ._EVAL_74(out_xbar__EVAL_74),
    ._EVAL_75(out_xbar__EVAL_75),
    ._EVAL_76(out_xbar__EVAL_76),
    ._EVAL_77(out_xbar__EVAL_77),
    ._EVAL_78(out_xbar__EVAL_78),
    ._EVAL_79(out_xbar__EVAL_79),
    ._EVAL_80(out_xbar__EVAL_80),
    ._EVAL_81(out_xbar__EVAL_81),
    ._EVAL_82(out_xbar__EVAL_82),
    ._EVAL_83(out_xbar__EVAL_83),
    ._EVAL_84(out_xbar__EVAL_84),
    ._EVAL_85(out_xbar__EVAL_85),
    ._EVAL_86(out_xbar__EVAL_86),
    ._EVAL_87(out_xbar__EVAL_87),
    ._EVAL_88(out_xbar__EVAL_88),
    ._EVAL_89(out_xbar__EVAL_89),
    ._EVAL_90(out_xbar__EVAL_90),
    ._EVAL_91(out_xbar__EVAL_91),
    ._EVAL_92(out_xbar__EVAL_92),
    ._EVAL_93(out_xbar__EVAL_93),
    ._EVAL_94(out_xbar__EVAL_94),
    ._EVAL_95(out_xbar__EVAL_95),
    ._EVAL_96(out_xbar__EVAL_96),
    ._EVAL_97(out_xbar__EVAL_97),
    ._EVAL_98(out_xbar__EVAL_98),
    ._EVAL_99(out_xbar__EVAL_99),
    ._EVAL_100(out_xbar__EVAL_100),
    ._EVAL_101(out_xbar__EVAL_101),
    ._EVAL_102(out_xbar__EVAL_102),
    ._EVAL_103(out_xbar__EVAL_103),
    ._EVAL_104(out_xbar__EVAL_104),
    ._EVAL_105(out_xbar__EVAL_105),
    ._EVAL_106(out_xbar__EVAL_106),
    ._EVAL_107(out_xbar__EVAL_107),
    ._EVAL_108(out_xbar__EVAL_108),
    ._EVAL_109(out_xbar__EVAL_109),
    ._EVAL_110(out_xbar__EVAL_110),
    ._EVAL_111(out_xbar__EVAL_111),
    ._EVAL_112(out_xbar__EVAL_112),
    ._EVAL_113(out_xbar__EVAL_113),
    ._EVAL_114(out_xbar__EVAL_114),
    ._EVAL_115(out_xbar__EVAL_115)
  );
  _EVAL_82 coupler_to_debug (
    ._EVAL(coupler_to_debug__EVAL),
    ._EVAL_0(coupler_to_debug__EVAL_0),
    ._EVAL_1(coupler_to_debug__EVAL_1),
    ._EVAL_2(coupler_to_debug__EVAL_2),
    ._EVAL_3(coupler_to_debug__EVAL_3),
    ._EVAL_4(coupler_to_debug__EVAL_4),
    ._EVAL_5(coupler_to_debug__EVAL_5),
    ._EVAL_6(coupler_to_debug__EVAL_6),
    ._EVAL_7(coupler_to_debug__EVAL_7),
    ._EVAL_8(coupler_to_debug__EVAL_8),
    ._EVAL_9(coupler_to_debug__EVAL_9),
    ._EVAL_10(coupler_to_debug__EVAL_10),
    ._EVAL_11(coupler_to_debug__EVAL_11),
    ._EVAL_12(coupler_to_debug__EVAL_12),
    ._EVAL_13(coupler_to_debug__EVAL_13),
    ._EVAL_14(coupler_to_debug__EVAL_14),
    ._EVAL_15(coupler_to_debug__EVAL_15),
    ._EVAL_16(coupler_to_debug__EVAL_16),
    ._EVAL_17(coupler_to_debug__EVAL_17),
    ._EVAL_18(coupler_to_debug__EVAL_18),
    ._EVAL_19(coupler_to_debug__EVAL_19),
    ._EVAL_20(coupler_to_debug__EVAL_20),
    ._EVAL_21(coupler_to_debug__EVAL_21),
    ._EVAL_22(coupler_to_debug__EVAL_22),
    ._EVAL_23(coupler_to_debug__EVAL_23),
    ._EVAL_24(coupler_to_debug__EVAL_24),
    ._EVAL_25(coupler_to_debug__EVAL_25),
    ._EVAL_26(coupler_to_debug__EVAL_26),
    ._EVAL_27(coupler_to_debug__EVAL_27),
    ._EVAL_28(coupler_to_debug__EVAL_28),
    ._EVAL_29(coupler_to_debug__EVAL_29),
    ._EVAL_30(coupler_to_debug__EVAL_30),
    ._EVAL_31(coupler_to_debug__EVAL_31),
    ._EVAL_32(coupler_to_debug__EVAL_32)
  );
  _EVAL_57 subsystem_cbus_clock_groups (
    ._EVAL_0(subsystem_cbus_clock_groups__EVAL_0),
    ._EVAL_4(subsystem_cbus_clock_groups__EVAL_4),
    ._EVAL_5(subsystem_cbus_clock_groups__EVAL_5),
    ._EVAL_6(subsystem_cbus_clock_groups__EVAL_6)
  );
  _EVAL_106 buffer_1 (
    ._EVAL(buffer_1__EVAL),
    ._EVAL_0(buffer_1__EVAL_0),
    ._EVAL_1(buffer_1__EVAL_1),
    ._EVAL_2(buffer_1__EVAL_2),
    ._EVAL_3(buffer_1__EVAL_3),
    ._EVAL_4(buffer_1__EVAL_4),
    ._EVAL_5(buffer_1__EVAL_5),
    ._EVAL_6(buffer_1__EVAL_6),
    ._EVAL_7(buffer_1__EVAL_7),
    ._EVAL_8(buffer_1__EVAL_8),
    ._EVAL_9(buffer_1__EVAL_9),
    ._EVAL_10(buffer_1__EVAL_10),
    ._EVAL_11(buffer_1__EVAL_11),
    ._EVAL_12(buffer_1__EVAL_12),
    ._EVAL_13(buffer_1__EVAL_13),
    ._EVAL_14(buffer_1__EVAL_14),
    ._EVAL_15(buffer_1__EVAL_15),
    ._EVAL_16(buffer_1__EVAL_16),
    ._EVAL_17(buffer_1__EVAL_17),
    ._EVAL_18(buffer_1__EVAL_18),
    ._EVAL_19(buffer_1__EVAL_19),
    ._EVAL_20(buffer_1__EVAL_20),
    ._EVAL_21(buffer_1__EVAL_21),
    ._EVAL_22(buffer_1__EVAL_22),
    ._EVAL_23(buffer_1__EVAL_23),
    ._EVAL_24(buffer_1__EVAL_24),
    ._EVAL_25(buffer_1__EVAL_25),
    ._EVAL_26(buffer_1__EVAL_26),
    ._EVAL_27(buffer_1__EVAL_27),
    ._EVAL_28(buffer_1__EVAL_28),
    ._EVAL_29(buffer_1__EVAL_29),
    ._EVAL_30(buffer_1__EVAL_30),
    ._EVAL_31(buffer_1__EVAL_31),
    ._EVAL_32(buffer_1__EVAL_32),
    ._EVAL_33(buffer_1__EVAL_33),
    ._EVAL_34(buffer_1__EVAL_34),
    ._EVAL_35(buffer_1__EVAL_35),
    ._EVAL_36(buffer_1__EVAL_36),
    ._EVAL_37(buffer_1__EVAL_37),
    ._EVAL_38(buffer_1__EVAL_38),
    ._EVAL_39(buffer_1__EVAL_39),
    ._EVAL_40(buffer_1__EVAL_40),
    ._EVAL_41(buffer_1__EVAL_41),
    ._EVAL_42(buffer_1__EVAL_42),
    ._EVAL_43(buffer_1__EVAL_43),
    ._EVAL_44(buffer_1__EVAL_44),
    ._EVAL_45(buffer_1__EVAL_45),
    ._EVAL_46(buffer_1__EVAL_46),
    ._EVAL_47(buffer_1__EVAL_47),
    ._EVAL_48(buffer_1__EVAL_48),
    ._EVAL_49(buffer_1__EVAL_49),
    ._EVAL_50(buffer_1__EVAL_50),
    ._EVAL_51(buffer_1__EVAL_51),
    ._EVAL_52(buffer_1__EVAL_52),
    ._EVAL_53(buffer_1__EVAL_53),
    ._EVAL_54(buffer_1__EVAL_54)
  );
  _EVAL_61 in_xbar (
    ._EVAL(in_xbar__EVAL),
    ._EVAL_0(in_xbar__EVAL_0),
    ._EVAL_1(in_xbar__EVAL_1),
    ._EVAL_2(in_xbar__EVAL_2),
    ._EVAL_3(in_xbar__EVAL_3),
    ._EVAL_4(in_xbar__EVAL_4),
    ._EVAL_5(in_xbar__EVAL_5),
    ._EVAL_6(in_xbar__EVAL_6),
    ._EVAL_7(in_xbar__EVAL_7),
    ._EVAL_8(in_xbar__EVAL_8),
    ._EVAL_9(in_xbar__EVAL_9),
    ._EVAL_10(in_xbar__EVAL_10),
    ._EVAL_11(in_xbar__EVAL_11),
    ._EVAL_12(in_xbar__EVAL_12),
    ._EVAL_13(in_xbar__EVAL_13),
    ._EVAL_14(in_xbar__EVAL_14),
    ._EVAL_15(in_xbar__EVAL_15),
    ._EVAL_16(in_xbar__EVAL_16),
    ._EVAL_17(in_xbar__EVAL_17),
    ._EVAL_18(in_xbar__EVAL_18),
    ._EVAL_19(in_xbar__EVAL_19),
    ._EVAL_20(in_xbar__EVAL_20),
    ._EVAL_21(in_xbar__EVAL_21),
    ._EVAL_22(in_xbar__EVAL_22),
    ._EVAL_23(in_xbar__EVAL_23),
    ._EVAL_24(in_xbar__EVAL_24),
    ._EVAL_25(in_xbar__EVAL_25),
    ._EVAL_26(in_xbar__EVAL_26),
    ._EVAL_27(in_xbar__EVAL_27),
    ._EVAL_28(in_xbar__EVAL_28),
    ._EVAL_29(in_xbar__EVAL_29),
    ._EVAL_30(in_xbar__EVAL_30),
    ._EVAL_31(in_xbar__EVAL_31),
    ._EVAL_32(in_xbar__EVAL_32),
    ._EVAL_33(in_xbar__EVAL_33),
    ._EVAL_34(in_xbar__EVAL_34),
    ._EVAL_35(in_xbar__EVAL_35),
    ._EVAL_36(in_xbar__EVAL_36),
    ._EVAL_37(in_xbar__EVAL_37),
    ._EVAL_38(in_xbar__EVAL_38),
    ._EVAL_39(in_xbar__EVAL_39),
    ._EVAL_40(in_xbar__EVAL_40),
    ._EVAL_41(in_xbar__EVAL_41),
    ._EVAL_42(in_xbar__EVAL_42),
    ._EVAL_43(in_xbar__EVAL_43),
    ._EVAL_44(in_xbar__EVAL_44),
    ._EVAL_45(in_xbar__EVAL_45),
    ._EVAL_46(in_xbar__EVAL_46),
    ._EVAL_47(in_xbar__EVAL_47),
    ._EVAL_48(in_xbar__EVAL_48),
    ._EVAL_49(in_xbar__EVAL_49),
    ._EVAL_50(in_xbar__EVAL_50),
    ._EVAL_51(in_xbar__EVAL_51),
    ._EVAL_52(in_xbar__EVAL_52),
    ._EVAL_53(in_xbar__EVAL_53),
    ._EVAL_54(in_xbar__EVAL_54)
  );
  _EVAL_0 clockGroup (
    ._EVAL(clockGroup__EVAL),
    ._EVAL_0(clockGroup__EVAL_0),
    ._EVAL_1(clockGroup__EVAL_1),
    ._EVAL_2(clockGroup__EVAL_2)
  );
  _EVAL_1 fixedClockNode (
    ._EVAL(fixedClockNode__EVAL),
    ._EVAL_0(fixedClockNode__EVAL_0),
    ._EVAL_1(fixedClockNode__EVAL_1),
    ._EVAL_2(fixedClockNode__EVAL_2)
  );
  _EVAL_69 atomics (
    ._EVAL(atomics__EVAL),
    ._EVAL_0(atomics__EVAL_0),
    ._EVAL_1(atomics__EVAL_1),
    ._EVAL_2(atomics__EVAL_2),
    ._EVAL_3(atomics__EVAL_3),
    ._EVAL_4(atomics__EVAL_4),
    ._EVAL_5(atomics__EVAL_5),
    ._EVAL_6(atomics__EVAL_6),
    ._EVAL_7(atomics__EVAL_7),
    ._EVAL_8(atomics__EVAL_8),
    ._EVAL_9(atomics__EVAL_9),
    ._EVAL_10(atomics__EVAL_10),
    ._EVAL_11(atomics__EVAL_11),
    ._EVAL_12(atomics__EVAL_12),
    ._EVAL_13(atomics__EVAL_13),
    ._EVAL_14(atomics__EVAL_14),
    ._EVAL_15(atomics__EVAL_15),
    ._EVAL_16(atomics__EVAL_16),
    ._EVAL_17(atomics__EVAL_17),
    ._EVAL_18(atomics__EVAL_18),
    ._EVAL_19(atomics__EVAL_19),
    ._EVAL_20(atomics__EVAL_20),
    ._EVAL_21(atomics__EVAL_21),
    ._EVAL_22(atomics__EVAL_22),
    ._EVAL_23(atomics__EVAL_23),
    ._EVAL_24(atomics__EVAL_24),
    ._EVAL_25(atomics__EVAL_25),
    ._EVAL_26(atomics__EVAL_26),
    ._EVAL_27(atomics__EVAL_27),
    ._EVAL_28(atomics__EVAL_28),
    ._EVAL_29(atomics__EVAL_29),
    ._EVAL_30(atomics__EVAL_30),
    ._EVAL_31(atomics__EVAL_31),
    ._EVAL_32(atomics__EVAL_32),
    ._EVAL_33(atomics__EVAL_33),
    ._EVAL_34(atomics__EVAL_34),
    ._EVAL_35(atomics__EVAL_35),
    ._EVAL_36(atomics__EVAL_36),
    ._EVAL_37(atomics__EVAL_37),
    ._EVAL_38(atomics__EVAL_38),
    ._EVAL_39(atomics__EVAL_39),
    ._EVAL_40(atomics__EVAL_40),
    ._EVAL_41(atomics__EVAL_41),
    ._EVAL_42(atomics__EVAL_42),
    ._EVAL_43(atomics__EVAL_43),
    ._EVAL_44(atomics__EVAL_44),
    ._EVAL_45(atomics__EVAL_45),
    ._EVAL_46(atomics__EVAL_46),
    ._EVAL_47(atomics__EVAL_47),
    ._EVAL_48(atomics__EVAL_48),
    ._EVAL_49(atomics__EVAL_49),
    ._EVAL_50(atomics__EVAL_50),
    ._EVAL_51(atomics__EVAL_51)
  );
  _EVAL_59 fixer (
    ._EVAL(fixer__EVAL),
    ._EVAL_0(fixer__EVAL_0),
    ._EVAL_1(fixer__EVAL_1),
    ._EVAL_2(fixer__EVAL_2),
    ._EVAL_3(fixer__EVAL_3),
    ._EVAL_4(fixer__EVAL_4),
    ._EVAL_5(fixer__EVAL_5),
    ._EVAL_6(fixer__EVAL_6),
    ._EVAL_7(fixer__EVAL_7),
    ._EVAL_8(fixer__EVAL_8),
    ._EVAL_9(fixer__EVAL_9),
    ._EVAL_10(fixer__EVAL_10),
    ._EVAL_11(fixer__EVAL_11),
    ._EVAL_12(fixer__EVAL_12),
    ._EVAL_13(fixer__EVAL_13),
    ._EVAL_14(fixer__EVAL_14),
    ._EVAL_15(fixer__EVAL_15),
    ._EVAL_16(fixer__EVAL_16),
    ._EVAL_17(fixer__EVAL_17),
    ._EVAL_18(fixer__EVAL_18),
    ._EVAL_19(fixer__EVAL_19),
    ._EVAL_20(fixer__EVAL_20),
    ._EVAL_21(fixer__EVAL_21),
    ._EVAL_22(fixer__EVAL_22),
    ._EVAL_23(fixer__EVAL_23),
    ._EVAL_24(fixer__EVAL_24),
    ._EVAL_25(fixer__EVAL_25),
    ._EVAL_26(fixer__EVAL_26),
    ._EVAL_27(fixer__EVAL_27),
    ._EVAL_28(fixer__EVAL_28),
    ._EVAL_29(fixer__EVAL_29),
    ._EVAL_30(fixer__EVAL_30),
    ._EVAL_31(fixer__EVAL_31),
    ._EVAL_32(fixer__EVAL_32),
    ._EVAL_33(fixer__EVAL_33),
    ._EVAL_34(fixer__EVAL_34),
    ._EVAL_35(fixer__EVAL_35),
    ._EVAL_36(fixer__EVAL_36),
    ._EVAL_37(fixer__EVAL_37),
    ._EVAL_38(fixer__EVAL_38),
    ._EVAL_39(fixer__EVAL_39),
    ._EVAL_40(fixer__EVAL_40),
    ._EVAL_41(fixer__EVAL_41),
    ._EVAL_42(fixer__EVAL_42),
    ._EVAL_43(fixer__EVAL_43),
    ._EVAL_44(fixer__EVAL_44),
    ._EVAL_45(fixer__EVAL_45),
    ._EVAL_46(fixer__EVAL_46),
    ._EVAL_47(fixer__EVAL_47),
    ._EVAL_48(fixer__EVAL_48)
  );
  assign out_xbar__EVAL_28 = wrapped_error_device__EVAL_10;
  assign fixer__EVAL_14 = out_xbar__EVAL_66;
  assign out_xbar__EVAL_35 = wrapped_error_device__EVAL_2;
  assign _EVAL_60 = buffer_1__EVAL_51;
  assign coupler_to_clic__EVAL_8 = _EVAL_38;
  assign buffer__EVAL_41 = atomics__EVAL_24;
  assign out_xbar__EVAL_114 = coupler_to_clic__EVAL_26;
  assign out_xbar__EVAL_108 = fixer__EVAL_29;
  assign coupler_to_clic__EVAL_6 = out_xbar__EVAL_83;
  assign coupler_to_debug__EVAL = fixedClockNode__EVAL_0;
  assign out_xbar__EVAL_96 = coupler_to_clic__EVAL_14;
  assign coupler_to_debug__EVAL_4 = out_xbar__EVAL_103;
  assign buffer__EVAL_48 = atomics__EVAL_41;
  assign fixer__EVAL_6 = out_xbar__EVAL_6;
  assign buffer__EVAL_23 = atomics__EVAL_40;
  assign atomics__EVAL_18 = in_xbar__EVAL_31;
  assign out_xbar__EVAL_61 = fixer__EVAL_2;
  assign coupler_to_port_named_ahb_periph_port__EVAL = out_xbar__EVAL_94;
  assign atomics__EVAL_14 = in_xbar__EVAL_8;
  assign coupler_to_port_named_ahb_periph_port__EVAL_17 = out_xbar__EVAL;
  assign buffer__EVAL_46 = fixer__EVAL_48;
  assign _EVAL_70 = fixedClockNode__EVAL_0;
  assign out_xbar__EVAL_57 = wrapped_error_device__EVAL_4;
  assign atomics__EVAL_21 = in_xbar__EVAL_34;
  assign coupler_to_clic__EVAL_17 = out_xbar__EVAL_27;
  assign _EVAL_77 = coupler_to_port_named_ahb_periph_port__EVAL_26;
  assign _EVAL_11 = buffer_1__EVAL_10;
  assign out_xbar__EVAL_30 = coupler_to_testIndicator__EVAL_2;
  assign in_xbar__EVAL_40 = buffer_1__EVAL_27;
  assign atomics__EVAL_2 = buffer__EVAL_22;
  assign buffer__EVAL_15 = fixer__EVAL_11;
  assign coupler_to_testIndicator__EVAL_10 = out_xbar__EVAL_64;
  assign out_xbar__EVAL_2 = wrapped_error_device__EVAL_12;
  assign _EVAL_78 = fixedClockNode__EVAL_2;
  assign coupler_to_testIndicator__EVAL_28 = fixedClockNode__EVAL_2;
  assign coupler_to_debug__EVAL_7 = fixedClockNode__EVAL_2;
  assign in_xbar__EVAL_22 = atomics__EVAL_30;
  assign coupler_to_port_named_ahb_periph_port__EVAL_4 = out_xbar__EVAL_48;
  assign fixer__EVAL_16 = buffer__EVAL_40;
  assign atomics__EVAL_5 = in_xbar__EVAL_45;
  assign out_xbar__EVAL_99 = coupler_to_testIndicator__EVAL_18;
  assign atomics__EVAL_13 = in_xbar__EVAL_9;
  assign fixer__EVAL_12 = fixedClockNode__EVAL_2;
  assign coupler_to_testIndicator__EVAL_14 = out_xbar__EVAL_34;
  assign atomics__EVAL_12 = in_xbar__EVAL_5;
  assign in_xbar__EVAL_35 = buffer_1__EVAL_48;
  assign coupler_to_debug__EVAL_0 = out_xbar__EVAL_89;
  assign coupler_to_debug__EVAL_9 = out_xbar__EVAL_109;
  assign wrapped_error_device__EVAL_5 = out_xbar__EVAL_56;
  assign _EVAL_36 = coupler_to_clic__EVAL_12;
  assign atomics__EVAL_9 = in_xbar__EVAL_21;
  assign coupler_to_port_named_ahb_periph_port__EVAL_30 = out_xbar__EVAL_72;
  assign coupler_to_port_named_ahb_periph_port__EVAL_8 = out_xbar__EVAL_0;
  assign coupler_to_testIndicator__EVAL = _EVAL_74;
  assign out_xbar__EVAL_63 = coupler_to_port_named_ahb_periph_port__EVAL_3;
  assign buffer_1__EVAL_17 = _EVAL_69;
  assign buffer_1__EVAL_47 = fixedClockNode__EVAL_2;
  assign in_xbar__EVAL = atomics__EVAL_7;
  assign out_xbar__EVAL_100 = coupler_to_testIndicator__EVAL_15;
  assign buffer__EVAL_31 = fixer__EVAL_9;
  assign out_xbar__EVAL_87 = coupler_to_debug__EVAL_10;
  assign out_xbar__EVAL_86 = fixedClockNode__EVAL_0;
  assign in_xbar__EVAL_28 = fixedClockNode__EVAL_2;
  assign out_xbar__EVAL_95 = fixer__EVAL_28;
  assign out_xbar__EVAL_52 = coupler_to_port_named_ahb_periph_port__EVAL_7;
  assign out_xbar__EVAL_12 = fixer__EVAL_35;
  assign buffer_1__EVAL_35 = _EVAL_80;
  assign buffer_1__EVAL_8 = in_xbar__EVAL_32;
  assign _EVAL_39 = coupler_to_testIndicator__EVAL_0;
  assign out_xbar__EVAL_5 = wrapped_error_device__EVAL_19;
  assign coupler_to_clic__EVAL_9 = out_xbar__EVAL_32;
  assign fixer__EVAL_3 = buffer__EVAL_47;
  assign _EVAL_27 = buffer_1__EVAL_14;
  assign wrapped_error_device__EVAL_18 = out_xbar__EVAL_65;
  assign coupler_to_testIndicator__EVAL_20 = out_xbar__EVAL_68;
  assign out_xbar__EVAL_90 = fixer__EVAL_17;
  assign out_xbar__EVAL_71 = coupler_to_debug__EVAL_29;
  assign out_xbar__EVAL_73 = coupler_to_debug__EVAL_25;
  assign coupler_to_clic__EVAL_1 = out_xbar__EVAL_24;
  assign _EVAL_82 = coupler_to_debug__EVAL_1;
  assign out_xbar__EVAL_107 = wrapped_error_device__EVAL_7;
  assign out_xbar__EVAL_98 = coupler_to_debug__EVAL_15;
  assign out_xbar__EVAL_19 = coupler_to_clic__EVAL_23;
  assign buffer_1__EVAL_7 = in_xbar__EVAL_49;
  assign fixer__EVAL_30 = buffer__EVAL_25;
  assign coupler_to_port_named_ahb_periph_port__EVAL_5 = out_xbar__EVAL_23;
  assign coupler_to_clic__EVAL_7 = fixedClockNode__EVAL_0;
  assign out_xbar__EVAL_45 = coupler_to_port_named_ahb_periph_port__EVAL_29;
  assign buffer__EVAL_16 = atomics__EVAL_48;
  assign _EVAL_18 = coupler_to_debug__EVAL_22;
  assign out_xbar__EVAL_37 = wrapped_error_device__EVAL_15;
  assign out_xbar__EVAL_110 = fixer__EVAL_39;
  assign atomics__EVAL_39 = in_xbar__EVAL_51;
  assign wrapped_error_device__EVAL_9 = out_xbar__EVAL_15;
  assign buffer_1__EVAL_2 = _EVAL_12;
  assign coupler_to_testIndicator__EVAL_19 = out_xbar__EVAL_59;
  assign coupler_to_debug__EVAL_19 = _EVAL_3;
  assign coupler_to_testIndicator__EVAL_31 = out_xbar__EVAL_18;
  assign wrapped_error_device__EVAL_8 = fixedClockNode__EVAL_0;
  assign in_xbar__EVAL_20 = buffer_1__EVAL_53;
  assign atomics__EVAL_35 = in_xbar__EVAL_15;
  assign _EVAL_65 = coupler_to_clic__EVAL_28;
  assign atomics__EVAL_45 = buffer__EVAL_27;
  assign atomics__EVAL_31 = in_xbar__EVAL_52;
  assign buffer_1__EVAL_4 = _EVAL_35;
  assign coupler_to_debug__EVAL_31 = _EVAL_54;
  assign out_xbar__EVAL_104 = wrapped_error_device__EVAL_16;
  assign atomics__EVAL_8 = buffer__EVAL_34;
  assign _EVAL_21 = coupler_to_testIndicator__EVAL_21;
  assign out_xbar__EVAL_58 = coupler_to_port_named_ahb_periph_port__EVAL_19;
  assign atomics__EVAL_0 = buffer__EVAL_44;
  assign buffer_1__EVAL_19 = _EVAL_62;
  assign buffer_1__EVAL_25 = in_xbar__EVAL_44;
  assign wrapped_error_device__EVAL_14 = out_xbar__EVAL_115;
  assign in_xbar__EVAL_7 = buffer_1__EVAL_21;
  assign _EVAL_8 = coupler_to_testIndicator__EVAL_23;
  assign out_xbar__EVAL_21 = coupler_to_port_named_ahb_periph_port__EVAL_21;
  assign fixer__EVAL_13 = out_xbar__EVAL_38;
  assign coupler_to_debug__EVAL_6 = out_xbar__EVAL_67;
  assign in_xbar__EVAL_14 = buffer_1__EVAL_5;
  assign buffer_1__EVAL_52 = _EVAL_49;
  assign _EVAL_44 = coupler_to_clic__EVAL;
  assign fixer__EVAL_37 = fixedClockNode__EVAL_0;
  assign atomics__EVAL_19 = buffer__EVAL_13;
  assign buffer_1__EVAL_33 = in_xbar__EVAL_50;
  assign coupler_to_clic__EVAL_22 = out_xbar__EVAL_85;
  assign _EVAL_52 = buffer_1__EVAL_54;
  assign _EVAL_13 = coupler_to_port_named_ahb_periph_port__EVAL_13;
  assign out_xbar__EVAL_39 = fixer__EVAL_45;
  assign coupler_to_port_named_ahb_periph_port__EVAL_31 = out_xbar__EVAL_54;
  assign _EVAL_64 = coupler_to_testIndicator__EVAL_27;
  assign buffer__EVAL_0 = fixer__EVAL_25;
  assign fixer__EVAL_18 = out_xbar__EVAL_69;
  assign coupler_to_port_named_ahb_periph_port__EVAL_18 = out_xbar__EVAL_33;
  assign fixer__EVAL_32 = buffer__EVAL_8;
  assign coupler_to_port_named_ahb_periph_port__EVAL_0 = _EVAL_88;
  assign in_xbar__EVAL_37 = buffer_1__EVAL_41;
  assign clockGroup__EVAL = subsystem_cbus_clock_groups__EVAL_0;
  assign in_xbar__EVAL_6 = buffer_1__EVAL_1;
  assign coupler_to_clic__EVAL_24 = _EVAL_17;
  assign atomics__EVAL_34 = fixedClockNode__EVAL_2;
  assign buffer__EVAL_43 = fixedClockNode__EVAL_0;
  assign out_xbar__EVAL_101 = coupler_to_port_named_ahb_periph_port__EVAL_20;
  assign atomics__EVAL_42 = fixedClockNode__EVAL_0;
  assign coupler_to_debug__EVAL_28 = _EVAL;
  assign atomics__EVAL_27 = in_xbar__EVAL_13;
  assign buffer_1__EVAL_43 = _EVAL_66;
  assign out_xbar__EVAL_22 = fixer__EVAL_34;
  assign atomics__EVAL_44 = buffer__EVAL_26;
  assign coupler_to_clic__EVAL_15 = fixedClockNode__EVAL_2;
  assign fixer__EVAL_0 = buffer__EVAL_38;
  assign atomics__EVAL_49 = buffer__EVAL_3;
  assign in_xbar__EVAL_36 = atomics__EVAL_10;
  assign _EVAL_31 = coupler_to_testIndicator__EVAL_24;
  assign atomics__EVAL_46 = buffer__EVAL_9;
  assign in_xbar__EVAL_42 = buffer_1__EVAL_36;
  assign out_xbar__EVAL_60 = fixer__EVAL_7;
  assign coupler_to_debug__EVAL_23 = out_xbar__EVAL_51;
  assign fixer__EVAL_8 = out_xbar__EVAL_44;
  assign out_xbar__EVAL_11 = coupler_to_port_named_ahb_periph_port__EVAL_10;
  assign out_xbar__EVAL_36 = fixer__EVAL_4;
  assign _EVAL_32 = coupler_to_clic__EVAL_25;
  assign _EVAL_29 = buffer_1__EVAL_23;
  assign coupler_to_testIndicator__EVAL_11 = out_xbar__EVAL_84;
  assign fixer__EVAL_41 = buffer__EVAL_11;
  assign _EVAL_76 = coupler_to_clic__EVAL_0;
  assign coupler_to_port_named_ahb_periph_port__EVAL_32 = out_xbar__EVAL_31;
  assign buffer_1__EVAL_9 = in_xbar__EVAL_18;
  assign atomics__EVAL_32 = in_xbar__EVAL_12;
  assign buffer__EVAL_2 = atomics__EVAL_47;
  assign out_xbar__EVAL_55 = coupler_to_debug__EVAL_26;
  assign wrapped_error_device__EVAL_13 = out_xbar__EVAL_111;
  assign buffer__EVAL_19 = atomics__EVAL_22;
  assign coupler_to_clic__EVAL_20 = out_xbar__EVAL_4;
  assign buffer_1__EVAL_32 = in_xbar__EVAL_30;
  assign buffer__EVAL_18 = fixer__EVAL_1;
  assign in_xbar__EVAL_48 = buffer_1__EVAL_24;
  assign _EVAL_90 = coupler_to_clic__EVAL_4;
  assign fixedClockNode__EVAL = clockGroup__EVAL_1;
  assign coupler_to_port_named_ahb_periph_port__EVAL_11 = fixedClockNode__EVAL_2;
  assign buffer__EVAL_36 = atomics__EVAL_50;
  assign _EVAL_68 = coupler_to_clic__EVAL_30;
  assign buffer_1__EVAL_16 = _EVAL_14;
  assign buffer_1__EVAL_20 = _EVAL_0;
  assign out_xbar__EVAL_77 = coupler_to_clic__EVAL_13;
  assign _EVAL_45 = buffer_1__EVAL_34;
  assign coupler_to_clic__EVAL_2 = out_xbar__EVAL_13;
  assign coupler_to_debug__EVAL_2 = out_xbar__EVAL_26;
  assign out_xbar__EVAL_14 = coupler_to_clic__EVAL_3;
  assign _EVAL_28 = coupler_to_debug__EVAL_24;
  assign in_xbar__EVAL_19 = buffer_1__EVAL_39;
  assign in_xbar__EVAL_25 = atomics__EVAL;
  assign out_xbar__EVAL_17 = wrapped_error_device__EVAL_17;
  assign coupler_to_clic__EVAL_29 = _EVAL_7;
  assign _EVAL_30 = coupler_to_debug__EVAL_13;
  assign in_xbar__EVAL_38 = atomics__EVAL_26;
  assign coupler_to_testIndicator__EVAL_22 = _EVAL_15;
  assign in_xbar__EVAL_39 = buffer_1__EVAL;
  assign _EVAL_20 = coupler_to_testIndicator__EVAL_9;
  assign buffer_1__EVAL_18 = _EVAL_59;
  assign buffer__EVAL_4 = atomics__EVAL_16;
  assign out_xbar__EVAL_79 = fixedClockNode__EVAL_2;
  assign _EVAL_26 = coupler_to_testIndicator__EVAL_3;
  assign wrapped_error_device__EVAL_0 = out_xbar__EVAL_9;
  assign coupler_to_testIndicator__EVAL_29 = out_xbar__EVAL_75;
  assign coupler_to_debug__EVAL_17 = _EVAL_34;
  assign coupler_to_testIndicator__EVAL_5 = out_xbar__EVAL_97;
  assign buffer_1__EVAL_22 = _EVAL_63;
  assign in_xbar__EVAL_16 = atomics__EVAL_4;
  assign fixer__EVAL_38 = buffer__EVAL_10;
  assign atomics__EVAL_28 = buffer__EVAL_21;
  assign buffer_1__EVAL_6 = fixedClockNode__EVAL_0;
  assign atomics__EVAL_43 = in_xbar__EVAL_43;
  assign buffer__EVAL_17 = atomics__EVAL_36;
  assign wrapped_error_device__EVAL = fixedClockNode__EVAL_2;
  assign atomics__EVAL_6 = in_xbar__EVAL_33;
  assign buffer_1__EVAL_29 = _EVAL_50;
  assign in_xbar__EVAL_29 = buffer_1__EVAL_12;
  assign fixer__EVAL_10 = out_xbar__EVAL_74;
  assign coupler_to_clic__EVAL_16 = _EVAL_89;
  assign coupler_to_port_named_ahb_periph_port__EVAL_24 = out_xbar__EVAL_76;
  assign buffer__EVAL_1 = atomics__EVAL_15;
  assign _EVAL_22 = coupler_to_debug__EVAL_27;
  assign coupler_to_clic__EVAL_10 = out_xbar__EVAL_113;
  assign buffer__EVAL = fixer__EVAL_47;
  assign wrapped_error_device__EVAL_3 = out_xbar__EVAL_47;
  assign fixer__EVAL_42 = buffer__EVAL_20;
  assign _EVAL_46 = coupler_to_clic__EVAL_18;
  assign wrapped_error_device__EVAL_6 = out_xbar__EVAL_25;
  assign buffer__EVAL_45 = fixer__EVAL_26;
  assign coupler_to_debug__EVAL_14 = out_xbar__EVAL_88;
  assign coupler_to_port_named_ahb_periph_port__EVAL_6 = out_xbar__EVAL_82;
  assign coupler_to_debug__EVAL_5 = _EVAL_75;
  assign fixer__EVAL_23 = buffer__EVAL_14;
  assign buffer_1__EVAL_49 = _EVAL_40;
  assign coupler_to_clic__EVAL_19 = _EVAL_42;
  assign _EVAL_73 = coupler_to_debug__EVAL_8;
  assign in_xbar__EVAL_26 = atomics__EVAL_29;
  assign fixer__EVAL = buffer__EVAL_39;
  assign in_xbar__EVAL_4 = buffer_1__EVAL_11;
  assign out_xbar__EVAL_3 = wrapped_error_device__EVAL_1;
  assign in_xbar__EVAL_47 = buffer_1__EVAL_40;
  assign buffer_1__EVAL_46 = _EVAL_23;
  assign in_xbar__EVAL_27 = atomics__EVAL_1;
  assign coupler_to_port_named_ahb_periph_port__EVAL_12 = _EVAL_84;
  assign _EVAL_24 = buffer_1__EVAL_42;
  assign coupler_to_testIndicator__EVAL_26 = _EVAL_41;
  assign in_xbar__EVAL_2 = atomics__EVAL_11;
  assign coupler_to_clic__EVAL_27 = out_xbar__EVAL_93;
  assign out_xbar__EVAL_40 = fixer__EVAL_15;
  assign out_xbar__EVAL_91 = coupler_to_port_named_ahb_periph_port__EVAL_22;
  assign fixer__EVAL_33 = out_xbar__EVAL_50;
  assign fixer__EVAL_44 = buffer__EVAL_24;
  assign coupler_to_debug__EVAL_32 = out_xbar__EVAL_105;
  assign buffer_1__EVAL_28 = _EVAL_4;
  assign coupler_to_testIndicator__EVAL_6 = fixedClockNode__EVAL_0;
  assign atomics__EVAL_51 = in_xbar__EVAL_41;
  assign _EVAL_2 = coupler_to_testIndicator__EVAL_16;
  assign fixer__EVAL_27 = buffer__EVAL_35;
  assign _EVAL_51 = coupler_to_debug__EVAL_16;
  assign _EVAL_47 = coupler_to_debug__EVAL_18;
  assign coupler_to_clic__EVAL_21 = out_xbar__EVAL_49;
  assign fixer__EVAL_40 = out_xbar__EVAL_10;
  assign clockGroup__EVAL_2 = subsystem_cbus_clock_groups__EVAL_5;
  assign _EVAL_87 = coupler_to_debug__EVAL_12;
  assign out_xbar__EVAL_8 = coupler_to_testIndicator__EVAL_32;
  assign out_xbar__EVAL_70 = fixer__EVAL_20;
  assign coupler_to_testIndicator__EVAL_25 = out_xbar__EVAL_78;
  assign buffer__EVAL_30 = atomics__EVAL_38;
  assign buffer__EVAL_7 = fixer__EVAL_24;
  assign coupler_to_debug__EVAL_20 = out_xbar__EVAL_92;
  assign _EVAL_25 = coupler_to_port_named_ahb_periph_port__EVAL_28;
  assign fixedClockNode__EVAL_1 = clockGroup__EVAL_0;
  assign coupler_to_testIndicator__EVAL_8 = _EVAL_83;
  assign buffer__EVAL_29 = fixer__EVAL_21;
  assign buffer__EVAL_32 = fixedClockNode__EVAL_2;
  assign in_xbar__EVAL_10 = buffer_1__EVAL_44;
  assign _EVAL_72 = coupler_to_port_named_ahb_periph_port__EVAL_9;
  assign in_xbar__EVAL_0 = buffer_1__EVAL_45;
  assign coupler_to_port_named_ahb_periph_port__EVAL_33 = fixedClockNode__EVAL_0;
  assign buffer__EVAL_12 = atomics__EVAL_17;
  assign in_xbar__EVAL_17 = buffer_1__EVAL_15;
  assign _EVAL_79 = coupler_to_port_named_ahb_periph_port__EVAL_27;
  assign coupler_to_port_named_ahb_periph_port__EVAL_15 = _EVAL_10;
  assign atomics__EVAL_3 = buffer__EVAL_42;
  assign wrapped_error_device__EVAL_11 = out_xbar__EVAL_42;
  assign out_xbar__EVAL_20 = fixer__EVAL_36;
  assign fixer__EVAL_22 = out_xbar__EVAL_112;
  assign atomics__EVAL_20 = in_xbar__EVAL_46;
  assign subsystem_cbus_clock_groups__EVAL_6 = _EVAL_16;
  assign coupler_to_debug__EVAL_11 = out_xbar__EVAL_102;
  assign in_xbar__EVAL_11 = fixedClockNode__EVAL_0;
  assign buffer_1__EVAL_31 = in_xbar__EVAL_53;
  assign _EVAL_56 = buffer_1__EVAL_37;
  assign coupler_to_testIndicator__EVAL_7 = _EVAL_57;
  assign out_xbar__EVAL_62 = coupler_to_testIndicator__EVAL_12;
  assign fixer__EVAL_19 = buffer__EVAL_33;
  assign _EVAL_85 = coupler_to_port_named_ahb_periph_port__EVAL_2;
  assign _EVAL_37 = buffer_1__EVAL_13;
  assign buffer_1__EVAL_0 = in_xbar__EVAL_3;
  assign subsystem_cbus_clock_groups__EVAL_4 = _EVAL_43;
  assign out_xbar__EVAL_106 = coupler_to_port_named_ahb_periph_port__EVAL_14;
  assign coupler_to_port_named_ahb_periph_port__EVAL_16 = out_xbar__EVAL_29;
  assign _EVAL_1 = coupler_to_clic__EVAL_5;
  assign out_xbar__EVAL_80 = coupler_to_testIndicator__EVAL_17;
  assign out_xbar__EVAL_7 = fixer__EVAL_43;
  assign buffer__EVAL_5 = atomics__EVAL_33;
  assign buffer_1__EVAL_50 = in_xbar__EVAL_1;
  assign out_xbar__EVAL_46 = coupler_to_debug__EVAL_30;
  assign _EVAL_58 = coupler_to_debug__EVAL_3;
  assign _EVAL_71 = coupler_to_testIndicator__EVAL_1;
  assign fixer__EVAL_31 = buffer__EVAL_28;
  assign in_xbar__EVAL_54 = atomics__EVAL_23;
  assign coupler_to_testIndicator__EVAL_4 = _EVAL_9;
  assign coupler_to_debug__EVAL_21 = _EVAL_19;
  assign coupler_to_testIndicator__EVAL_13 = out_xbar__EVAL_43;
  assign buffer__EVAL_37 = atomics__EVAL_25;
  assign buffer_1__EVAL_3 = in_xbar__EVAL_24;
  assign buffer_1__EVAL_38 = _EVAL_61;
  assign buffer__EVAL_6 = fixer__EVAL_5;
  assign out_xbar__EVAL_1 = coupler_to_port_named_ahb_periph_port__EVAL_25;
  assign buffer_1__EVAL_30 = _EVAL_67;
  assign out_xbar__EVAL_53 = coupler_to_clic__EVAL_11;
  assign _EVAL_86 = coupler_to_clic__EVAL_31;
  assign atomics__EVAL_37 = in_xbar__EVAL_23;
  assign fixer__EVAL_46 = out_xbar__EVAL_81;
  assign coupler_to_port_named_ahb_periph_port__EVAL_1 = out_xbar__EVAL_41;
  assign _EVAL_81 = coupler_to_testIndicator__EVAL_30;
  assign coupler_to_port_named_ahb_periph_port__EVAL_23 = out_xbar__EVAL_16;
  assign coupler_to_clic__EVAL_32 = _EVAL_48;
  assign _EVAL_55 = buffer_1__EVAL_26;
endmodule
