//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_28(
  input  [2:0]  _EVAL,
  output [1:0]  _EVAL_0,
  output [2:0]  _EVAL_1,
  input  [3:0]  _EVAL_2,
  output        _EVAL_3,
  output [30:0] _EVAL_4,
  input         _EVAL_5,
  output [3:0]  _EVAL_6,
  output        _EVAL_7,
  input  [2:0]  _EVAL_8,
  output [2:0]  _EVAL_9,
  output        _EVAL_10,
  output        _EVAL_11,
  input         _EVAL_12,
  output        _EVAL_13,
  output        _EVAL_14,
  input  [1:0]  _EVAL_15,
  output [31:0] _EVAL_16,
  input         _EVAL_17,
  input  [30:0] _EVAL_18,
  output        _EVAL_19,
  input  [31:0] _EVAL_20,
  input         _EVAL_21,
  output [2:0]  _EVAL_22,
  input  [2:0]  _EVAL_23,
  input  [2:0]  _EVAL_24,
  input         _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  output [2:0]  _EVAL_28,
  input  [2:0]  _EVAL_29,
  output [2:0]  _EVAL_30,
  input  [2:0]  _EVAL_31,
  input         _EVAL_32,
  output [2:0]  _EVAL_33,
  output        _EVAL_34,
  output [31:0] _EVAL_35,
  output        _EVAL_36,
  input         _EVAL_37,
  input         _EVAL_38,
  input  [31:0] _EVAL_39,
  input  [2:0]  _EVAL_40,
  output        _EVAL_41,
  input         _EVAL_42,
  output        _EVAL_43,
  input         _EVAL_44,
  input         _EVAL_45,
  output        _EVAL_46,
  input         _EVAL_47,
  output [2:0]  _EVAL_48
);
  assign _EVAL_4 = _EVAL_18;
  assign _EVAL_11 = _EVAL_32;
  assign _EVAL_46 = _EVAL_45;
  assign _EVAL_22 = _EVAL_31;
  assign _EVAL_34 = _EVAL_12;
  assign _EVAL_10 = _EVAL_26;
  assign _EVAL_7 = _EVAL_42;
  assign _EVAL_28 = _EVAL_29;
  assign _EVAL_48 = _EVAL_8;
  assign _EVAL_43 = _EVAL_5;
  assign _EVAL_30 = _EVAL_40;
  assign _EVAL_13 = _EVAL_17;
  assign _EVAL_33 = _EVAL_23;
  assign _EVAL_0 = _EVAL_15;
  assign _EVAL_14 = _EVAL_38;
  assign _EVAL_3 = _EVAL_25;
  assign _EVAL_35 = _EVAL_39;
  assign _EVAL_16 = _EVAL_20;
  assign _EVAL_41 = _EVAL_27;
  assign _EVAL_9 = _EVAL;
  assign _EVAL_1 = _EVAL_24;
  assign _EVAL_19 = _EVAL_21;
  assign _EVAL_6 = _EVAL_2;
  assign _EVAL_36 = _EVAL_47;
endmodule
