//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_40_assert(
  input  [3:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input  [3:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [1:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input  [3:0]  _EVAL_15,
  input  [2:0]  _EVAL_16,
  input  [31:0] _EVAL_17
);
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  reg [2:0] _EVAL_22;
  reg [31:0] _RAND_0;
  wire [32:0] _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire [6:0] _EVAL_39;
  wire [32:0] _EVAL_40;
  wire  _EVAL_41;
  wire [7:0] _EVAL_42;
  wire [1:0] _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire [5:0] _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_61;
  wire  _EVAL_63;
  reg [5:0] _EVAL_64;
  reg [31:0] _RAND_1;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire [32:0] _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  reg  _EVAL_77;
  reg [31:0] _RAND_2;
  reg [31:0] _EVAL_78;
  reg [31:0] _RAND_3;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire [6:0] _EVAL_83;
  wire  _EVAL_84;
  wire [32:0] _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire [1:0] _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  reg [5:0] _EVAL_94;
  reg [31:0] _RAND_4;
  wire [31:0] _EVAL_95;
  wire  _EVAL_96;
  wire [32:0] _EVAL_97;
  wire [5:0] _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_103;
  wire [32:0] _EVAL_104;
  wire [32:0] _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire [32:0] _EVAL_114;
  wire  _EVAL_115;
  wire [1:0] _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire [1:0] _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire [5:0] _EVAL_138;
  wire  _EVAL_139;
  wire [1:0] _EVAL_140;
  wire  _EVAL_141;
  wire [31:0] _EVAL_142;
  wire  _EVAL_143;
  reg [5:0] _EVAL_144;
  reg [31:0] _RAND_5;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire [32:0] _EVAL_153;
  reg [2:0] _EVAL_154;
  reg [31:0] _RAND_6;
  wire  _EVAL_155;
  wire  _EVAL_156;
  reg  _EVAL_157;
  reg [31:0] _RAND_7;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire [31:0] _EVAL_165;
  wire  _EVAL_166;
  wire [6:0] _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire [3:0] _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  reg [1:0] _EVAL_181;
  reg [31:0] _RAND_8;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  reg [31:0] _EVAL_185;
  reg [31:0] _RAND_9;
  reg  _EVAL_186;
  reg [31:0] _RAND_10;
  wire [31:0] _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_195;
  wire [32:0] _EVAL_196;
  wire  _EVAL_197;
  wire [32:0] _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire [32:0] _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire [32:0] _EVAL_209;
  wire  _EVAL_210;
  wire [32:0] _EVAL_211;
  wire  _EVAL_212;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire [5:0] _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire [6:0] _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  reg [5:0] _EVAL_226;
  reg [31:0] _RAND_11;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  reg [3:0] _EVAL_230;
  reg [31:0] _RAND_12;
  wire  _EVAL_231;
  wire [5:0] _EVAL_232;
  wire  _EVAL_233;
  wire [7:0] _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire [31:0] _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire [32:0] _EVAL_249;
  wire [32:0] _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire [5:0] _EVAL_256;
  wire [22:0] _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire [31:0] _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire [32:0] _EVAL_265;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire [3:0] _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire [32:0] _EVAL_276;
  wire  _EVAL_277;
  reg  _EVAL_278;
  reg [31:0] _RAND_13;
  wire [31:0] _EVAL_279;
  wire [7:0] _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire [32:0] _EVAL_283;
  wire  _EVAL_284;
  wire [22:0] _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire [3:0] _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire [3:0] _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  reg [2:0] _EVAL_303;
  reg [31:0] _RAND_14;
  reg [3:0] _EVAL_304;
  reg [31:0] _RAND_15;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire [31:0] _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire [7:0] _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire  _EVAL_318;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_159 = _EVAL_20 | _EVAL_79;
  assign _EVAL_67 = _EVAL_1 & _EVAL_238;
  assign _EVAL_106 = ~_EVAL_210;
  assign _EVAL_241 = _EVAL_78 < plusarg_reader_out;
  assign _EVAL_305 = _EVAL_5 == _EVAL_186;
  assign _EVAL_28 = ~_EVAL_9;
  assign _EVAL_155 = ~_EVAL_222;
  assign _EVAL_316 = ~_EVAL_126;
  assign _EVAL_129 = ~_EVAL_133;
  assign _EVAL_135 = _EVAL_6 == _EVAL_304;
  assign _EVAL_237 = _EVAL_114[31:0];
  assign _EVAL_92 = _EVAL_12 & _EVAL_93;
  assign _EVAL_296 = _EVAL_11 == _EVAL_181;
  assign _EVAL_252 = _EVAL_6 <= 4'h8;
  assign _EVAL_101 = _EVAL_212 & _EVAL_37;
  assign _EVAL_136 = _EVAL_65 | _EVAL_301;
  assign _EVAL_143 = _EVAL_49 | _EVAL_7;
  assign _EVAL_163 = _EVAL_291 & _EVAL_50;
  assign _EVAL_158 = _EVAL_292 | _EVAL_7;
  assign _EVAL_262 = ~_EVAL_169;
  assign _EVAL_85 = $signed(_EVAL_40) & -33'sh1000;
  assign _EVAL_299 = _EVAL_15 >= 4'h2;
  assign _EVAL_285 = 23'hff << _EVAL_15;
  assign _EVAL_114 = _EVAL_78 + 32'h1;
  assign _EVAL_283 = _EVAL_265;
  assign _EVAL_27 = _EVAL_172 | _EVAL_7;
  assign _EVAL_81 = _EVAL_16 <= 3'h2;
  assign _EVAL_91 = _EVAL_4 == 3'h5;
  assign _EVAL_59 = ~_EVAL_195;
  assign _EVAL_240 = _EVAL_247 | _EVAL_7;
  assign _EVAL_187 = _EVAL_17 ^ 32'h40000000;
  assign _EVAL_76 = _EVAL_157 | _EVAL_32;
  assign _EVAL_39 = _EVAL_226 - 6'h1;
  assign _EVAL_195 = _EVAL_299 | _EVAL_7;
  assign _EVAL_258 = ~_EVAL_127;
  assign _EVAL_300 = _EVAL & _EVAL_171;
  assign _EVAL_41 = _EVAL_10 == _EVAL_22;
  assign _EVAL_317 = _EVAL_318 | _EVAL_7;
  assign _EVAL_95 = _EVAL_17 ^ 32'h3000;
  assign _EVAL_232 = _EVAL_39[5:0];
  assign _EVAL_63 = _EVAL_191 | _EVAL_26;
  assign _EVAL_147 = ~_EVAL_54;
  assign _EVAL_118 = $signed(_EVAL_250) == 33'sh0;
  assign _EVAL_287 = ~_EVAL_53;
  assign _EVAL_88 = _EVAL_113 | _EVAL_7;
  assign _EVAL_236 = _EVAL_245 | _EVAL_86;
  assign _EVAL_115 = _EVAL == _EVAL_295;
  assign _EVAL_32 = _EVAL_116[0];
  assign _EVAL_52 = _EVAL_42[7:2];
  assign _EVAL_24 = ~_EVAL_72;
  assign _EVAL_166 = _EVAL_66 | _EVAL_7;
  assign _EVAL_288 = ~_EVAL_25;
  assign _EVAL_105 = $signed(_EVAL_23) & -33'sh1000000;
  assign _EVAL_200 = _EVAL_16 <= 3'h1;
  assign _EVAL_233 = _EVAL_12 & _EVAL_213;
  assign _EVAL_295 = {_EVAL_19,_EVAL_36,_EVAL_89,_EVAL_145};
  assign _EVAL_112 = _EVAL_229 & _EVAL_152;
  assign _EVAL_55 = ~_EVAL_74;
  assign _EVAL_87 = _EVAL_2 == _EVAL_77;
  assign _EVAL_73 = _EVAL_251 | _EVAL_96;
  assign _EVAL_178 = _EVAL_11 != 2'h2;
  assign _EVAL_89 = _EVAL_297 | _EVAL_273;
  assign _EVAL_93 = _EVAL_10 == 3'h5;
  assign _EVAL_34 = _EVAL_11 <= 2'h2;
  assign _EVAL_213 = _EVAL_10 == 3'h1;
  assign _EVAL_248 = _EVAL_10 == 3'h4;
  assign _EVAL_110 = _EVAL_45 | _EVAL_30;
  assign _EVAL_311 = _EVAL_17 ^ 32'h80000000;
  assign _EVAL_255 = $signed(_EVAL_196) == 33'sh0;
  assign _EVAL_293 = _EVAL_189 | _EVAL_7;
  assign _EVAL_142 = _EVAL_17 ^ 32'h2000000;
  assign _EVAL_231 = ~_EVAL_306;
  assign _EVAL_204 = _EVAL_4 <= 3'h6;
  assign _EVAL_275 = ~_EVAL_120;
  assign _EVAL_145 = _EVAL_297 | _EVAL_131;
  assign _EVAL_188 = _EVAL_41 | _EVAL_7;
  assign _EVAL_123 = _EVAL_212 & _EVAL_50;
  assign _EVAL_160 = ~_EVAL_2;
  assign _EVAL_308 = _EVAL_251 & _EVAL_312;
  assign _EVAL_251 = _EVAL_8 & _EVAL_12;
  assign _EVAL_301 = $signed(_EVAL_283) == 33'sh0;
  assign _EVAL_72 = _EVAL_236 | _EVAL_7;
  assign _EVAL_180 = _EVAL_260 == 32'h0;
  assign _EVAL_235 = _EVAL_10[2];
  assign _EVAL_40 = {1'b0,$signed(_EVAL_95)};
  assign _EVAL_18 = ~_EVAL_70;
  assign _EVAL_315 = _EVAL_4[0];
  assign _EVAL_210 = _EVAL_226 == 6'h0;
  assign _EVAL_42 = ~_EVAL_314;
  assign _EVAL_221 = _EVAL_81 | _EVAL_7;
  assign _EVAL_257 = 23'hff << _EVAL_6;
  assign _EVAL_193 = ~_EVAL_0;
  assign _EVAL_314 = _EVAL_285[7:0];
  assign _EVAL_268 = _EVAL_16 <= 3'h4;
  assign _EVAL_30 = _EVAL_44 & _EVAL_118;
  assign _EVAL_273 = _EVAL_229 & _EVAL_101;
  assign _EVAL_208 = _EVAL_298 | _EVAL_7;
  assign _EVAL_250 = _EVAL_249;
  assign _EVAL_58 = ~_EVAL_310;
  assign _EVAL_47 = ~_EVAL_177;
  assign _EVAL_98 = _EVAL_220[5:0];
  assign _EVAL_107 = _EVAL_28 | _EVAL_7;
  assign _EVAL_310 = _EVAL_242 | _EVAL_7;
  assign _EVAL_126 = _EVAL_64 == 6'h0;
  assign _EVAL_131 = _EVAL_229 & _EVAL_123;
  assign _EVAL_54 = _EVAL_178 | _EVAL_7;
  assign _EVAL_234 = _EVAL_257[7:0];
  assign _EVAL_74 = _EVAL_263 | _EVAL_7;
  assign _EVAL_83 = _EVAL_64 - 6'h1;
  assign _EVAL_103 = ~_EVAL_143;
  assign _EVAL_265 = $signed(_EVAL_201) & -33'sh2000;
  assign _EVAL_247 = _EVAL_16 == _EVAL_154;
  assign _EVAL_23 = {1'b0,$signed(_EVAL_142)};
  assign _EVAL_290 = _EVAL_1 & _EVAL_289;
  assign _EVAL_214 = _EVAL_170 | _EVAL_7;
  assign _EVAL_139 = _EVAL_160 | _EVAL_9;
  assign _EVAL_149 = _EVAL_1 & _EVAL_134;
  assign _EVAL_223 = _EVAL_229 & _EVAL_163;
  assign _EVAL_165 = {{24'd0}, _EVAL_280};
  assign _EVAL_242 = _EVAL_110 | _EVAL_79;
  assign _EVAL_171 = ~_EVAL_295;
  assign _EVAL_31 = ~_EVAL_221;
  assign _EVAL_267 = _EVAL_10 == 3'h3;
  assign _EVAL_238 = _EVAL_4 == 3'h4;
  assign _EVAL_199 = _EVAL_307 | _EVAL_272;
  assign _EVAL_51 = ~_EVAL_158;
  assign _EVAL_100 = ~_EVAL_128;
  assign _EVAL_121 = _EVAL_12 & _EVAL_259;
  assign _EVAL_134 = _EVAL_4 == 3'h1;
  assign _EVAL_82 = _EVAL_4 == 3'h2;
  assign _EVAL_280 = ~_EVAL_234;
  assign _EVAL_56 = _EVAL_30 | _EVAL_79;
  assign _EVAL_281 = _EVAL_140[1];
  assign _EVAL_245 = _EVAL_32 != _EVAL_127;
  assign _EVAL_218 = ~_EVAL_88;
  assign _EVAL_45 = _EVAL_192 & _EVAL_61;
  assign _EVAL_249 = $signed(_EVAL_211) & -33'sh2000;
  assign _EVAL_151 = _EVAL_197 & _EVAL_231;
  assign _EVAL_70 = _EVAL_204 | _EVAL_7;
  assign _EVAL_43 = 2'h1 << _EVAL_0;
  assign _EVAL_271 = ~_EVAL;
  assign _EVAL_65 = _EVAL_199 | _EVAL_26;
  assign _EVAL_277 = _EVAL_180 | _EVAL_7;
  assign _EVAL_292 = _EVAL_15 == _EVAL_230;
  assign _EVAL_122 = _EVAL_300 == 4'h0;
  assign _EVAL_50 = ~_EVAL_37;
  assign _EVAL_243 = ~_EVAL_157;
  assign _EVAL_84 = ~_EVAL_254;
  assign _EVAL_119 = _EVAL_225 | _EVAL_99;
  assign _EVAL_174 = _EVAL_157 >> _EVAL_0;
  assign _EVAL_97 = $signed(_EVAL_153) & -33'shc000;
  assign _EVAL_222 = _EVAL_274 | _EVAL_7;
  assign _EVAL_152 = _EVAL_291 & _EVAL_37;
  assign _EVAL_276 = _EVAL_105;
  assign _EVAL_274 = _EVAL_271 == 4'h0;
  assign _EVAL_169 = _EVAL_34 | _EVAL_7;
  assign _EVAL_57 = _EVAL_38 | _EVAL_7;
  assign _EVAL_161 = ~_EVAL_166;
  assign _EVAL_294 = _EVAL_243 | _EVAL_111;
  assign _EVAL_172 = _EVAL_0 == _EVAL_278;
  assign _EVAL_220 = _EVAL_94 - 6'h1;
  assign _EVAL_179 = ~_EVAL_13;
  assign _EVAL_26 = $signed(_EVAL_198) == 33'sh0;
  assign _EVAL_198 = _EVAL_209;
  assign _EVAL_128 = _EVAL_200 | _EVAL_7;
  assign _EVAL_153 = {1'b0,$signed(_EVAL_311)};
  assign _EVAL_177 = _EVAL_268 | _EVAL_7;
  assign _EVAL_141 = _EVAL_203 | _EVAL_7;
  assign _EVAL_261 = ~_EVAL_7;
  assign _EVAL_289 = _EVAL_4 == 3'h0;
  assign _EVAL_61 = _EVAL_63 | _EVAL_301;
  assign _EVAL_284 = _EVAL_179 | _EVAL_7;
  assign _EVAL_291 = _EVAL_17[1];
  assign _EVAL_207 = ~_EVAL_188;
  assign _EVAL_253 = _EVAL_144 == 6'h0;
  assign _EVAL_19 = _EVAL_119 | _EVAL_112;
  assign _EVAL_20 = _EVAL_192 & _EVAL_63;
  assign _EVAL_138 = _EVAL_167[5:0];
  assign _EVAL_184 = ~_EVAL_57;
  assign _EVAL_312 = _EVAL_94 == 6'h0;
  assign _EVAL_318 = _EVAL_56 | _EVAL_146;
  assign _EVAL_164 = ~_EVAL_109;
  assign _EVAL_170 = _EVAL_192 & _EVAL_136;
  assign _EVAL_38 = _EVAL_11 == 2'h0;
  assign _EVAL_191 = _EVAL_255 | _EVAL_272;
  assign _EVAL_269 = _EVAL_10 == 3'h2;
  assign _EVAL_150 = _EVAL_115 | _EVAL_7;
  assign _EVAL_36 = _EVAL_119 | _EVAL_223;
  assign _EVAL_133 = _EVAL_305 | _EVAL_7;
  assign _EVAL_175 = _EVAL_1 & _EVAL_306;
  assign _EVAL_96 = _EVAL_14 & _EVAL_1;
  assign _EVAL_282 = _EVAL_160 | _EVAL_7;
  assign _EVAL_286 = ~_EVAL_277;
  assign _EVAL_69 = _EVAL_85;
  assign _EVAL_33 = _EVAL_10 == 3'h7;
  assign _EVAL_239 = _EVAL_12 & _EVAL_33;
  assign _EVAL_86 = ~_EVAL_32;
  assign _EVAL_80 = _EVAL_96 & _EVAL_210;
  assign _EVAL_137 = _EVAL_32 | _EVAL_157;
  assign _EVAL_79 = _EVAL_252 & _EVAL_307;
  assign _EVAL_113 = _EVAL_17 == _EVAL_185;
  assign _EVAL_264 = ~_EVAL_27;
  assign _EVAL_270 = _EVAL_12 & _EVAL_309;
  assign _EVAL_246 = _EVAL_12 & _EVAL_316;
  assign _EVAL_263 = _EVAL_294 | _EVAL_241;
  assign _EVAL_90 = _EVAL_151 ? 2'h1 : 2'h0;
  assign _EVAL_176 = _EVAL_87 | _EVAL_7;
  assign _EVAL_127 = _EVAL_90[0];
  assign _EVAL_224 = _EVAL_12 & _EVAL_269;
  assign _EVAL_71 = _EVAL_193 | _EVAL_7;
  assign _EVAL_211 = {1'b0,$signed(_EVAL_187)};
  assign _EVAL_108 = _EVAL_12 & _EVAL_267;
  assign _EVAL_203 = _EVAL_4 == _EVAL_303;
  assign _EVAL_190 = _EVAL_225 | _EVAL_7;
  assign _EVAL_35 = ~_EVAL_208;
  assign _EVAL_68 = _EVAL_6[0];
  assign _EVAL_217 = _EVAL_280[7:2];
  assign _EVAL_225 = _EVAL_6 >= 4'h2;
  assign _EVAL_49 = _EVAL_16 == 3'h0;
  assign _EVAL_272 = $signed(_EVAL_276) == 33'sh0;
  assign _EVAL_111 = plusarg_reader_out == 32'h0;
  assign _EVAL_46 = _EVAL_12 & _EVAL_248;
  assign _EVAL_192 = _EVAL_6 <= 4'h2;
  assign _EVAL_25 = _EVAL_135 | _EVAL_7;
  assign _EVAL_201 = {1'b0,$signed(_EVAL_279)};
  assign _EVAL_182 = _EVAL_1 & _EVAL_91;
  assign _EVAL_205 = ~_EVAL_317;
  assign _EVAL_140 = _EVAL_124 | 2'h1;
  assign _EVAL_215 = ~_EVAL_293;
  assign _EVAL_117 = _EVAL_1 & _EVAL_82;
  assign _EVAL_259 = _EVAL_10 == 3'h6;
  assign _EVAL_37 = _EVAL_17[0];
  assign _EVAL_124 = 2'h1 << _EVAL_68;
  assign _EVAL_29 = ~_EVAL_190;
  assign _EVAL_306 = _EVAL_4 == 3'h6;
  assign _EVAL_189 = _EVAL_16 <= 3'h3;
  assign _EVAL_228 = ~_EVAL_240;
  assign _EVAL_104 = {1'b0,$signed(_EVAL_17)};
  assign _EVAL_196 = _EVAL_97;
  assign _EVAL_279 = _EVAL_17 ^ 32'h20000000;
  assign _EVAL_219 = _EVAL_251 & _EVAL_126;
  assign _EVAL_313 = _EVAL_1 & _EVAL_106;
  assign _EVAL_307 = $signed(_EVAL_69) == 33'sh0;
  assign _EVAL_44 = _EVAL_6 <= 4'h6;
  assign _EVAL_202 = ~_EVAL_284;
  assign _EVAL_212 = ~_EVAL_291;
  assign _EVAL_216 = ~_EVAL_141;
  assign _EVAL_125 = ~_EVAL_282;
  assign _EVAL_132 = ~_EVAL_150;
  assign _EVAL_21 = ~_EVAL_214;
  assign _EVAL_256 = _EVAL_83[5:0];
  assign _EVAL_229 = _EVAL_140[0];
  assign _EVAL_116 = _EVAL_308 ? _EVAL_43 : 2'h0;
  assign _EVAL_297 = _EVAL_225 | _EVAL_302;
  assign _EVAL_260 = _EVAL_17 & _EVAL_165;
  assign _EVAL_309 = _EVAL_10 == 3'h0;
  assign _EVAL_168 = ~_EVAL_235;
  assign _EVAL_75 = _EVAL_296 | _EVAL_7;
  assign _EVAL_120 = _EVAL_159 | _EVAL_7;
  assign _EVAL_197 = _EVAL_96 & _EVAL_253;
  assign _EVAL_48 = _EVAL_76 & _EVAL_258;
  assign _EVAL_209 = $signed(_EVAL_104) & -33'sh5000;
  assign _EVAL_298 = ~_EVAL_174;
  assign _EVAL_227 = ~_EVAL_71;
  assign _EVAL_167 = _EVAL_144 - 6'h1;
  assign _EVAL_173 = ~_EVAL_107;
  assign _EVAL_66 = _EVAL_16 != 3'h0;
  assign _EVAL_183 = ~_EVAL_75;
  assign _EVAL_302 = _EVAL_281 & _EVAL_212;
  assign _EVAL_109 = _EVAL_139 | _EVAL_7;
  assign _EVAL_53 = _EVAL_122 | _EVAL_7;
  assign _EVAL_156 = ~_EVAL_176;
  assign _EVAL_254 = _EVAL_137 | _EVAL_7;
  assign _EVAL_99 = _EVAL_281 & _EVAL_291;
  assign _EVAL_146 = _EVAL_192 & _EVAL_301;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_22 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_64 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_77 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_78 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_94 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_144 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_154 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_157 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_181 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_185 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_186 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_226 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_230 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_278 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_303 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_304 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_3) begin
    if (_EVAL_219) begin
      _EVAL_22 <= _EVAL_10;
    end
    if (_EVAL_7) begin
      _EVAL_64 <= 6'h0;
    end else if (_EVAL_251) begin
      if (_EVAL_126) begin
        if (_EVAL_168) begin
          _EVAL_64 <= _EVAL_217;
        end else begin
          _EVAL_64 <= 6'h0;
        end
      end else begin
        _EVAL_64 <= _EVAL_256;
      end
    end
    if (_EVAL_80) begin
      _EVAL_77 <= _EVAL_2;
    end
    if (_EVAL_7) begin
      _EVAL_78 <= 32'h0;
    end else if (_EVAL_73) begin
      _EVAL_78 <= 32'h0;
    end else begin
      _EVAL_78 <= _EVAL_237;
    end
    if (_EVAL_7) begin
      _EVAL_94 <= 6'h0;
    end else if (_EVAL_251) begin
      if (_EVAL_312) begin
        if (_EVAL_168) begin
          _EVAL_94 <= _EVAL_217;
        end else begin
          _EVAL_94 <= 6'h0;
        end
      end else begin
        _EVAL_94 <= _EVAL_98;
      end
    end
    if (_EVAL_7) begin
      _EVAL_144 <= 6'h0;
    end else if (_EVAL_96) begin
      if (_EVAL_253) begin
        if (_EVAL_315) begin
          _EVAL_144 <= _EVAL_52;
        end else begin
          _EVAL_144 <= 6'h0;
        end
      end else begin
        _EVAL_144 <= _EVAL_138;
      end
    end
    if (_EVAL_219) begin
      _EVAL_154 <= _EVAL_16;
    end
    if (_EVAL_7) begin
      _EVAL_157 <= 1'h0;
    end else begin
      _EVAL_157 <= _EVAL_48;
    end
    if (_EVAL_80) begin
      _EVAL_181 <= _EVAL_11;
    end
    if (_EVAL_219) begin
      _EVAL_185 <= _EVAL_17;
    end
    if (_EVAL_80) begin
      _EVAL_186 <= _EVAL_5;
    end
    if (_EVAL_7) begin
      _EVAL_226 <= 6'h0;
    end else if (_EVAL_96) begin
      if (_EVAL_210) begin
        if (_EVAL_315) begin
          _EVAL_226 <= _EVAL_52;
        end else begin
          _EVAL_226 <= 6'h0;
        end
      end else begin
        _EVAL_226 <= _EVAL_232;
      end
    end
    if (_EVAL_80) begin
      _EVAL_230 <= _EVAL_15;
    end
    if (_EVAL_219) begin
      _EVAL_278 <= _EVAL_0;
    end
    if (_EVAL_80) begin
      _EVAL_303 <= _EVAL_4;
    end
    if (_EVAL_219) begin
      _EVAL_304 <= _EVAL_6;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(deefc4fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c045b10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d41d7a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(788be241)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_31) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3aadc74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2c26e6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27cd3594)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f7a370b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_275) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ded6317e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_31) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70184fc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3148404)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68d5993a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91563fcb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(456e29ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4588881d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a1aefcb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35e4796a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(998d1c37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e02605c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc08c451)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(923d4d5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c54f1588)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89020e9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66d3bf75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_288) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ddb4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24ff4942)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26403382)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0c26c86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(525354d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d03f4f9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6f99c14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_264) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_288) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27ebf185)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b06458e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_31) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e43d3f5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b32545a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86778e23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6d4cefe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5091346)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(148f949)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f38558b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57cbab58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8f0cce8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d51e7448)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f37d9d0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66cb9a43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_287) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(158c208c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29f94eb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a898ab5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0920e6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ea44e47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15d90829)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63dbc405)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(492a9121)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(615849fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f69f7af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de510041)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c15f1b2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64d413c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fd6b8a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ca0e850)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3704f0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_275) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96f45313)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1feef216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_31) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b7f685)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(622d40ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(750350)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5b3c06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26e86f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e217562d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_287) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61fb980d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_264) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35edce6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(baf0bfe4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(939dbe0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13897c50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(741e8778)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(536044aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa578dd3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f89e45ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(517ee29d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e54ec1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71f28c1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0415e9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(568561de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70fbb9d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
