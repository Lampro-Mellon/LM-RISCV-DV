//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_156(
  input         _EVAL,
  output        _EVAL_0,
  input  [31:0] _EVAL_1,
  input  [1:0]  _EVAL_2,
  input         _EVAL_3,
  output        _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [29:0] _EVAL_10,
  input  [1:0]  _EVAL_11,
  input  [31:0] _EVAL_12,
  input         _EVAL_13,
  input  [29:0] _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [29:0] _EVAL_17,
  input         _EVAL_18,
  input  [31:0] _EVAL_19,
  input  [1:0]  _EVAL_20,
  input         _EVAL_21,
  input         _EVAL_22,
  input  [1:0]  _EVAL_23,
  output        _EVAL_24,
  input  [29:0] _EVAL_25,
  input  [31:0] _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  input  [1:0]  _EVAL_30,
  input         _EVAL_31,
  input  [31:0] _EVAL_32,
  input         _EVAL_33
);
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire [31:0] _EVAL_37;
  wire  _EVAL_39;
  wire  _EVAL_41;
  wire [31:0] _EVAL_43;
  wire  _EVAL_44;
  wire [31:0] _EVAL_49;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire [31:0] _EVAL_63;
  wire [31:0] _EVAL_66;
  wire [31:0] _EVAL_67;
  wire [31:0] _EVAL_69;
  wire  _EVAL_72;
  wire [31:0] _EVAL_75;
  wire [31:0] _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire [31:0] _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_83;
  wire [31:0] _EVAL_84;
  wire [31:0] _EVAL_85;
  wire  _EVAL_88;
  wire [31:0] _EVAL_89;
  wire [31:0] _EVAL_91;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_101;
  wire [31:0] _EVAL_102;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_113;
  wire [31:0] _EVAL_116;
  wire  _EVAL_118;
  wire  _EVAL_120;
  wire [31:0] _EVAL_121;
  wire  _EVAL_123;
  wire  _EVAL_125;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire [31:0] _EVAL_139;
  wire [31:0] _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire [31:0] _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_150;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire [31:0] _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_167;
  wire  _EVAL_169;
  wire [31:0] _EVAL_170;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire [31:0] _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_178;
  wire [31:0] _EVAL_179;
  wire [31:0] _EVAL_181;
  wire [31:0] _EVAL_182;
  wire [31:0] _EVAL_184;
  wire  _EVAL_187;
  wire  _EVAL_193;
  wire  _EVAL_195;
  wire [31:0] _EVAL_196;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  assign _EVAL_184 = _EVAL_179 | 32'h3;
  assign _EVAL_178 = ~_EVAL_8;
  assign _EVAL_160 = _EVAL_13 | _EVAL_54;
  assign _EVAL_84 = _EVAL_32 ^ _EVAL_76;
  assign _EVAL_157 = _EVAL_7 | _EVAL_94;
  assign _EVAL_91 = _EVAL_147 | 32'h3;
  assign _EVAL_69 = ~_EVAL_175;
  assign _EVAL_97 = _EVAL_11[1];
  assign _EVAL_202 = _EVAL_167 ? _EVAL_105 : _EVAL_145;
  assign _EVAL_174 = _EVAL_49 == 32'h0;
  assign _EVAL_139 = {_EVAL_17, 2'h0};
  assign _EVAL_193 = ~_EVAL_3;
  assign _EVAL_55 = ~_EVAL_22;
  assign _EVAL_61 = ~_EVAL_148;
  assign _EVAL_113 = _EVAL_2[0];
  assign _EVAL_181 = _EVAL_32 ^ _EVAL_121;
  assign _EVAL_137 = _EVAL_58 & _EVAL_148;
  assign _EVAL_72 = ~_EVAL_33;
  assign _EVAL_62 = _EVAL_32 < _EVAL_85;
  assign _EVAL_143 = _EVAL_44 ? _EVAL_160 : _EVAL_146;
  assign _EVAL_81 = _EVAL_32 < _EVAL_76;
  assign _EVAL_44 = _EVAL_101 ? _EVAL_174 : _EVAL_150;
  assign _EVAL_76 = ~_EVAL_91;
  assign _EVAL_116 = ~_EVAL_139;
  assign _EVAL_43 = {_EVAL_10, 2'h0};
  assign _EVAL_125 = _EVAL_20[0];
  assign _EVAL_96 = _EVAL_167 ? _EVAL_157 : _EVAL_41;
  assign _EVAL_176 = _EVAL_120 & _EVAL_161;
  assign _EVAL_159 = _EVAL_181 & _EVAL_140;
  assign _EVAL_106 = _EVAL_30[1];
  assign _EVAL_39 = _EVAL_15 | _EVAL_54;
  assign _EVAL_0 = _EVAL_57 ? _EVAL_93 : _EVAL_202;
  assign _EVAL_120 = ~_EVAL_62;
  assign _EVAL_131 = _EVAL_34 & _EVAL_176;
  assign _EVAL_167 = _EVAL_106 ? _EVAL_123 : _EVAL_131;
  assign _EVAL_66 = _EVAL_32 ^ _EVAL_69;
  assign _EVAL_102 = ~_EVAL_12;
  assign _EVAL_141 = _EVAL_16 | _EVAL_94;
  assign _EVAL_123 = _EVAL_159 == 32'h0;
  assign _EVAL_67 = ~_EVAL_26;
  assign _EVAL_37 = _EVAL_32 ^ _EVAL_85;
  assign _EVAL_85 = ~_EVAL_75;
  assign _EVAL_130 = _EVAL_78 ? _EVAL_142 : _EVAL_198;
  assign _EVAL_150 = _EVAL_113 & _EVAL_156;
  assign _EVAL_80 = {_EVAL_25, 2'h0};
  assign _EVAL_118 = _EVAL_146 & _EVAL_193;
  assign _EVAL_142 = _EVAL_27 | _EVAL_169;
  assign _EVAL_196 = {_EVAL_14, 2'h0};
  assign _EVAL_94 = _EVAL_146 & _EVAL_72;
  assign _EVAL_195 = _EVAL_11[0];
  assign _EVAL_199 = _EVAL_195 & _EVAL_62;
  assign _EVAL_49 = _EVAL_84 & _EVAL_170;
  assign _EVAL_187 = _EVAL_44 ? _EVAL_39 : _EVAL_146;
  assign _EVAL_98 = _EVAL_5 | _EVAL_54;
  assign _EVAL_140 = ~_EVAL_19;
  assign _EVAL_170 = ~_EVAL_1;
  assign _EVAL_101 = _EVAL_2[1];
  assign _EVAL_77 = _EVAL_20[1];
  assign _EVAL_148 = _EVAL_32 < _EVAL_69;
  assign _EVAL_54 = _EVAL_146 & _EVAL_55;
  assign _EVAL_83 = _EVAL_29 | _EVAL_169;
  assign _EVAL_105 = _EVAL_31 | _EVAL_94;
  assign _EVAL_75 = _EVAL_116 | 32'h3;
  assign _EVAL_179 = ~_EVAL_196;
  assign _EVAL_175 = _EVAL_182 | 32'h3;
  assign _EVAL_121 = ~_EVAL_184;
  assign _EVAL_24 = _EVAL_57 ? _EVAL_132 : _EVAL_96;
  assign _EVAL_182 = ~_EVAL_43;
  assign _EVAL_34 = _EVAL_30[0];
  assign _EVAL_89 = _EVAL_37 & _EVAL_67;
  assign _EVAL_4 = _EVAL_57 ? _EVAL_88 : _EVAL_138;
  assign _EVAL_200 = _EVAL_21 | _EVAL_169;
  assign _EVAL_57 = _EVAL_97 ? _EVAL_35 : _EVAL_199;
  assign _EVAL_173 = _EVAL_125 & _EVAL_137;
  assign _EVAL_63 = _EVAL_66 & _EVAL_102;
  assign _EVAL_145 = _EVAL_78 ? _EVAL_200 : _EVAL_187;
  assign _EVAL_58 = ~_EVAL_161;
  assign _EVAL_93 = _EVAL_18 | _EVAL_118;
  assign _EVAL_198 = _EVAL_44 ? _EVAL_98 : _EVAL_146;
  assign _EVAL_78 = _EVAL_77 ? _EVAL_201 : _EVAL_173;
  assign _EVAL_146 = _EVAL_23 > 2'h1;
  assign _EVAL_88 = _EVAL_9 | _EVAL_118;
  assign _EVAL_169 = _EVAL_146 & _EVAL_178;
  assign _EVAL_201 = _EVAL_63 == 32'h0;
  assign _EVAL_161 = _EVAL_32 < _EVAL_121;
  assign _EVAL_138 = _EVAL_167 ? _EVAL_141 : _EVAL_130;
  assign _EVAL_147 = ~_EVAL_80;
  assign _EVAL_41 = _EVAL_78 ? _EVAL_83 : _EVAL_143;
  assign _EVAL_132 = _EVAL_6 | _EVAL_118;
  assign _EVAL_35 = _EVAL_89 == 32'h0;
  assign _EVAL_156 = _EVAL_61 & _EVAL_81;
endmodule
