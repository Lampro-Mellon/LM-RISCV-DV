//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_7_assert(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [31:0] _EVAL_7,
  input  [2:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [3:0]  _EVAL_13,
  input  [3:0]  _EVAL_14,
  input  [3:0]  _EVAL_15,
  input  [1:0]  _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18
);
  wire  _EVAL_19;
  reg [5:0] _EVAL_20;
  reg [31:0] _RAND_0;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire [1:0] _EVAL_29;
  wire  _EVAL_30;
  wire [22:0] _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  reg  _EVAL_34;
  reg [31:0] _RAND_1;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire [7:0] _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire [31:0] _EVAL_41;
  wire  _EVAL_42;
  wire [32:0] _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire [31:0] _EVAL_46;
  wire [5:0] _EVAL_47;
  wire  _EVAL_48;
  wire [5:0] _EVAL_49;
  wire  _EVAL_50;
  reg [2:0] _EVAL_51;
  reg [31:0] _RAND_2;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire [32:0] _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire [31:0] _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_72;
  reg [1:0] _EVAL_73;
  reg [31:0] _RAND_3;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire [1:0] _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire [1:0] _EVAL_79;
  wire [31:0] _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire [32:0] _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire [31:0] _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  reg [31:0] _EVAL_97;
  reg [31:0] _RAND_4;
  reg [5:0] _EVAL_98;
  reg [31:0] _RAND_5;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire [31:0] _EVAL_102;
  wire [6:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire [32:0] _EVAL_110;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  reg [5:0] _EVAL_117;
  reg [31:0] _RAND_6;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  reg [31:0] _EVAL_124;
  reg [31:0] _RAND_7;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire [32:0] _EVAL_128;
  wire  _EVAL_129;
  reg [5:0] _EVAL_130;
  reg [31:0] _RAND_8;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  reg [3:0] _EVAL_135;
  reg [31:0] _RAND_9;
  wire [3:0] _EVAL_136;
  wire [32:0] _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire [5:0] _EVAL_145;
  wire  _EVAL_146;
  wire [31:0] _EVAL_148;
  reg  _EVAL_149;
  reg [31:0] _RAND_10;
  wire [3:0] _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  reg [2:0] _EVAL_155;
  reg [31:0] _RAND_11;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire [1:0] _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  reg [1:0] _EVAL_165;
  reg [31:0] _RAND_12;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire [6:0] _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire [32:0] _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire [1:0] _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire [32:0] _EVAL_182;
  wire [7:0] _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire [32:0] _EVAL_189;
  wire [22:0] _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire [32:0] _EVAL_200;
  reg [3:0] _EVAL_201;
  reg [31:0] _RAND_13;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire [1:0] _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire [5:0] _EVAL_211;
  wire  _EVAL_212;
  wire [1:0] _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire [32:0] _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire [1:0] _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire [6:0] _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire [1:0] _EVAL_232;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire [1:0] _EVAL_248;
  wire [1:0] _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire [3:0] _EVAL_263;
  wire [32:0] _EVAL_264;
  wire  _EVAL_265;
  wire [32:0] _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  reg  _EVAL_276;
  reg [31:0] _RAND_14;
  wire  _EVAL_277;
  wire [32:0] _EVAL_278;
  wire  _EVAL_279;
  wire [3:0] _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire [5:0] _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  reg [2:0] _EVAL_290;
  reg [31:0] _RAND_15;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire [32:0] _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire [31:0] _EVAL_297;
  wire  _EVAL_298;
  wire [32:0] _EVAL_299;
  reg  _EVAL_300;
  reg [31:0] _RAND_16;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire [32:0] _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire [1:0] _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire [7:0] _EVAL_311;
  wire [5:0] _EVAL_312;
  wire [7:0] _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire [32:0] _EVAL_316;
  wire  _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire [6:0] _EVAL_321;
  wire [32:0] _EVAL_322;
  wire  _EVAL_323;
  wire  _EVAL_324;
  wire  _EVAL_325;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_153 = _EVAL_121 | _EVAL_11;
  assign _EVAL_214 = ~_EVAL_294;
  assign _EVAL_102 = _EVAL_7 ^ 32'h3000;
  assign _EVAL_196 = _EVAL_152 | _EVAL_185;
  assign _EVAL_231 = ~_EVAL_38;
  assign _EVAL_158 = ~_EVAL_216;
  assign _EVAL_143 = ~_EVAL_28;
  assign _EVAL_110 = _EVAL_322;
  assign _EVAL_67 = _EVAL_125 | _EVAL_27;
  assign _EVAL_240 = _EVAL_146 & _EVAL_27;
  assign _EVAL_221 = _EVAL_142 | _EVAL_11;
  assign _EVAL_310 = _EVAL_13 <= 4'h6;
  assign _EVAL_264 = _EVAL_124 + 32'h1;
  assign _EVAL_243 = _EVAL_9[0];
  assign _EVAL_107 = _EVAL_324 | _EVAL_11;
  assign _EVAL_170 = _EVAL_6 & _EVAL_238;
  assign _EVAL_162 = _EVAL_79 | _EVAL_165;
  assign _EVAL_281 = _EVAL_295 | _EVAL_178;
  assign _EVAL_185 = _EVAL_310 & _EVAL_66;
  assign _EVAL_305 = _EVAL_130 == 6'h0;
  assign _EVAL_322 = $signed(_EVAL_176) & -33'sh5000;
  assign _EVAL_95 = _EVAL_14 == _EVAL_201;
  assign _EVAL_286 = $signed(_EVAL_110) == 33'sh0;
  assign _EVAL_48 = _EVAL_9 == 3'h4;
  assign _EVAL_128 = $signed(_EVAL_293) & -33'sh2000;
  assign _EVAL_74 = ~_EVAL_30;
  assign _EVAL_154 = ~_EVAL_221;
  assign _EVAL_267 = _EVAL_281 | _EVAL_195;
  assign _EVAL_172 = _EVAL_98 - 6'h1;
  assign _EVAL_244 = _EVAL_255 | _EVAL_11;
  assign _EVAL_261 = _EVAL_35 & _EVAL_62;
  assign _EVAL_284 = _EVAL_9 == 3'h2;
  assign _EVAL_257 = _EVAL_5 == _EVAL_34;
  assign _EVAL_22 = _EVAL_185 | _EVAL_151;
  assign _EVAL_87 = ~_EVAL_288;
  assign _EVAL_180 = _EVAL_6 & _EVAL_75;
  assign _EVAL_72 = _EVAL_146 & _EVAL_125;
  assign _EVAL_236 = _EVAL_7[0];
  assign _EVAL_303 = _EVAL_43;
  assign _EVAL_45 = _EVAL_9 == 3'h1;
  assign _EVAL_256 = ~_EVAL_10;
  assign _EVAL_24 = _EVAL_257 | _EVAL_11;
  assign _EVAL_58 = {1'b0,$signed(_EVAL_80)};
  assign _EVAL_298 = ~_EVAL_244;
  assign _EVAL_89 = ~_EVAL_138;
  assign _EVAL_166 = _EVAL_212 | _EVAL_11;
  assign _EVAL_191 = _EVAL_230 | _EVAL_259;
  assign _EVAL_200 = _EVAL_299;
  assign _EVAL_186 = ~_EVAL_246;
  assign _EVAL_26 = _EVAL <= 3'h4;
  assign _EVAL_99 = ~_EVAL_197;
  assign _EVAL_146 = _EVAL_13 <= 4'h2;
  assign _EVAL_192 = ~_EVAL_131;
  assign _EVAL_138 = _EVAL_69 | _EVAL_11;
  assign _EVAL_250 = ~_EVAL_260;
  assign _EVAL_189 = $signed(_EVAL_83) & -33'sh1000000;
  assign _EVAL_36 = _EVAL_256 | _EVAL_11;
  assign _EVAL_122 = _EVAL != 3'h0;
  assign _EVAL_142 = _EVAL == 3'h0;
  assign _EVAL_277 = _EVAL_18 & _EVAL_284;
  assign _EVAL_275 = ~_EVAL_234;
  assign _EVAL_223 = ~_EVAL_107;
  assign _EVAL_148 = _EVAL_7 & _EVAL_297;
  assign _EVAL_88 = _EVAL_117 == 6'h0;
  assign _EVAL_220 = _EVAL_189;
  assign _EVAL_91 = _EVAL_271 | _EVAL_11;
  assign _EVAL_179 = ~_EVAL_248;
  assign _EVAL_248 = _EVAL_261 ? _EVAL_213 : 2'h0;
  assign _EVAL_176 = {1'b0,$signed(_EVAL_7)};
  assign _EVAL_255 = _EVAL_64 | _EVAL_3;
  assign _EVAL_271 = _EVAL_8 == _EVAL_290;
  assign _EVAL_260 = _EVAL_292 | _EVAL_11;
  assign _EVAL_84 = _EVAL_20 == 6'h0;
  assign _EVAL_232 = 2'h1 << _EVAL_1;
  assign _EVAL_212 = _EVAL_148 == 32'h0;
  assign _EVAL_174 = _EVAL_124 < plusarg_reader_out;
  assign _EVAL_254 = _EVAL_249[0];
  assign _EVAL_104 = _EVAL_309 | _EVAL_11;
  assign _EVAL_70 = _EVAL_150 == 4'h0;
  assign _EVAL_205 = _EVAL_16 <= 2'h2;
  assign _EVAL_125 = _EVAL_198 | _EVAL_286;
  assign _EVAL_263 = {_EVAL_100,_EVAL_199,_EVAL_267,_EVAL_141};
  assign _EVAL_266 = $signed(_EVAL_278) & -33'sh2000;
  assign _EVAL_141 = _EVAL_281 | _EVAL_160;
  assign _EVAL_121 = _EVAL_17 == _EVAL_300;
  assign _EVAL_44 = _EVAL_159 | _EVAL_11;
  assign _EVAL_105 = _EVAL_52 | _EVAL_11;
  assign _EVAL_159 = _EVAL_13 == _EVAL_135;
  assign _EVAL_112 = _EVAL_9 <= 3'h6;
  assign _EVAL_80 = _EVAL_7 ^ 32'h80000000;
  assign _EVAL_151 = _EVAL_56 & _EVAL_94;
  assign _EVAL_178 = _EVAL_253 & _EVAL_262;
  assign _EVAL_47 = _EVAL_228[5:0];
  assign _EVAL_59 = ~_EVAL_305;
  assign _EVAL_239 = _EVAL_6 & _EVAL_318;
  assign _EVAL_173 = _EVAL_94 | _EVAL_320;
  assign _EVAL_289 = _EVAL_22 | _EVAL_240;
  assign _EVAL_315 = _EVAL_280 == 4'h0;
  assign _EVAL_150 = ~_EVAL_15;
  assign _EVAL_37 = ~_EVAL_183;
  assign _EVAL_258 = _EVAL_193 | _EVAL_11;
  assign _EVAL_288 = _EVAL_26 | _EVAL_11;
  assign _EVAL_76 = _EVAL_165 | _EVAL_79;
  assign _EVAL_273 = _EVAL_6 & _EVAL_219;
  assign _EVAL_237 = _EVAL_163 & _EVAL_317;
  assign _EVAL_216 = _EVAL_181 | _EVAL_11;
  assign _EVAL_195 = _EVAL_254 & _EVAL_118;
  assign _EVAL_242 = ~_EVAL_91;
  assign _EVAL_123 = ~_EVAL_302;
  assign _EVAL_115 = ~_EVAL_106;
  assign _EVAL_137 = _EVAL_266;
  assign _EVAL_321 = _EVAL_130 - 6'h1;
  assign _EVAL_21 = _EVAL_253 & _EVAL_163;
  assign _EVAL_323 = _EVAL <= 3'h1;
  assign _EVAL_218 = _EVAL_9 == 3'h6;
  assign _EVAL_230 = _EVAL_0 & _EVAL_6;
  assign _EVAL_82 = ~_EVAL_11;
  assign _EVAL_168 = ~_EVAL_229;
  assign _EVAL_126 = _EVAL_16 == _EVAL_73;
  assign _EVAL_318 = _EVAL_8 == 3'h7;
  assign _EVAL_229 = _EVAL_245 | _EVAL_11;
  assign _EVAL_103 = _EVAL_20 - 6'h1;
  assign _EVAL_210 = _EVAL == _EVAL_155;
  assign _EVAL_27 = $signed(_EVAL_316) == 33'sh0;
  assign _EVAL_131 = _EVAL_101 | _EVAL_11;
  assign _EVAL_193 = _EVAL_14 >= 4'h2;
  assign _EVAL_197 = _EVAL_139 | _EVAL_11;
  assign _EVAL_68 = _EVAL_295 | _EVAL_11;
  assign _EVAL_118 = _EVAL_262 & _EVAL_236;
  assign _EVAL_213 = 2'h1 << _EVAL_5;
  assign _EVAL_75 = _EVAL_8 == 3'h6;
  assign _EVAL_246 = _EVAL_165 != 2'h0;
  assign _EVAL_219 = _EVAL_8 == 3'h1;
  assign _EVAL_144 = ~_EVAL_53;
  assign _EVAL_32 = _EVAL_8 == 3'h3;
  assign _EVAL_49 = _EVAL_172[5:0];
  assign _EVAL_160 = _EVAL_254 & _EVAL_50;
  assign _EVAL_40 = _EVAL_72 | _EVAL_151;
  assign _EVAL_90 = ~_EVAL_287;
  assign _EVAL_316 = _EVAL_128;
  assign _EVAL_228 = _EVAL_117 - 6'h1;
  assign _EVAL_169 = _EVAL_188 | _EVAL_11;
  assign _EVAL_235 = _EVAL_259 & _EVAL_305;
  assign _EVAL_269 = _EVAL_9 == 3'h0;
  assign _EVAL_301 = ~_EVAL_215;
  assign _EVAL_33 = ~_EVAL_166;
  assign _EVAL_252 = _EVAL_8 == 3'h2;
  assign _EVAL_253 = _EVAL_249[1];
  assign _EVAL_293 = {1'b0,$signed(_EVAL_92)};
  assign _EVAL_127 = _EVAL_13[0];
  assign _EVAL_100 = _EVAL_132 | _EVAL_247;
  assign _EVAL_62 = ~_EVAL_218;
  assign _EVAL_167 = ~_EVAL_77;
  assign _EVAL_94 = $signed(_EVAL_303) == 33'sh0;
  assign _EVAL_19 = _EVAL_225[0];
  assign _EVAL_208 = _EVAL_165 >> _EVAL_1;
  assign _EVAL_114 = _EVAL_18 & _EVAL_269;
  assign _EVAL_136 = ~_EVAL_263;
  assign _EVAL_206 = _EVAL_6 & _EVAL_140;
  assign _EVAL_177 = _EVAL_291 | _EVAL_11;
  assign _EVAL_225 = _EVAL_162 >> _EVAL_5;
  assign _EVAL_53 = _EVAL_323 | _EVAL_11;
  assign _EVAL_57 = _EVAL_60 | _EVAL_174;
  assign _EVAL_106 = _EVAL_40 | _EVAL_11;
  assign _EVAL_54 = ~_EVAL_258;
  assign _EVAL_291 = _EVAL_1 == _EVAL_276;
  assign _EVAL_182 = {1'b0,$signed(_EVAL_102)};
  assign _EVAL_324 = _EVAL_7 == _EVAL_97;
  assign _EVAL_198 = _EVAL_81 | _EVAL_320;
  assign _EVAL_238 = _EVAL_8 == 3'h5;
  assign _EVAL_65 = ~_EVAL_304;
  assign _EVAL_312 = _EVAL_103[5:0];
  assign _EVAL_320 = $signed(_EVAL_220) == 33'sh0;
  assign _EVAL_204 = _EVAL_18 & _EVAL_45;
  assign _EVAL_56 = _EVAL_13 <= 4'h8;
  assign _EVAL_224 = _EVAL_6 & _EVAL_217;
  assign _EVAL_79 = _EVAL_314 ? _EVAL_232 : 2'h0;
  assign _EVAL_183 = _EVAL_31[7:0];
  assign _EVAL_63 = _EVAL_7 ^ 32'h40000000;
  assign _EVAL_209 = ~_EVAL_296;
  assign _EVAL_28 = _EVAL_93 | _EVAL_11;
  assign _EVAL_278 = {1'b0,$signed(_EVAL_63)};
  assign _EVAL_140 = _EVAL_8 == 3'h4;
  assign _EVAL_302 = _EVAL_126 | _EVAL_11;
  assign _EVAL_297 = {{24'd0}, _EVAL_37};
  assign _EVAL_60 = _EVAL_186 | _EVAL_161;
  assign _EVAL_279 = ~_EVAL_169;
  assign _EVAL_157 = _EVAL_163 & _EVAL_236;
  assign _EVAL_227 = ~_EVAL_177;
  assign _EVAL_306 = ~_EVAL_119;
  assign _EVAL_314 = _EVAL_230 & _EVAL_84;
  assign _EVAL_133 = _EVAL_8[2];
  assign _EVAL_311 = ~_EVAL_313;
  assign _EVAL_163 = _EVAL_7[1];
  assign _EVAL_64 = ~_EVAL_2;
  assign _EVAL_211 = _EVAL_37[7:2];
  assign _EVAL_93 = ~_EVAL_3;
  assign _EVAL_134 = _EVAL_18 & _EVAL_129;
  assign _EVAL_69 = _EVAL_16 != 2'h2;
  assign _EVAL_283 = _EVAL_311[7:2];
  assign _EVAL_120 = ~_EVAL_308;
  assign _EVAL_202 = _EVAL_18 & _EVAL_48;
  assign _EVAL_265 = ~_EVAL_153;
  assign _EVAL_304 = _EVAL_315 | _EVAL_11;
  assign _EVAL_308 = _EVAL_70 | _EVAL_11;
  assign _EVAL_31 = 23'hff << _EVAL_13;
  assign _EVAL_319 = _EVAL_79 != _EVAL_248;
  assign _EVAL_164 = ~_EVAL_133;
  assign _EVAL_190 = 23'hff << _EVAL_14;
  assign _EVAL_295 = _EVAL_13 >= 4'h2;
  assign _EVAL_282 = _EVAL_208[0];
  assign _EVAL_249 = _EVAL_29 | 2'h1;
  assign _EVAL_299 = $signed(_EVAL_58) & -33'shc000;
  assign _EVAL_25 = ~_EVAL_268;
  assign _EVAL_29 = 2'h1 << _EVAL_127;
  assign _EVAL_181 = _EVAL_9 == _EVAL_51;
  assign _EVAL_42 = ~_EVAL_68;
  assign _EVAL_92 = _EVAL_7 ^ 32'h20000000;
  assign _EVAL_317 = ~_EVAL_236;
  assign _EVAL_85 = _EVAL_173 | _EVAL_286;
  assign _EVAL_292 = _EVAL_146 & _EVAL_270;
  assign _EVAL_139 = _EVAL_16 == 2'h0;
  assign _EVAL_41 = _EVAL_264[31:0];
  assign _EVAL_35 = _EVAL_259 & _EVAL_88;
  assign _EVAL_285 = ~_EVAL_171;
  assign _EVAL_187 = ~_EVAL_104;
  assign _EVAL_188 = _EVAL_319 | _EVAL_275;
  assign _EVAL_52 = _EVAL <= 3'h2;
  assign _EVAL_77 = _EVAL_210 | _EVAL_11;
  assign _EVAL_108 = ~_EVAL_44;
  assign _EVAL_203 = _EVAL_15 == _EVAL_263;
  assign _EVAL_215 = _EVAL_98 == 6'h0;
  assign _EVAL_294 = _EVAL_122 | _EVAL_11;
  assign _EVAL_50 = _EVAL_262 & _EVAL_317;
  assign _EVAL_247 = _EVAL_254 & _EVAL_157;
  assign _EVAL_30 = _EVAL_64 | _EVAL_11;
  assign _EVAL_113 = _EVAL_57 | _EVAL_11;
  assign _EVAL_96 = ~_EVAL_105;
  assign _EVAL_296 = _EVAL_19 | _EVAL_11;
  assign _EVAL_226 = _EVAL_6 & _EVAL_301;
  assign _EVAL_78 = ~_EVAL_113;
  assign _EVAL_270 = _EVAL_85 | _EVAL_27;
  assign _EVAL_287 = _EVAL_112 | _EVAL_11;
  assign _EVAL_161 = plusarg_reader_out == 32'h0;
  assign _EVAL_119 = _EVAL_203 | _EVAL_11;
  assign _EVAL_81 = $signed(_EVAL_200) == 33'sh0;
  assign _EVAL_145 = _EVAL_321[5:0];
  assign _EVAL_325 = _EVAL_18 & _EVAL_218;
  assign _EVAL_245 = _EVAL <= 3'h3;
  assign _EVAL_101 = _EVAL_196 | _EVAL_151;
  assign _EVAL_313 = _EVAL_190[7:0];
  assign _EVAL_234 = _EVAL_79 != 2'h0;
  assign _EVAL_66 = $signed(_EVAL_137) == 33'sh0;
  assign _EVAL_280 = _EVAL_15 & _EVAL_136;
  assign _EVAL_23 = _EVAL_6 & _EVAL_32;
  assign _EVAL_129 = _EVAL_9 == 3'h5;
  assign _EVAL_38 = _EVAL_205 | _EVAL_11;
  assign _EVAL_217 = _EVAL_8 == 3'h0;
  assign _EVAL_259 = _EVAL_12 & _EVAL_18;
  assign _EVAL_241 = ~_EVAL_274;
  assign _EVAL_268 = _EVAL_95 | _EVAL_11;
  assign _EVAL_175 = _EVAL_230 & _EVAL_215;
  assign _EVAL_171 = _EVAL_222 | _EVAL_11;
  assign _EVAL_199 = _EVAL_132 | _EVAL_61;
  assign _EVAL_184 = ~_EVAL_24;
  assign _EVAL_43 = $signed(_EVAL_182) & -33'sh1000;
  assign _EVAL_61 = _EVAL_254 & _EVAL_237;
  assign _EVAL_86 = _EVAL_18 & _EVAL_59;
  assign _EVAL_83 = {1'b0,$signed(_EVAL_46)};
  assign _EVAL_309 = ~_EVAL_282;
  assign _EVAL_46 = _EVAL_7 ^ 32'h2000000;
  assign _EVAL_307 = _EVAL_76 & _EVAL_179;
  assign _EVAL_262 = ~_EVAL_163;
  assign _EVAL_55 = ~_EVAL_36;
  assign _EVAL_132 = _EVAL_295 | _EVAL_21;
  assign _EVAL_152 = _EVAL_146 & _EVAL_67;
  assign _EVAL_274 = _EVAL_289 | _EVAL_11;
  assign _EVAL_39 = _EVAL_6 & _EVAL_252;
  assign _EVAL_222 = _EVAL_2 == _EVAL_149;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_20 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_34 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_51 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_73 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_97 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_98 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_117 = _RAND_6[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_124 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_130 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_135 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_149 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_155 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_165 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_201 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_276 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_290 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_300 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_4) begin
    if (_EVAL_11) begin
      _EVAL_20 <= 6'h0;
    end else if (_EVAL_230) begin
      if (_EVAL_84) begin
        if (_EVAL_164) begin
          _EVAL_20 <= _EVAL_211;
        end else begin
          _EVAL_20 <= 6'h0;
        end
      end else begin
        _EVAL_20 <= _EVAL_312;
      end
    end
    if (_EVAL_235) begin
      _EVAL_34 <= _EVAL_5;
    end
    if (_EVAL_235) begin
      _EVAL_51 <= _EVAL_9;
    end
    if (_EVAL_235) begin
      _EVAL_73 <= _EVAL_16;
    end
    if (_EVAL_175) begin
      _EVAL_97 <= _EVAL_7;
    end
    if (_EVAL_11) begin
      _EVAL_98 <= 6'h0;
    end else if (_EVAL_230) begin
      if (_EVAL_215) begin
        if (_EVAL_164) begin
          _EVAL_98 <= _EVAL_211;
        end else begin
          _EVAL_98 <= 6'h0;
        end
      end else begin
        _EVAL_98 <= _EVAL_49;
      end
    end
    if (_EVAL_11) begin
      _EVAL_117 <= 6'h0;
    end else if (_EVAL_259) begin
      if (_EVAL_88) begin
        if (_EVAL_243) begin
          _EVAL_117 <= _EVAL_283;
        end else begin
          _EVAL_117 <= 6'h0;
        end
      end else begin
        _EVAL_117 <= _EVAL_47;
      end
    end
    if (_EVAL_11) begin
      _EVAL_124 <= 32'h0;
    end else if (_EVAL_191) begin
      _EVAL_124 <= 32'h0;
    end else begin
      _EVAL_124 <= _EVAL_41;
    end
    if (_EVAL_11) begin
      _EVAL_130 <= 6'h0;
    end else if (_EVAL_259) begin
      if (_EVAL_305) begin
        if (_EVAL_243) begin
          _EVAL_130 <= _EVAL_283;
        end else begin
          _EVAL_130 <= 6'h0;
        end
      end else begin
        _EVAL_130 <= _EVAL_145;
      end
    end
    if (_EVAL_175) begin
      _EVAL_135 <= _EVAL_13;
    end
    if (_EVAL_235) begin
      _EVAL_149 <= _EVAL_2;
    end
    if (_EVAL_175) begin
      _EVAL_155 <= _EVAL;
    end
    if (_EVAL_11) begin
      _EVAL_165 <= 2'h0;
    end else begin
      _EVAL_165 <= _EVAL_307;
    end
    if (_EVAL_235) begin
      _EVAL_201 <= _EVAL_14;
    end
    if (_EVAL_175) begin
      _EVAL_276 <= _EVAL_1;
    end
    if (_EVAL_175) begin
      _EVAL_290 <= _EVAL_8;
    end
    if (_EVAL_235) begin
      _EVAL_300 <= _EVAL_17;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_325 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39f1cef3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(482088d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abff3733)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbadd8a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_325 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_325 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4402918)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b741dac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3db62be7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_265) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffdb2e9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(112e5d9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74c81c3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_325 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c6ecf8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e02022c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48f8d9c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_314 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce9ae3f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e2d1434)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d6ce7ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f05169b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_325 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(294086d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(990a428a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96104023)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3070a9f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51418ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dbd5836)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1db7cb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6858e05d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e2d3cc7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_314 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_265) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3861fca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(166ab2b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30446e5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_298) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7869b24f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97a4c842)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afbb60dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18d19b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48e1ff91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edae4cd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b562b1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d371f933)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b973059)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(947a2dc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de5b818d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_325 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7538c50c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30fe2580)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ef51a9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3067ea40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bce2d140)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3117b061)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd594426)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48402f50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c3cdb2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17edb9d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5071669a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ada9dc59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4db8e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd87f9c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3337819e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e14bb3d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48846ca1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(851239e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_298) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae3e7213)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74365aab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73dc9fb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48adebe9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63e2d7c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce496b56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be531509)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_298) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f264d4ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(291f0fa7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d85cc32a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b05448ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1375c66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_325 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2896b9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_298) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b4f8896)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5502f9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(217e219e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7e087a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ab2c7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb3c298)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_325 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
