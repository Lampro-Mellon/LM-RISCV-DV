//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_47(
  output [2:0]  _EVAL,
  input         _EVAL_0,
  output        _EVAL_1,
  output [31:0] _EVAL_2,
  output        _EVAL_3,
  output        _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  output [31:0] _EVAL_7,
  input  [3:0]  _EVAL_8,
  output        _EVAL_9,
  output        _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  output        _EVAL_13,
  input  [31:0] _EVAL_14,
  input         _EVAL_15,
  output        _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  output        _EVAL_20,
  output        _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  output        _EVAL_24,
  input         _EVAL_25,
  output [3:0]  _EVAL_26,
  output        _EVAL_27,
  output        _EVAL_28,
  input  [31:0] _EVAL_29,
  output        _EVAL_30,
  output [2:0]  _EVAL_31,
  input  [2:0]  _EVAL_32,
  output [1:0]  _EVAL_33,
  input         _EVAL_34,
  input         _EVAL_35,
  input  [3:0]  _EVAL_36,
  input  [1:0]  _EVAL_37,
  input         _EVAL_38,
  input  [3:0]  _EVAL_39,
  input         _EVAL_40,
  input  [31:0] _EVAL_41,
  input         _EVAL_42,
  output        _EVAL_43,
  output [3:0]  _EVAL_44,
  output [3:0]  _EVAL_45,
  output [31:0] _EVAL_46
);
  assign _EVAL_45 = _EVAL_39;
  assign _EVAL_16 = _EVAL_17;
  assign _EVAL_4 = _EVAL_25;
  assign _EVAL_3 = _EVAL_15;
  assign _EVAL_33 = _EVAL_37;
  assign _EVAL_13 = _EVAL_22;
  assign _EVAL_21 = _EVAL_0;
  assign _EVAL_7 = _EVAL_41;
  assign _EVAL_27 = _EVAL_6;
  assign _EVAL_30 = _EVAL_11;
  assign _EVAL_43 = _EVAL_38;
  assign _EVAL_44 = _EVAL_36;
  assign _EVAL_1 = _EVAL_42;
  assign _EVAL_24 = _EVAL_18;
  assign _EVAL = _EVAL_32;
  assign _EVAL_2 = _EVAL_14;
  assign _EVAL_46 = _EVAL_29;
  assign _EVAL_20 = _EVAL_19;
  assign _EVAL_28 = _EVAL_40;
  assign _EVAL_10 = _EVAL_23;
  assign _EVAL_31 = _EVAL_5;
  assign _EVAL_9 = _EVAL_35;
  assign _EVAL_26 = _EVAL_8;
endmodule
