//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_50(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  output        _EVAL_2,
  input         _EVAL_3,
  input  [1:0]  _EVAL_4,
  input  [31:0] _EVAL_5,
  output [2:0]  _EVAL_6,
  output        _EVAL_7,
  output [3:0]  _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  output [31:0] _EVAL_11,
  input         _EVAL_12,
  output        _EVAL_13,
  output        _EVAL_14,
  output        _EVAL_15,
  input         _EVAL_16,
  output        _EVAL_17,
  output [31:0] _EVAL_18,
  input  [31:0] _EVAL_19,
  input         _EVAL_20,
  input  [2:0]  _EVAL_21,
  output        _EVAL_22,
  output        _EVAL_23,
  output [3:0]  _EVAL_24,
  output        _EVAL_25,
  output        _EVAL_26,
  input  [3:0]  _EVAL_27,
  input  [31:0] _EVAL_28,
  output [31:0] _EVAL_29,
  input         _EVAL_30
);
  reg [31:0] _EVAL_31;
  reg [31:0] _RAND_0;
  wire  _EVAL_32;
  wire [2:0] _EVAL_33;
  wire  _EVAL_34;
  reg  _EVAL_35;
  reg [31:0] _RAND_1;
  wire [31:0] _EVAL_37;
  wire [32:0] _EVAL_38;
  wire [32:0] _EVAL_39;
  reg  _EVAL_40;
  reg [31:0] _RAND_2;
  wire  _EVAL_41;
  reg  _EVAL_43;
  reg [31:0] _RAND_3;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire [4:0] _EVAL_46;
  reg  _EVAL_47;
  reg [31:0] _RAND_4;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire [32:0] _EVAL_52;
  wire [1:0] _EVAL_53;
  wire  _EVAL_54;
  wire [32:0] _EVAL_56;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire [1:0] _EVAL_60;
  wire [5:0] _EVAL_61;
  wire  _EVAL_62;
  wire [32:0] _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire [2:0] _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire [31:0] _EVAL_75;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire [31:0] _EVAL_81;
  wire  _EVAL_82;
  wire [5:0] _EVAL_83;
  reg [31:0] _EVAL_85;
  reg [31:0] _RAND_5;
  wire  _EVAL_86;
  reg [3:0] _EVAL_88;
  reg [31:0] _RAND_6;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire [32:0] _EVAL_93;
  wire [32:0] _EVAL_94;
  wire [32:0] _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_100;
  wire [31:0] _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_106;
  wire [2:0] _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_112;
  wire  _EVAL_113;
  reg  _EVAL_114;
  reg [31:0] _RAND_7;
  wire [32:0] _EVAL_115;
  wire  _EVAL_116;
  wire [5:0] _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  reg  _EVAL_121;
  reg [31:0] _RAND_8;
  wire [32:0] _EVAL_122;
  wire [32:0] _EVAL_123;
  wire  _EVAL_124;
  reg [3:0] _EVAL_125;
  reg [31:0] _RAND_9;
  wire [2:0] _EVAL_127;
  wire  _EVAL_128;
  wire [32:0] _EVAL_131;
  wire  _EVAL_133;
  wire [32:0] _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire [3:0] _EVAL_140;
  wire  _EVAL_141;
  reg  _EVAL_142;
  reg [31:0] _RAND_10;
  wire [2:0] _EVAL_143;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire [1:0] _EVAL_151;
  wire  _EVAL_153;
  wire [5:0] _EVAL_154;
  wire [32:0] _EVAL_155;
  wire  _EVAL_156;
  wire [31:0] _EVAL_157;
  wire [1:0] _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire [2:0] _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire [31:0] _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire [32:0] _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [5:0] _EVAL_174;
  wire [31:0] _EVAL_175;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire [5:0] _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  reg  _EVAL_182;
  reg [31:0] _RAND_11;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire [32:0] _EVAL_192;
  reg  _EVAL_193;
  reg [31:0] _RAND_12;
  reg  _EVAL_196;
  reg [31:0] _RAND_13;
  wire  _EVAL_197;
  wire [3:0] _EVAL_198;
  wire  _EVAL_199;
  wire [32:0] _EVAL_200;
  reg  _EVAL_201;
  reg [31:0] _RAND_14;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire [32:0] _EVAL_204;
  wire  _EVAL_205;
  wire [2:0] _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_210;
  wire  _EVAL_212;
  assign _EVAL_134 = _EVAL_204;
  assign _EVAL_188 = _EVAL_27[0];
  assign _EVAL_13 = _EVAL_142;
  assign _EVAL_140 = _EVAL_179[5:2];
  assign _EVAL_64 = _EVAL_89 & _EVAL_68;
  assign _EVAL_181 = ~_EVAL_188;
  assign _EVAL_73 = _EVAL_4 == 2'h3;
  assign _EVAL_49 = _EVAL_31[1];
  assign _EVAL_149 = _EVAL_210 | _EVAL_73;
  assign _EVAL_24 = {_EVAL_53,_EVAL_60};
  assign _EVAL_135 = _EVAL_150 | _EVAL_58;
  assign _EVAL_68 = _EVAL_86 & _EVAL_156;
  assign _EVAL_178 = _EVAL_9 & _EVAL_100;
  assign _EVAL_18 = _EVAL_19;
  assign _EVAL_145 = _EVAL_40 ? _EVAL_65 : _EVAL_97;
  assign _EVAL_106 = $signed(_EVAL_134) == 33'sh0;
  assign _EVAL_124 = _EVAL_88 == 4'h0;
  assign _EVAL_177 = _EVAL_166 | _EVAL_106;
  assign _EVAL_78 = _EVAL_20 ? _EVAL_103 : _EVAL_103;
  assign _EVAL_147 = _EVAL_66 & _EVAL_49;
  assign _EVAL_117 = 3'h2 == _EVAL_10 ? 6'hf : 6'h3;
  assign _EVAL_133 = ~_EVAL_201;
  assign _EVAL_174 = 3'h4 == _EVAL_10 ? 6'h1f : _EVAL_61;
  assign _EVAL_17 = _EVAL_182;
  assign _EVAL_15 = _EVAL_201;
  assign _EVAL_136 = _EVAL_120 & _EVAL_121;
  assign _EVAL_109 = _EVAL_98 & _EVAL_54;
  assign _EVAL_148 = _EVAL_116 & _EVAL_79;
  assign _EVAL_169 = $signed(_EVAL_93) == 33'sh0;
  assign _EVAL_138 = _EVAL_3 & _EVAL;
  assign _EVAL_150 = ~_EVAL_20;
  assign _EVAL_167 = _EVAL_30 ? 1'h0 : _EVAL_193;
  assign _EVAL_45 = _EVAL_128 | _EVAL_64;
  assign _EVAL_123 = $signed(_EVAL_96) & -33'sh1000000;
  assign _EVAL_104 = _EVAL_197 & _EVAL_190;
  assign _EVAL_139 = _EVAL_20 ? _EVAL_92 : _EVAL_92;
  assign _EVAL_155 = {1'b0,$signed(_EVAL_175)};
  assign _EVAL_112 = $signed(_EVAL_115) == 33'sh0;
  assign _EVAL_199 = _EVAL_173 | _EVAL_172;
  assign _EVAL_207 = _EVAL_107 <= 3'h6;
  assign _EVAL_53 = {_EVAL_90,_EVAL_74};
  assign _EVAL_159 = 2'h1 << _EVAL_185;
  assign _EVAL_41 = _EVAL_34 ? 1'h0 : _EVAL_121;
  assign _EVAL_14 = _EVAL_43;
  assign _EVAL_89 = _EVAL_151[0];
  assign _EVAL_50 = _EVAL_21 == 3'h2;
  assign _EVAL_168 = _EVAL_5 ^ 32'h40000000;
  assign _EVAL_189 = _EVAL_203 | _EVAL_147;
  assign _EVAL_63 = _EVAL_122;
  assign _EVAL_202 = _EVAL_49 & _EVAL_80;
  assign _EVAL_154 = 3'h5 == _EVAL_10 ? 6'h1f : _EVAL_174;
  assign _EVAL_65 = _EVAL_110 & _EVAL_161;
  assign _EVAL_119 = _EVAL_89 & _EVAL_70;
  assign _EVAL_204 = $signed(_EVAL_39) & -33'sh5000;
  assign _EVAL_96 = {1'b0,$signed(_EVAL_157)};
  assign _EVAL_185 = _EVAL_125[0];
  assign _EVAL_161 = _EVAL_108 | _EVAL_9;
  assign _EVAL_206 = 3'h6 == _EVAL_10 ? 3'h6 : _EVAL_67;
  assign _EVAL_102 = _EVAL_27[3];
  assign _EVAL_34 = _EVAL_145 & _EVAL_120;
  assign _EVAL_128 = _EVAL_203 | _EVAL_141;
  assign _EVAL_93 = _EVAL_192;
  assign _EVAL_23 = _EVAL_196;
  assign _EVAL_90 = _EVAL_189 | _EVAL_205;
  assign _EVAL_143 = 3'h3 == _EVAL_10 ? 3'h4 : _EVAL_33;
  assign _EVAL_92 = _EVAL_71 | _EVAL_186;
  assign _EVAL_94 = _EVAL_52;
  assign _EVAL_79 = _EVAL_177 | _EVAL_186;
  assign _EVAL_69 = _EVAL_10 != 3'h1;
  assign _EVAL_83 = 3'h6 == _EVAL_10 ? 6'h3f : _EVAL_154;
  assign _EVAL_58 = _EVAL_9 ? 1'h0 : _EVAL_201;
  assign _EVAL_2 = _EVAL_193;
  assign _EVAL_25 = _EVAL_47;
  assign _EVAL_210 = _EVAL_4 == 2'h2;
  assign _EVAL_200 = {1'b0,$signed(_EVAL_75)};
  assign _EVAL_165 = ~_EVAL_193;
  assign _EVAL_203 = _EVAL_125 >= 4'h2;
  assign _EVAL_91 = _EVAL_124 & _EVAL_3;
  assign _EVAL_160 = _EVAL_89 & _EVAL_72;
  assign _EVAL_75 = _EVAL_5 ^ 32'h3000;
  assign _EVAL_37 = {{26'd0}, _EVAL_179};
  assign _EVAL_39 = {1'b0,$signed(_EVAL_5)};
  assign _EVAL_141 = _EVAL_66 & _EVAL_86;
  assign _EVAL_101 = _EVAL_5 & _EVAL_37;
  assign _EVAL_108 = _EVAL_82 | _EVAL_133;
  assign _EVAL_54 = ~_EVAL_91;
  assign _EVAL_11 = _EVAL_31;
  assign _EVAL_32 = _EVAL_27[1];
  assign _EVAL_205 = _EVAL_89 & _EVAL_202;
  assign _EVAL_52 = $signed(_EVAL_171) & -33'shc000;
  assign _EVAL_61 = 3'h3 == _EVAL_10 ? 6'hf : _EVAL_117;
  assign _EVAL_67 = 3'h5 == _EVAL_10 ? 3'h5 : _EVAL_162;
  assign _EVAL_22 = _EVAL_145 & _EVAL_163;
  assign _EVAL_162 = 3'h4 == _EVAL_10 ? 3'h5 : _EVAL_143;
  assign _EVAL_81 = _EVAL_5 ^ 32'h80000000;
  assign _EVAL_190 = ~_EVAL_139;
  assign _EVAL_198 = _EVAL_46[3:0];
  assign _EVAL_127 = _EVAL_59 ? _EVAL_107 : _EVAL_21;
  assign _EVAL_60 = {_EVAL_170,_EVAL_45};
  assign _EVAL_110 = _EVAL_165 | _EVAL_30;
  assign _EVAL_115 = _EVAL_123;
  assign _EVAL_173 = $signed(_EVAL_94) == 33'sh0;
  assign _EVAL_98 = _EVAL_114 | _EVAL_178;
  assign _EVAL_59 = _EVAL_62 & _EVAL_78;
  assign _EVAL_153 = _EVAL_124 | _EVAL_41;
  assign _EVAL_120 = _EVAL_98 & _EVAL_124;
  assign _EVAL_137 = _EVAL_109 | _EVAL_104;
  assign _EVAL_66 = _EVAL_151[1];
  assign _EVAL_6 = _EVAL_40 ? 3'h0 : 3'h4;
  assign _EVAL_175 = _EVAL_5 ^ 32'h20000000;
  assign _EVAL_186 = $signed(_EVAL_63) == 33'sh0;
  assign _EVAL_118 = _EVAL_210 & _EVAL_50;
  assign _EVAL_192 = $signed(_EVAL_200) & -33'sh1000;
  assign _EVAL_146 = _EVAL_199 | _EVAL_169;
  assign _EVAL_116 = _EVAL_107 <= 3'h2;
  assign _EVAL_33 = 3'h2 == _EVAL_10 ? 3'h4 : 3'h2;
  assign _EVAL_80 = _EVAL_31[0];
  assign _EVAL_197 = _EVAL_138 & _EVAL_149;
  assign _EVAL_71 = _EVAL_183 | _EVAL_106;
  assign _EVAL_62 = _EVAL_184 & _EVAL_69;
  assign _EVAL_163 = ~_EVAL_136;
  assign _EVAL_100 = _EVAL_12 | _EVAL_0;
  assign _EVAL_131 = _EVAL_56;
  assign _EVAL_72 = _EVAL_86 & _EVAL_80;
  assign _EVAL_113 = _EVAL_197 ? _EVAL_153 : _EVAL_41;
  assign _EVAL_86 = ~_EVAL_49;
  assign _EVAL_46 = _EVAL_88 - 4'h1;
  assign _EVAL_8 = _EVAL_125;
  assign _EVAL_44 = _EVAL_148 | _EVAL_212;
  assign _EVAL_156 = ~_EVAL_80;
  assign _EVAL_97 = _EVAL_9 | _EVAL_133;
  assign _EVAL_151 = _EVAL_159 | 2'h1;
  assign _EVAL_170 = _EVAL_128 | _EVAL_160;
  assign _EVAL_184 = _EVAL_118 & _EVAL_187;
  assign _EVAL_183 = _EVAL_146 | _EVAL_112;
  assign _EVAL_122 = $signed(_EVAL_155) & -33'sh2000;
  assign _EVAL_157 = _EVAL_5 ^ 32'h2000000;
  assign _EVAL_56 = $signed(_EVAL_38) & -33'sh2000;
  assign _EVAL_103 = _EVAL_44 | _EVAL_169;
  assign _EVAL_172 = $signed(_EVAL_131) == 33'sh0;
  assign _EVAL_171 = {1'b0,$signed(_EVAL_81)};
  assign _EVAL_191 = _EVAL_27[2];
  assign _EVAL_29 = _EVAL_201 ? _EVAL_28 : _EVAL_85;
  assign _EVAL_180 = _EVAL_20 | _EVAL_167;
  assign _EVAL_26 = _EVAL_35;
  assign _EVAL_107 = 3'h7 == _EVAL_10 ? 3'h6 : _EVAL_206;
  assign _EVAL_7 = _EVAL_145 & _EVAL_120;
  assign _EVAL_212 = _EVAL_207 & _EVAL_172;
  assign _EVAL_166 = _EVAL_173 | _EVAL_112;
  assign _EVAL_179 = 3'h7 == _EVAL_10 ? 6'h3f : _EVAL_83;
  assign _EVAL_38 = {1'b0,$signed(_EVAL_168)};
  assign _EVAL_82 = ~_EVAL_124;
  assign _EVAL_70 = _EVAL_49 & _EVAL_156;
  assign _EVAL_187 = _EVAL_101 == 32'h0;
  assign _EVAL_74 = _EVAL_189 | _EVAL_119;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_31 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_35 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_40 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_43 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_47 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_85 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_88 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_114 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_121 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_125 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_142 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_182 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_193 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_196 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_201 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_16) begin
    if (_EVAL_197) begin
      if (_EVAL_124) begin
        _EVAL_31 <= _EVAL_5;
      end
    end
    if (_EVAL_197) begin
      if (_EVAL_124) begin
        _EVAL_35 <= _EVAL_181;
      end
    end
    if (_EVAL_1) begin
      _EVAL_40 <= 1'h0;
    end else if (_EVAL_197) begin
      if (_EVAL_124) begin
        _EVAL_40 <= _EVAL_20;
      end
    end
    if (_EVAL_197) begin
      if (_EVAL_124) begin
        _EVAL_43 <= _EVAL_32;
      end
    end
    if (_EVAL_197) begin
      if (_EVAL_124) begin
        _EVAL_47 <= _EVAL_102;
      end
    end
    if (_EVAL_201) begin
      _EVAL_85 <= _EVAL_28;
    end
    if (_EVAL_1) begin
      _EVAL_88 <= 4'h0;
    end else if (_EVAL_197) begin
      if (_EVAL_124) begin
        if (_EVAL_59) begin
          _EVAL_88 <= _EVAL_140;
        end else begin
          _EVAL_88 <= 4'h0;
        end
      end else begin
        _EVAL_88 <= _EVAL_198;
      end
    end
    if (_EVAL_1) begin
      _EVAL_114 <= 1'h0;
    end else begin
      _EVAL_114 <= _EVAL_137;
    end
    _EVAL_121 <= _EVAL_1 | _EVAL_113;
    if (_EVAL_197) begin
      if (_EVAL_124) begin
        _EVAL_125 <= {{1'd0}, _EVAL_127};
      end
    end
    if (_EVAL_197) begin
      if (_EVAL_124) begin
        _EVAL_142 <= _EVAL_102;
      end
    end
    if (_EVAL_197) begin
      if (_EVAL_124) begin
        _EVAL_182 <= _EVAL_191;
      end
    end
    if (_EVAL_1) begin
      _EVAL_193 <= 1'h0;
    end else if (_EVAL_197) begin
      if (_EVAL_124) begin
        if (_EVAL_20) begin
          _EVAL_193 <= _EVAL_92;
        end else begin
          _EVAL_193 <= _EVAL_92;
        end
      end else begin
        _EVAL_193 <= _EVAL_180;
      end
    end else if (_EVAL_30) begin
      _EVAL_193 <= 1'h0;
    end
    if (_EVAL_197) begin
      if (_EVAL_124) begin
        _EVAL_196 <= _EVAL_102;
      end
    end
    if (_EVAL_1) begin
      _EVAL_201 <= 1'h0;
    end else if (_EVAL_197) begin
      if (_EVAL_124) begin
        if (_EVAL_20) begin
          _EVAL_201 <= _EVAL_92;
        end else begin
          _EVAL_201 <= _EVAL_92;
        end
      end else begin
        _EVAL_201 <= _EVAL_135;
      end
    end else if (_EVAL_9) begin
      _EVAL_201 <= 1'h0;
    end
  end
endmodule
