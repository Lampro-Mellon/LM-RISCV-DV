//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_138_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input  [3:0]  _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [1:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input  [11:0] _EVAL_8,
  input  [1:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [2:0]  _EVAL_14
);
  wire [7:0] _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire [4:0] _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  reg [2:0] _EVAL_51;
  reg [31:0] _RAND_0;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  reg [1:0] _EVAL_69;
  reg [31:0] _RAND_1;
  reg  _EVAL_70;
  reg [31:0] _RAND_2;
  wire  _EVAL_71;
  wire [1:0] _EVAL_72;
  wire  _EVAL_73;
  wire [12:0] _EVAL_74;
  wire  _EVAL_75;
  wire [3:0] _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  reg  _EVAL_79;
  reg [31:0] _RAND_3;
  wire [12:0] _EVAL_80;
  reg [2:0] _EVAL_81;
  reg [31:0] _RAND_4;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_95;
  wire [7:0] _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire [4:0] _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire [4:0] _EVAL_105;
  reg [31:0] _EVAL_106;
  reg [31:0] _RAND_5;
  wire [7:0] _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  reg  _EVAL_121;
  reg [31:0] _RAND_6;
  wire  _EVAL_122;
  wire [1:0] _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  reg [2:0] _EVAL_127;
  reg [31:0] _RAND_7;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire [4:0] _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire [12:0] _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire [3:0] _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire [1:0] _EVAL_157;
  wire [4:0] _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire [1:0] _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire [11:0] _EVAL_166;
  wire  _EVAL_167;
  wire [3:0] _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire [4:0] _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [4:0] _EVAL_174;
  wire  _EVAL_175;
  wire [1:0] _EVAL_176;
  wire  _EVAL_177;
  wire [7:0] _EVAL_178;
  wire [4:0] _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire [11:0] _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire [1:0] _EVAL_195;
  wire  _EVAL_196;
  reg [1:0] _EVAL_197;
  reg [31:0] _RAND_8;
  reg [11:0] _EVAL_198;
  reg [31:0] _RAND_9;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire [3:0] _EVAL_202;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_203;
  wire [1:0] _EVAL_204;
  wire  _EVAL_205;
  wire [1:0] _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire [32:0] _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  reg [4:0] _EVAL_219;
  reg [31:0] _RAND_10;
  wire [31:0] _EVAL_220;
  wire  _EVAL_222;
  reg [2:0] _EVAL_223;
  reg [31:0] _RAND_11;
  wire  _EVAL_224;
  reg  _EVAL_225;
  reg [31:0] _RAND_12;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  reg [2:0] _EVAL_233;
  reg [31:0] _RAND_13;
  wire [4:0] _EVAL_234;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_202 = ~_EVAL_168;
  assign _EVAL_186 = _EVAL_9 == _EVAL_197;
  assign _EVAL_97 = _EVAL_110 & _EVAL_36;
  assign _EVAL_183 = _EVAL_55 | _EVAL_1;
  assign _EVAL_19 = _EVAL_0 & _EVAL_213;
  assign _EVAL_192 = _EVAL_34 & _EVAL_122;
  assign _EVAL_72 = _EVAL_79 - 1'h1;
  assign _EVAL_130 = _EVAL_106 < plusarg_reader_out;
  assign _EVAL_199 = _EVAL_156 | _EVAL_1;
  assign _EVAL_133 = _EVAL_187 == 12'h0;
  assign _EVAL_187 = _EVAL_8 & _EVAL_166;
  assign _EVAL_65 = _EVAL_186 | _EVAL_1;
  assign _EVAL_63 = _EVAL_8 == _EVAL_198;
  assign _EVAL_228 = _EVAL_0 & _EVAL_230;
  assign _EVAL_68 = _EVAL_6 == 3'h1;
  assign _EVAL_135 = ~_EVAL_67;
  assign _EVAL_115 = _EVAL & _EVAL_182;
  assign _EVAL_62 = _EVAL_208 | _EVAL_1;
  assign _EVAL_60 = _EVAL_17 | _EVAL_1;
  assign _EVAL_209 = _EVAL_6 == _EVAL_51;
  assign _EVAL_131 = ~_EVAL_46;
  assign _EVAL_194 = _EVAL_47 | _EVAL_1;
  assign _EVAL_215 = ~_EVAL_175;
  assign _EVAL_191 = _EVAL_14 == 3'h7;
  assign _EVAL_208 = _EVAL_76 == 4'h0;
  assign _EVAL_124 = _EVAL & _EVAL_229;
  assign _EVAL_76 = _EVAL_3 & _EVAL_202;
  assign _EVAL_31 = _EVAL_111 | _EVAL_1;
  assign _EVAL_140 = ~_EVAL_121;
  assign _EVAL_15 = _EVAL_172 ? _EVAL_96 : 8'h0;
  assign _EVAL_29 = _EVAL_14 == 3'h6;
  assign _EVAL_87 = _EVAL_0 & _EVAL_160;
  assign _EVAL_44 = _EVAL_119 | _EVAL_1;
  assign _EVAL_46 = _EVAL_89 | _EVAL_1;
  assign _EVAL_85 = _EVAL_63 | _EVAL_1;
  assign _EVAL_216 = _EVAL_34 & _EVAL_181;
  assign _EVAL_145 = _EVAL_210 | _EVAL_1;
  assign _EVAL_102 = _EVAL_0 & _EVAL_214;
  assign _EVAL_195 = ~_EVAL_206;
  assign _EVAL_160 = _EVAL_6 == 3'h5;
  assign _EVAL_201 = _EVAL_54 | _EVAL_1;
  assign _EVAL_189 = ~_EVAL_141;
  assign _EVAL_107 = _EVAL_18 ? _EVAL_178 : 8'h0;
  assign _EVAL_99 = _EVAL_72[0];
  assign _EVAL_59 = _EVAL_118 | _EVAL_190;
  assign _EVAL_105 = _EVAL_219 >> _EVAL_4;
  assign _EVAL_18 = _EVAL_118 & _EVAL_73;
  assign _EVAL_210 = _EVAL_9 >= 2'h2;
  assign _EVAL_41 = _EVAL_219 | _EVAL_171;
  assign _EVAL_98 = ~_EVAL_112;
  assign _EVAL_205 = ~_EVAL_231;
  assign _EVAL_226 = ~_EVAL_36;
  assign _EVAL_89 = _EVAL_10 <= 3'h4;
  assign _EVAL_161 = _EVAL_6 == 3'h2;
  assign _EVAL_17 = ~_EVAL_7;
  assign _EVAL_206 = _EVAL_179[1:0];
  assign _EVAL_134 = _EVAL_48 | _EVAL_1;
  assign _EVAL_32 = _EVAL_226 & _EVAL_112;
  assign _EVAL_185 = _EVAL_154 == 4'h0;
  assign _EVAL_148 = ~_EVAL_31;
  assign _EVAL_188 = ~_EVAL_193;
  assign _EVAL_212 = ~_EVAL_199;
  assign _EVAL_21 = _EVAL_190 & _EVAL_30;
  assign _EVAL_167 = _EVAL_204[0];
  assign _EVAL_163 = plusarg_reader_out == 32'h0;
  assign _EVAL_159 = _EVAL_0 & _EVAL_161;
  assign _EVAL_157 = _EVAL_123 | 2'h1;
  assign _EVAL_179 = 5'h3 << _EVAL_5;
  assign _EVAL_38 = ~_EVAL_214;
  assign _EVAL_214 = _EVAL_6 == 3'h6;
  assign _EVAL_24 = _EVAL_162[0];
  assign _EVAL_39 = _EVAL_4 <= 3'h4;
  assign _EVAL_64 = ~_EVAL_95;
  assign _EVAL_173 = _EVAL_4 == _EVAL_81;
  assign _EVAL_231 = _EVAL_113 | _EVAL_1;
  assign _EVAL_28 = _EVAL_3 == _EVAL_168;
  assign _EVAL_36 = _EVAL_8[1];
  assign _EVAL_103 = ~_EVAL_136;
  assign _EVAL_182 = ~_EVAL_140;
  assign _EVAL_58 = _EVAL_14 == 3'h1;
  assign _EVAL_77 = ~_EVAL_70;
  assign _EVAL_139 = _EVAL_15[4:0];
  assign _EVAL_126 = _EVAL_190 & _EVAL_77;
  assign _EVAL_35 = _EVAL_105[0];
  assign _EVAL_166 = {{10'd0}, _EVAL_195};
  assign _EVAL_75 = ~_EVAL_201;
  assign _EVAL_23 = _EVAL_113 | _EVAL_117;
  assign _EVAL_213 = ~_EVAL_30;
  assign _EVAL_203 = ~_EVAL_134;
  assign _EVAL_67 = _EVAL_39 | _EVAL_1;
  assign _EVAL_55 = _EVAL_10 == _EVAL_223;
  assign _EVAL_80 = $signed(_EVAL_147) & -13'sh1000;
  assign _EVAL_143 = ~_EVAL_37;
  assign _EVAL_196 = _EVAL_152 | _EVAL_1;
  assign _EVAL_48 = _EVAL_174[0];
  assign _EVAL_96 = 8'h1 << _EVAL_11;
  assign _EVAL_170 = _EVAL_50 | _EVAL_1;
  assign _EVAL_227 = ~_EVAL_232;
  assign _EVAL_144 = _EVAL_0 & _EVAL_68;
  assign _EVAL_155 = _EVAL & _EVAL_93;
  assign _EVAL_177 = ~_EVAL_170;
  assign _EVAL_138 = _EVAL_6 == 3'h0;
  assign _EVAL_169 = ~_EVAL_60;
  assign _EVAL_22 = ~_EVAL_62;
  assign _EVAL_112 = _EVAL_8[0];
  assign _EVAL_217 = _EVAL & _EVAL_66;
  assign _EVAL_27 = ~_EVAL_1;
  assign _EVAL_104 = _EVAL_209 | _EVAL_1;
  assign _EVAL_88 = _EVAL_14 == 3'h2;
  assign _EVAL_54 = _EVAL_10 == 3'h0;
  assign _EVAL_172 = _EVAL_126 & _EVAL_38;
  assign _EVAL_34 = _EVAL_157[0];
  assign _EVAL_175 = _EVAL_219 != 5'h0;
  assign _EVAL_152 = _EVAL_11 <= 3'h4;
  assign _EVAL_73 = ~_EVAL_225;
  assign _EVAL_114 = _EVAL_132 | _EVAL_216;
  assign _EVAL_150 = _EVAL_34 & _EVAL_32;
  assign _EVAL_119 = _EVAL_10 != 3'h0;
  assign _EVAL_146 = _EVAL_34 & _EVAL_200;
  assign _EVAL_43 = _EVAL_132 | _EVAL_146;
  assign _EVAL_117 = _EVAL_110 & _EVAL_226;
  assign _EVAL_132 = _EVAL_113 | _EVAL_97;
  assign _EVAL_193 = _EVAL_218 | _EVAL_1;
  assign _EVAL_234 = _EVAL_171 | _EVAL_219;
  assign _EVAL_57 = _EVAL_165 | _EVAL_1;
  assign _EVAL_52 = _EVAL & _EVAL_29;
  assign _EVAL_180 = ~_EVAL_44;
  assign _EVAL_125 = _EVAL_11 == _EVAL_233;
  assign _EVAL_53 = _EVAL_6 <= 3'h6;
  assign _EVAL_142 = $signed(_EVAL_74) == 13'sh0;
  assign _EVAL_74 = _EVAL_80;
  assign _EVAL_56 = _EVAL_5[0];
  assign _EVAL_66 = _EVAL_14 == 3'h5;
  assign _EVAL_151 = _EVAL_176[0];
  assign _EVAL_92 = ~_EVAL_40;
  assign _EVAL_122 = _EVAL_226 & _EVAL_98;
  assign _EVAL_147 = {1'b0,$signed(_EVAL_8)};
  assign _EVAL_84 = ~_EVAL_196;
  assign _EVAL_232 = _EVAL_133 | _EVAL_1;
  assign _EVAL_181 = _EVAL_36 & _EVAL_98;
  assign _EVAL_111 = _EVAL_10 <= 3'h2;
  assign _EVAL_128 = ~_EVAL_57;
  assign _EVAL_118 = _EVAL_12 & _EVAL;
  assign _EVAL_141 = _EVAL_53 | _EVAL_1;
  assign _EVAL_211 = _EVAL_106 + 32'h1;
  assign _EVAL_158 = _EVAL_41 & _EVAL_100;
  assign _EVAL_42 = _EVAL & _EVAL_88;
  assign _EVAL_61 = _EVAL_0 & _EVAL_138;
  assign _EVAL_224 = _EVAL_10 <= 3'h3;
  assign _EVAL_49 = _EVAL_224 | _EVAL_1;
  assign _EVAL_220 = _EVAL_211[31:0];
  assign _EVAL_113 = _EVAL_5 >= 2'h2;
  assign _EVAL_47 = _EVAL_10 <= 3'h1;
  assign _EVAL_149 = _EVAL_23 | _EVAL_192;
  assign _EVAL_222 = _EVAL_215 | _EVAL_163;
  assign _EVAL_230 = _EVAL_6 == 3'h4;
  assign _EVAL_136 = _EVAL_86 | _EVAL_1;
  assign _EVAL_86 = _EVAL_5 == _EVAL_69;
  assign _EVAL_171 = _EVAL_107[4:0];
  assign _EVAL_30 = ~_EVAL_79;
  assign _EVAL_90 = _EVAL & _EVAL_137;
  assign _EVAL_101 = ~_EVAL_65;
  assign _EVAL_156 = _EVAL_14 == _EVAL_127;
  assign _EVAL_108 = ~_EVAL_183;
  assign _EVAL_204 = _EVAL_121 - 1'h1;
  assign _EVAL_109 = ~_EVAL_145;
  assign _EVAL_165 = _EVAL_222 | _EVAL_130;
  assign _EVAL_200 = _EVAL_36 & _EVAL_112;
  assign _EVAL_162 = _EVAL_70 - 1'h1;
  assign _EVAL_176 = _EVAL_225 - 1'h1;
  assign _EVAL_33 = _EVAL_5 <= 2'h2;
  assign _EVAL_110 = _EVAL_157[1];
  assign _EVAL_178 = 8'h1 << _EVAL_4;
  assign _EVAL_50 = _EVAL_33 & _EVAL_142;
  assign _EVAL_100 = ~_EVAL_139;
  assign _EVAL_207 = _EVAL_173 | _EVAL_1;
  assign _EVAL_71 = ~_EVAL_49;
  assign _EVAL_229 = _EVAL_14 == 3'h3;
  assign _EVAL_153 = ~_EVAL_85;
  assign _EVAL_218 = ~_EVAL_35;
  assign _EVAL_116 = _EVAL_23 | _EVAL_150;
  assign _EVAL_129 = ~_EVAL_104;
  assign _EVAL_154 = ~_EVAL_3;
  assign _EVAL_16 = _EVAL & _EVAL_191;
  assign _EVAL_93 = _EVAL_14 == 3'h0;
  assign _EVAL_95 = _EVAL_28 | _EVAL_1;
  assign _EVAL_168 = {_EVAL_43,_EVAL_114,_EVAL_116,_EVAL_149};
  assign _EVAL_83 = _EVAL & _EVAL_58;
  assign _EVAL_82 = ~_EVAL_194;
  assign _EVAL_78 = ~_EVAL_207;
  assign _EVAL_37 = _EVAL_185 | _EVAL_1;
  assign _EVAL_123 = 2'h1 << _EVAL_56;
  assign _EVAL_174 = _EVAL_234 >> _EVAL_11;
  assign _EVAL_40 = _EVAL_125 | _EVAL_1;
  assign _EVAL_137 = _EVAL_14 == 3'h4;
  assign _EVAL_190 = _EVAL_2 & _EVAL_0;
  assign _EVAL_164 = _EVAL_118 & _EVAL_140;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_51 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_69 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_70 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_79 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_81 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_106 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_121 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_127 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_197 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_198 = _RAND_9[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_219 = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_223 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_225 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_233 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_13) begin
    if (_EVAL_21) begin
      _EVAL_51 <= _EVAL_6;
    end
    if (_EVAL_164) begin
      _EVAL_69 <= _EVAL_5;
    end
    if (_EVAL_1) begin
      _EVAL_70 <= 1'h0;
    end else if (_EVAL_190) begin
      if (_EVAL_77) begin
        _EVAL_70 <= 1'h0;
      end else begin
        _EVAL_70 <= _EVAL_24;
      end
    end
    if (_EVAL_1) begin
      _EVAL_79 <= 1'h0;
    end else if (_EVAL_190) begin
      if (_EVAL_30) begin
        _EVAL_79 <= 1'h0;
      end else begin
        _EVAL_79 <= _EVAL_99;
      end
    end
    if (_EVAL_164) begin
      _EVAL_81 <= _EVAL_4;
    end
    if (_EVAL_1) begin
      _EVAL_106 <= 32'h0;
    end else if (_EVAL_59) begin
      _EVAL_106 <= 32'h0;
    end else begin
      _EVAL_106 <= _EVAL_220;
    end
    if (_EVAL_1) begin
      _EVAL_121 <= 1'h0;
    end else if (_EVAL_118) begin
      if (_EVAL_140) begin
        _EVAL_121 <= 1'h0;
      end else begin
        _EVAL_121 <= _EVAL_167;
      end
    end
    if (_EVAL_164) begin
      _EVAL_127 <= _EVAL_14;
    end
    if (_EVAL_21) begin
      _EVAL_197 <= _EVAL_9;
    end
    if (_EVAL_164) begin
      _EVAL_198 <= _EVAL_8;
    end
    if (_EVAL_1) begin
      _EVAL_219 <= 5'h0;
    end else begin
      _EVAL_219 <= _EVAL_158;
    end
    if (_EVAL_164) begin
      _EVAL_223 <= _EVAL_10;
    end
    if (_EVAL_1) begin
      _EVAL_225 <= 1'h0;
    end else if (_EVAL_118) begin
      if (_EVAL_73) begin
        _EVAL_225 <= 1'h0;
      end else begin
        _EVAL_225 <= _EVAL_151;
      end
    end
    if (_EVAL_21) begin
      _EVAL_233 <= _EVAL_11;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3af92aae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c943f913)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11e5814e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69f4adda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(848d37b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94aad787)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18d188ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0357842)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c47af12d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e690a16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cbbe0c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d3333a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2156a9be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f06fa14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4c1c52d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(509e3633)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a48db70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8970a7b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df7cb923)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c010461d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23e7e767)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68195bef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c11f71ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(829c30e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b36470a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(203c3edb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8287bf90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf9ee803)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84a8df5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17ece8c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a52153a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3dcd14b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdf186ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e310a22d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4c60e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f0f5694)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(450bacda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88809ebf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e58db3d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0e1ccf7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9da9db35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(505027c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a8802aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(381b4134)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ea145a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b8648e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48d8d4bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e95a6cab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8586e4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9cfda6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac0a7aa4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebb55527)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3d2de44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef1480bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f75fe505)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dde5043b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61265ebe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee0cf295)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69709334)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9913cd59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c9317b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf7bcbe1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26ff04e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce7735a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cde716c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b90473e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f7edc10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ebe3b94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(819f45b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ce5b256)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a33173e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df99b32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
