//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_83_assert(
  input         _EVAL,
  input  [29:0] _EVAL_0,
  input  [3:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input  [1:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [1:0]  _EVAL_12,
  input         _EVAL_13,
  input  [1:0]  _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18
);
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  reg [2:0] _EVAL_32;
  reg [31:0] _RAND_0;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire [4:0] _EVAL_43;
  reg  _EVAL_44;
  reg [31:0] _RAND_1;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  reg [2:0] _EVAL_50;
  reg [31:0] _RAND_2;
  wire  _EVAL_51;
  wire [4:0] _EVAL_52;
  wire  _EVAL_53;
  reg [2:0] _EVAL_54;
  reg [31:0] _RAND_3;
  wire [30:0] _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire [3:0] _EVAL_58;
  wire [4:0] _EVAL_60;
  wire  _EVAL_61;
  wire [29:0] _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  reg [2:0] _EVAL_69;
  reg [31:0] _RAND_4;
  wire  _EVAL_71;
  wire  _EVAL_72;
  reg  _EVAL_73;
  reg [31:0] _RAND_5;
  wire [4:0] _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire [3:0] _EVAL_92;
  wire [29:0] _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire [1:0] _EVAL_102;
  wire [31:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire [3:0] _EVAL_117;
  wire  _EVAL_118;
  wire [1:0] _EVAL_119;
  wire  _EVAL_120;
  wire [4:0] _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire [4:0] _EVAL_135;
  wire  _EVAL_136;
  wire [3:0] _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  reg  _EVAL_142;
  reg [31:0] _RAND_6;
  wire  _EVAL_143;
  reg [4:0] _EVAL_144;
  reg [31:0] _RAND_7;
  wire  _EVAL_145;
  wire [32:0] _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  reg  _EVAL_152;
  reg [31:0] _RAND_8;
  reg [29:0] _EVAL_153;
  reg [31:0] _RAND_9;
  wire  _EVAL_154;
  reg [1:0] _EVAL_155;
  reg [31:0] _RAND_10;
  wire  _EVAL_156;
  wire [1:0] _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  reg [31:0] _EVAL_165;
  reg [31:0] _RAND_11;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  reg [1:0] _EVAL_170;
  reg [31:0] _RAND_12;
  wire  _EVAL_171;
  wire [4:0] _EVAL_172;
  wire  _EVAL_173;
  wire [1:0] _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire [30:0] _EVAL_186;
  wire [7:0] _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  reg [1:0] _EVAL_191;
  reg [31:0] _RAND_13;
  wire [29:0] _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire [1:0] _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_201;
  wire [7:0] _EVAL_202;
  wire  _EVAL_203;
  wire [1:0] _EVAL_204;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire [7:0] _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire [7:0] _EVAL_230;
  wire  _EVAL_232;
  reg  _EVAL_233;
  reg [31:0] _RAND_14;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire [1:0] _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  reg  _EVAL_249;
  reg [31:0] _RAND_15;
  wire [30:0] _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire [4:0] _EVAL_255;
  wire  _EVAL_256;
  wire [4:0] _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire [1:0] _EVAL_261;
  reg [2:0] _EVAL_262;
  reg [31:0] _RAND_16;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_90 = _EVAL_14 == _EVAL_170;
  assign _EVAL_171 = _EVAL_131 | _EVAL_217;
  assign _EVAL_218 = _EVAL_2 == 3'h1;
  assign _EVAL_25 = ~_EVAL_265;
  assign _EVAL_227 = ~_EVAL_147;
  assign _EVAL_270 = _EVAL_35 | _EVAL_13;
  assign _EVAL_180 = $signed(_EVAL_250) == 31'sh0;
  assign _EVAL_132 = _EVAL_148 | _EVAL_13;
  assign _EVAL_157 = _EVAL_119 | 2'h1;
  assign _EVAL_151 = _EVAL_60[0];
  assign _EVAL_87 = _EVAL_8 != 2'h2;
  assign _EVAL_101 = _EVAL_5 & _EVAL_30;
  assign _EVAL_42 = _EVAL_157[0];
  assign _EVAL_100 = ~_EVAL_95;
  assign _EVAL_75 = ~_EVAL_72;
  assign _EVAL_193 = _EVAL_264 | _EVAL_13;
  assign _EVAL_267 = ~_EVAL_244;
  assign _EVAL_222 = ~_EVAL_78;
  assign _EVAL_226 = _EVAL_87 | _EVAL_13;
  assign _EVAL_33 = _EVAL_9 <= 3'h1;
  assign _EVAL_137 = {_EVAL_37,_EVAL_177,_EVAL_167,_EVAL_237};
  assign _EVAL_186 = {1'b0,$signed(_EVAL_192)};
  assign _EVAL_49 = ~_EVAL_161;
  assign _EVAL_248 = _EVAL_134 | _EVAL_13;
  assign _EVAL_35 = ~_EVAL_7;
  assign _EVAL_220 = _EVAL_16 & _EVAL_218;
  assign _EVAL_234 = _EVAL_12 == _EVAL_155;
  assign _EVAL_79 = ~_EVAL_76;
  assign _EVAL_95 = ~_EVAL_152;
  assign _EVAL_23 = ~_EVAL_142;
  assign _EVAL_173 = ~_EVAL_226;
  assign _EVAL_258 = ~_EVAL_246;
  assign _EVAL_114 = _EVAL_33 | _EVAL_13;
  assign _EVAL_145 = _EVAL_0 == _EVAL_153;
  assign _EVAL_96 = ~_EVAL;
  assign _EVAL_111 = ~_EVAL_245;
  assign _EVAL_268 = _EVAL_4 <= 3'h4;
  assign _EVAL_252 = ~_EVAL_207;
  assign _EVAL_138 = _EVAL_165 < plusarg_reader_out;
  assign _EVAL_65 = _EVAL_247 & _EVAL_180;
  assign _EVAL_275 = _EVAL_145 | _EVAL_13;
  assign _EVAL_41 = _EVAL_94 | _EVAL_66;
  assign _EVAL_146 = _EVAL_165 + 32'h1;
  assign _EVAL_235 = ~_EVAL_127;
  assign _EVAL_163 = _EVAL_62 == 30'h0;
  assign _EVAL_149 = _EVAL_144 != 5'h0;
  assign _EVAL_202 = _EVAL_38 ? _EVAL_230 : 8'h0;
  assign _EVAL_117 = ~_EVAL_1;
  assign _EVAL_62 = _EVAL_0 & _EVAL_93;
  assign _EVAL_47 = ~_EVAL_208;
  assign _EVAL_198 = ~_EVAL_29;
  assign _EVAL_221 = _EVAL_92 == 4'h0;
  assign _EVAL_166 = _EVAL_26 | _EVAL_13;
  assign _EVAL_21 = _EVAL_8 == 2'h0;
  assign _EVAL_201 = _EVAL_3 <= 3'h6;
  assign _EVAL_72 = _EVAL_163 | _EVAL_13;
  assign _EVAL_58 = ~_EVAL_137;
  assign _EVAL_236 = _EVAL_73 - 1'h1;
  assign _EVAL_27 = ~_EVAL_139;
  assign _EVAL_78 = _EVAL_110 | _EVAL_13;
  assign _EVAL_123 = _EVAL_135 != 5'h0;
  assign _EVAL_128 = _EVAL_104 & _EVAL_95;
  assign _EVAL_129 = _EVAL_51 | _EVAL_13;
  assign _EVAL_83 = ~_EVAL_115;
  assign _EVAL_224 = _EVAL_64 | _EVAL_13;
  assign _EVAL_31 = _EVAL_16 & _EVAL_91;
  assign _EVAL_175 = ~_EVAL_13;
  assign _EVAL_164 = _EVAL_42 & _EVAL_241;
  assign _EVAL_273 = _EVAL_2 == 3'h7;
  assign _EVAL_159 = _EVAL_199 | _EVAL_13;
  assign _EVAL_245 = _EVAL_196 | _EVAL_13;
  assign _EVAL_55 = $signed(_EVAL_186) & -31'sh2000;
  assign _EVAL_259 = ~_EVAL_143;
  assign _EVAL_274 = _EVAL_151 | _EVAL_13;
  assign _EVAL_29 = _EVAL_154 | _EVAL_13;
  assign _EVAL_206 = _EVAL_204[0];
  assign _EVAL_160 = _EVAL_5 & _EVAL_195;
  assign _EVAL_104 = _EVAL_10 & _EVAL_5;
  assign _EVAL_84 = ~_EVAL_251;
  assign _EVAL_169 = _EVAL_9 != 3'h0;
  assign _EVAL_110 = _EVAL_9 <= 3'h3;
  assign _EVAL_39 = _EVAL_238 & _EVAL_139;
  assign _EVAL_214 = _EVAL_20 | _EVAL_13;
  assign _EVAL_56 = ~_EVAL_132;
  assign _EVAL_20 = _EVAL_6 == _EVAL_54;
  assign _EVAL_188 = _EVAL_158 | _EVAL_13;
  assign _EVAL_246 = _EVAL_74[0];
  assign _EVAL_30 = _EVAL_3 == 3'h2;
  assign _EVAL_197 = _EVAL_233 - 1'h1;
  assign _EVAL_210 = _EVAL_98 | _EVAL_13;
  assign _EVAL_134 = _EVAL_1 == _EVAL_137;
  assign _EVAL_141 = _EVAL_2 == 3'h4;
  assign _EVAL_229 = ~_EVAL_68;
  assign _EVAL_182 = ~_EVAL_193;
  assign _EVAL_36 = _EVAL_80 | _EVAL_13;
  assign _EVAL_130 = _EVAL_183 & _EVAL_22;
  assign _EVAL_269 = _EVAL_252 & _EVAL_79;
  assign _EVAL_103 = _EVAL_146[31:0];
  assign _EVAL_237 = _EVAL_133 | _EVAL_48;
  assign _EVAL_119 = 2'h1 << _EVAL_86;
  assign _EVAL_161 = _EVAL_21 | _EVAL_13;
  assign _EVAL_51 = _EVAL_18 == _EVAL_249;
  assign _EVAL_116 = ~_EVAL_123;
  assign _EVAL_241 = _EVAL_207 & _EVAL_79;
  assign _EVAL_168 = ~_EVAL_270;
  assign _EVAL_194 = _EVAL_16 & _EVAL_27;
  assign _EVAL_232 = _EVAL_3 == 3'h1;
  assign _EVAL_176 = _EVAL_2 == 3'h6;
  assign _EVAL_260 = _EVAL_5 & _EVAL_81;
  assign _EVAL_225 = _EVAL_238 | _EVAL_104;
  assign _EVAL_243 = _EVAL_157[1];
  assign _EVAL_86 = _EVAL_12[0];
  assign _EVAL_213 = _EVAL_3 == 3'h5;
  assign _EVAL_257 = _EVAL_135 | _EVAL_144;
  assign _EVAL_211 = _EVAL_42 & _EVAL_89;
  assign _EVAL_172 = ~_EVAL_121;
  assign _EVAL_122 = _EVAL_16 & _EVAL_53;
  assign _EVAL_216 = _EVAL_16 & _EVAL_176;
  assign _EVAL_77 = _EVAL_24 | _EVAL_13;
  assign _EVAL_271 = _EVAL_201 | _EVAL_13;
  assign _EVAL_184 = _EVAL_117 == 4'h0;
  assign _EVAL_261 = ~_EVAL_174;
  assign _EVAL_205 = _EVAL_3 == 3'h4;
  assign _EVAL_52 = 5'h3 << _EVAL_12;
  assign _EVAL_208 = _EVAL_190 | _EVAL_13;
  assign _EVAL_192 = _EVAL_0 ^ 30'h20000000;
  assign _EVAL_125 = _EVAL_105 | _EVAL_13;
  assign _EVAL_190 = _EVAL_97 | _EVAL_116;
  assign _EVAL_150 = ~_EVAL_214;
  assign _EVAL_80 = _EVAL_9 <= 3'h4;
  assign _EVAL_81 = _EVAL_3 == 3'h0;
  assign _EVAL_148 = _EVAL_3 == _EVAL_69;
  assign _EVAL_256 = _EVAL_169 | _EVAL_13;
  assign _EVAL_266 = ~_EVAL_275;
  assign _EVAL_185 = _EVAL_5 & _EVAL_205;
  assign _EVAL_179 = _EVAL_9 <= 3'h2;
  assign _EVAL_238 = _EVAL_11 & _EVAL_16;
  assign _EVAL_228 = ~_EVAL_188;
  assign _EVAL_209 = _EVAL_162 | _EVAL_13;
  assign _EVAL_131 = _EVAL_12 >= 2'h2;
  assign _EVAL_102 = _EVAL_152 - 1'h1;
  assign _EVAL_26 = _EVAL_9 == _EVAL_32;
  assign _EVAL_223 = ~_EVAL_274;
  assign _EVAL_133 = _EVAL_131 | _EVAL_112;
  assign _EVAL_143 = _EVAL_90 | _EVAL_13;
  assign _EVAL_48 = _EVAL_42 & _EVAL_269;
  assign _EVAL_68 = _EVAL_258 | _EVAL_13;
  assign _EVAL_40 = ~_EVAL_256;
  assign _EVAL_24 = _EVAL_4 == _EVAL_50;
  assign _EVAL_212 = _EVAL_207 & _EVAL_76;
  assign _EVAL_57 = _EVAL_16 & _EVAL_273;
  assign _EVAL_94 = ~_EVAL_149;
  assign _EVAL_85 = ~_EVAL_63;
  assign _EVAL_250 = _EVAL_55;
  assign _EVAL_219 = ~_EVAL_248;
  assign _EVAL_272 = ~_EVAL_166;
  assign _EVAL_135 = _EVAL_202[4:0];
  assign _EVAL_242 = _EVAL_14 >= 2'h2;
  assign _EVAL_217 = _EVAL_243 & _EVAL_207;
  assign _EVAL_121 = _EVAL_215[4:0];
  assign _EVAL_156 = ~_EVAL_210;
  assign _EVAL_43 = _EVAL_144 | _EVAL_135;
  assign _EVAL_120 = _EVAL_236[0];
  assign _EVAL_139 = ~_EVAL_233;
  assign _EVAL_265 = _EVAL_234 | _EVAL_13;
  assign _EVAL_244 = _EVAL_131 | _EVAL_13;
  assign _EVAL_255 = _EVAL_43 & _EVAL_172;
  assign _EVAL_207 = _EVAL_0[1];
  assign _EVAL_53 = _EVAL_2 == 3'h0;
  assign _EVAL_203 = ~_EVAL_129;
  assign _EVAL_247 = _EVAL_12 <= 2'h2;
  assign _EVAL_45 = _EVAL_5 & _EVAL_100;
  assign _EVAL_112 = _EVAL_243 & _EVAL_252;
  assign _EVAL_19 = _EVAL_197[0];
  assign _EVAL_37 = _EVAL_171 | _EVAL_82;
  assign _EVAL_28 = ~_EVAL_99;
  assign _EVAL_127 = _EVAL_221 | _EVAL_13;
  assign _EVAL_158 = _EVAL_8 <= 2'h2;
  assign _EVAL_93 = {{28'd0}, _EVAL_261};
  assign _EVAL_22 = ~_EVAL_195;
  assign _EVAL_195 = _EVAL_3 == 3'h6;
  assign _EVAL_154 = _EVAL_6 <= 3'h4;
  assign _EVAL_181 = _EVAL_16 & _EVAL_141;
  assign _EVAL_76 = _EVAL_0[0];
  assign _EVAL_183 = _EVAL_104 & _EVAL_23;
  assign _EVAL_97 = _EVAL_135 != _EVAL_121;
  assign _EVAL_177 = _EVAL_171 | _EVAL_164;
  assign _EVAL_124 = ~_EVAL_271;
  assign _EVAL_174 = _EVAL_52[1:0];
  assign _EVAL_92 = _EVAL_1 & _EVAL_58;
  assign _EVAL_162 = _EVAL_41 | _EVAL_138;
  assign _EVAL_239 = _EVAL_2 == 3'h5;
  assign _EVAL_264 = _EVAL_2 == _EVAL_262;
  assign _EVAL_34 = ~_EVAL_159;
  assign _EVAL_64 = _EVAL_8 == _EVAL_191;
  assign _EVAL_240 = ~_EVAL_114;
  assign _EVAL_263 = _EVAL_102[0];
  assign _EVAL_136 = ~_EVAL_125;
  assign _EVAL_199 = _EVAL_9 == 3'h0;
  assign _EVAL_215 = _EVAL_130 ? _EVAL_187 : 8'h0;
  assign _EVAL_63 = _EVAL_179 | _EVAL_13;
  assign _EVAL_254 = _EVAL_16 & _EVAL_239;
  assign _EVAL_46 = _EVAL_268 | _EVAL_13;
  assign _EVAL_99 = _EVAL_96 | _EVAL_13;
  assign _EVAL_106 = _EVAL_16 & _EVAL_189;
  assign _EVAL_91 = _EVAL_2 == 3'h2;
  assign _EVAL_115 = _EVAL_65 | _EVAL_13;
  assign _EVAL_253 = _EVAL_5 & _EVAL_213;
  assign _EVAL_189 = _EVAL_2 == 3'h3;
  assign _EVAL_147 = _EVAL_184 | _EVAL_13;
  assign _EVAL_187 = 8'h1 << _EVAL_6;
  assign _EVAL_82 = _EVAL_42 & _EVAL_212;
  assign _EVAL_66 = plusarg_reader_out == 32'h0;
  assign _EVAL_196 = _EVAL_98 | _EVAL_7;
  assign _EVAL_60 = _EVAL_257 >> _EVAL_6;
  assign _EVAL_167 = _EVAL_133 | _EVAL_211;
  assign _EVAL_204 = _EVAL_142 - 1'h1;
  assign _EVAL_74 = _EVAL_144 >> _EVAL_4;
  assign _EVAL_108 = ~_EVAL_46;
  assign _EVAL_38 = _EVAL_238 & _EVAL_109;
  assign _EVAL_118 = ~_EVAL_224;
  assign _EVAL_251 = _EVAL_242 | _EVAL_13;
  assign _EVAL_67 = ~_EVAL_77;
  assign _EVAL_89 = _EVAL_252 & _EVAL_76;
  assign _EVAL_140 = ~_EVAL_209;
  assign _EVAL_109 = ~_EVAL_73;
  assign _EVAL_71 = ~_EVAL_36;
  assign _EVAL_230 = 8'h1 << _EVAL_4;
  assign _EVAL_98 = ~_EVAL_17;
  assign _EVAL_105 = _EVAL_17 == _EVAL_44;
  assign _EVAL_61 = _EVAL_5 & _EVAL_232;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_32 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_44 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_50 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_54 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_69 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_73 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_142 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_144 = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_152 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_153 = _RAND_9[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_155 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_165 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_170 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_191 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_233 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_249 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_262 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_15) begin
    if (_EVAL_39) begin
      _EVAL_32 <= _EVAL_9;
    end
    if (_EVAL_128) begin
      _EVAL_44 <= _EVAL_17;
    end
    if (_EVAL_39) begin
      _EVAL_50 <= _EVAL_4;
    end
    if (_EVAL_128) begin
      _EVAL_54 <= _EVAL_6;
    end
    if (_EVAL_128) begin
      _EVAL_69 <= _EVAL_3;
    end
    if (_EVAL_13) begin
      _EVAL_73 <= 1'h0;
    end else if (_EVAL_238) begin
      if (_EVAL_109) begin
        _EVAL_73 <= 1'h0;
      end else begin
        _EVAL_73 <= _EVAL_120;
      end
    end
    if (_EVAL_13) begin
      _EVAL_142 <= 1'h0;
    end else if (_EVAL_104) begin
      if (_EVAL_23) begin
        _EVAL_142 <= 1'h0;
      end else begin
        _EVAL_142 <= _EVAL_206;
      end
    end
    if (_EVAL_13) begin
      _EVAL_144 <= 5'h0;
    end else begin
      _EVAL_144 <= _EVAL_255;
    end
    if (_EVAL_13) begin
      _EVAL_152 <= 1'h0;
    end else if (_EVAL_104) begin
      if (_EVAL_95) begin
        _EVAL_152 <= 1'h0;
      end else begin
        _EVAL_152 <= _EVAL_263;
      end
    end
    if (_EVAL_39) begin
      _EVAL_153 <= _EVAL_0;
    end
    if (_EVAL_39) begin
      _EVAL_155 <= _EVAL_12;
    end
    if (_EVAL_13) begin
      _EVAL_165 <= 32'h0;
    end else if (_EVAL_225) begin
      _EVAL_165 <= 32'h0;
    end else begin
      _EVAL_165 <= _EVAL_103;
    end
    if (_EVAL_128) begin
      _EVAL_170 <= _EVAL_14;
    end
    if (_EVAL_128) begin
      _EVAL_191 <= _EVAL_8;
    end
    if (_EVAL_13) begin
      _EVAL_233 <= 1'h0;
    end else if (_EVAL_238) begin
      if (_EVAL_139) begin
        _EVAL_233 <= 1'h0;
      end else begin
        _EVAL_233 <= _EVAL_19;
      end
    end
    if (_EVAL_128) begin
      _EVAL_249 <= _EVAL_18;
    end
    if (_EVAL_39) begin
      _EVAL_262 <= _EVAL_2;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89b4180c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f353f76a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f17cc5da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56e66161)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37257089)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ffc0fa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41b51cd3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c3b3069)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d382ae4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4803a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15a43a06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2454b4cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8eb19de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b3ea07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0fa8014)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eac3de42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(980ece4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f43446b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37fabf26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20404cfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e26d7bff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3186991)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b27362a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98a4f20b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a77b44c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b838acb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afe9f6ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8376e8d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b5e0f08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd91bd60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5dee85a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cca589f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63d1c7fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(466b38ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d224afa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72e2a460)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ef9558)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6cd8631)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c4049c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e287356)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(488436d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d6726df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6abf053f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de3c2aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35322e59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec931edf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e15f098f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abd05652)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f84cdc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(483e7f00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(590d9e45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cb98bdb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(961ea605)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7f25708)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(312e8867)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14688790)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4bb78d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efd736bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c20bac25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a83f307)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a5c9f45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7778c9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6219529)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7a19f06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff52e9c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d05c9ce5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93b23275)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fc29ea2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d03546bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(195033b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f419768e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38160c67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd6da60f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18fef165)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66d6b6c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1050a5a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27e63d80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(241911d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cef39e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20fa6765)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d15adcd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fdd9336)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cb8af92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5599809)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45cf6de5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c93fa97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec52c56f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9be6ca0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81b526a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5b0cde8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3173ca34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1150393)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24c45af3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
