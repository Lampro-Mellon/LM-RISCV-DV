//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_94_assert(
  input         _EVAL,
  input  [1:0]  _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [1:0]  _EVAL_4,
  input         _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input  [1:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  input  [3:0]  _EVAL_11,
  input         _EVAL_12,
  input  [29:0] _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18
);
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire [31:0] _EVAL_22;
  reg  _EVAL_23;
  reg [31:0] _RAND_0;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire [3:0] _EVAL_28;
  reg [31:0] _EVAL_29;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_30;
  reg [31:0] _RAND_2;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire [4:0] _EVAL_47;
  wire [32:0] _EVAL_48;
  wire [4:0] _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire [1:0] _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire [7:0] _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  reg [4:0] _EVAL_77;
  reg [31:0] _RAND_3;
  wire [30:0] _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire [7:0] _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire [3:0] _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire [4:0] _EVAL_95;
  wire [1:0] _EVAL_96;
  reg  _EVAL_97;
  reg [31:0] _RAND_4;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire [1:0] _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_104;
  wire [30:0] _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire [4:0] _EVAL_115;
  reg  _EVAL_116;
  reg [31:0] _RAND_5;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire [3:0] _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire [1:0] _EVAL_122;
  wire  _EVAL_123;
  wire [1:0] _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  reg  _EVAL_130;
  reg [31:0] _RAND_6;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [4:0] _EVAL_143;
  reg  _EVAL_144;
  reg [31:0] _RAND_7;
  wire  _EVAL_145;
  wire  _EVAL_146;
  reg [1:0] _EVAL_147;
  reg [31:0] _RAND_8;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  reg [1:0] _EVAL_155;
  reg [31:0] _RAND_9;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  reg  _EVAL_161;
  reg [31:0] _RAND_10;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire [29:0] _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire [1:0] _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire [7:0] _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  reg [2:0] _EVAL_183;
  reg [31:0] _RAND_11;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  reg [29:0] _EVAL_189;
  reg [31:0] _RAND_12;
  wire  _EVAL_190;
  wire [29:0] _EVAL_191;
  wire [3:0] _EVAL_192;
  wire [30:0] _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  reg [2:0] _EVAL_197;
  reg [31:0] _RAND_13;
  wire [4:0] _EVAL_198;
  wire  _EVAL_199;
  wire [1:0] _EVAL_200;
  reg [2:0] _EVAL_201;
  reg [31:0] _RAND_14;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire [4:0] _EVAL_205;
  wire  _EVAL_206;
  wire [1:0] _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  reg [1:0] _EVAL_227;
  reg [31:0] _RAND_15;
  wire [7:0] _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire [4:0] _EVAL_233;
  wire [29:0] _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire [1:0] _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire [4:0] _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire [1:0] _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  reg [2:0] _EVAL_279;
  reg [31:0] _RAND_16;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_37 = _EVAL_16 & _EVAL_117;
  assign _EVAL_131 = _EVAL_276 & _EVAL_27;
  assign _EVAL_31 = ~_EVAL_252;
  assign _EVAL_47 = _EVAL_205 | _EVAL_77;
  assign _EVAL_149 = _EVAL_9 <= 3'h4;
  assign _EVAL_61 = ~_EVAL_97;
  assign _EVAL_74 = ~_EVAL_107;
  assign _EVAL_244 = _EVAL_11 == _EVAL_28;
  assign _EVAL_33 = _EVAL_150 | _EVAL_217;
  assign _EVAL_145 = ~_EVAL_237;
  assign _EVAL_191 = {{28'd0}, _EVAL_54};
  assign _EVAL_92 = ~_EVAL_11;
  assign _EVAL_213 = _EVAL_38 | _EVAL_5;
  assign _EVAL_174 = _EVAL_13 == _EVAL_189;
  assign _EVAL_199 = _EVAL_49[0];
  assign _EVAL_236 = _EVAL_217 & _EVAL_126;
  assign _EVAL_224 = _EVAL_243 | _EVAL_5;
  assign _EVAL_151 = _EVAL_245 | _EVAL_5;
  assign _EVAL_165 = ~_EVAL_86;
  assign _EVAL_233 = _EVAL_246 & _EVAL_198;
  assign _EVAL_157 = _EVAL_2 == 3'h4;
  assign _EVAL_228 = _EVAL_283 ? _EVAL_89 : 8'h0;
  assign _EVAL_113 = _EVAL_18 == _EVAL_23;
  assign _EVAL_282 = _EVAL_16 & _EVAL_50;
  assign _EVAL_180 = _EVAL_150 & _EVAL_61;
  assign _EVAL_248 = _EVAL_1 <= 3'h6;
  assign _EVAL_121 = ~_EVAL_152;
  assign _EVAL_79 = _EVAL_29 < plusarg_reader_out;
  assign _EVAL_88 = _EVAL_120 | _EVAL_5;
  assign _EVAL_122 = _EVAL_170 | 2'h1;
  assign _EVAL_65 = _EVAL_3 == 3'h7;
  assign _EVAL_271 = _EVAL_2[2:1];
  assign _EVAL_273 = _EVAL_256 | _EVAL_118;
  assign _EVAL_62 = _EVAL_110 | _EVAL_5;
  assign _EVAL_156 = _EVAL_122[0];
  assign _EVAL_246 = _EVAL_77 | _EVAL_205;
  assign _EVAL_83 = _EVAL_3 == _EVAL_183;
  assign _EVAL_163 = ~_EVAL_17;
  assign _EVAL_190 = ~_EVAL_194;
  assign _EVAL_207 = _EVAL_130 - 1'h1;
  assign _EVAL_238 = ~_EVAL_5;
  assign _EVAL_53 = _EVAL_137 | _EVAL_278;
  assign _EVAL_219 = _EVAL_4 == _EVAL_147;
  assign _EVAL_195 = ~_EVAL_166;
  assign _EVAL_91 = _EVAL_9 == 3'h0;
  assign _EVAL_54 = ~_EVAL_242;
  assign _EVAL_105 = _EVAL_193;
  assign _EVAL_208 = _EVAL_4 == 2'h0;
  assign _EVAL_285 = _EVAL_96 == 2'h1;
  assign _EVAL_125 = ~_EVAL_266;
  assign _EVAL_112 = ~_EVAL_116;
  assign _EVAL_200 = _EVAL_116 - 1'h1;
  assign _EVAL_178 = _EVAL_223 | _EVAL_5;
  assign _EVAL_119 = ~_EVAL_28;
  assign _EVAL_34 = ~_EVAL_230;
  assign _EVAL_226 = ~_EVAL_130;
  assign _EVAL_66 = _EVAL_200[0];
  assign _EVAL_179 = _EVAL_51 | _EVAL_5;
  assign _EVAL_221 = ~_EVAL_153;
  assign _EVAL_284 = ~_EVAL_67;
  assign _EVAL_241 = ~_EVAL_169;
  assign _EVAL_60 = ~_EVAL_226;
  assign _EVAL_154 = ~_EVAL_178;
  assign _EVAL_283 = _EVAL_150 & _EVAL_112;
  assign _EVAL_258 = _EVAL_12 & _EVAL_265;
  assign _EVAL_25 = ~_EVAL_44;
  assign _EVAL_252 = _EVAL_254 | _EVAL_5;
  assign _EVAL_142 = _EVAL_12 & _EVAL_138;
  assign _EVAL_108 = _EVAL_16 & _EVAL_76;
  assign _EVAL_22 = _EVAL_48[31:0];
  assign _EVAL_20 = _EVAL_6 == 3'h4;
  assign _EVAL_206 = _EVAL_12 & _EVAL_109;
  assign _EVAL_93 = _EVAL_199 | _EVAL_5;
  assign _EVAL_64 = _EVAL_156 & _EVAL_267;
  assign _EVAL_150 = _EVAL_7 & _EVAL_16;
  assign _EVAL_32 = _EVAL_2 == _EVAL_279;
  assign _EVAL_216 = _EVAL_16 & _EVAL_75;
  assign _EVAL_58 = _EVAL_156 & _EVAL_225;
  assign _EVAL_260 = _EVAL_205 != _EVAL_115;
  assign _EVAL_36 = _EVAL_4 <= 2'h2;
  assign _EVAL_242 = _EVAL_95[1:0];
  assign _EVAL_235 = _EVAL_122[1];
  assign _EVAL_264 = _EVAL_208 | _EVAL_5;
  assign _EVAL_172 = _EVAL_16 & _EVAL_261;
  assign _EVAL_43 = _EVAL_271 == 2'h1;
  assign _EVAL_276 = ~_EVAL_90;
  assign _EVAL_115 = _EVAL_175[4:0];
  assign _EVAL_275 = ~_EVAL_136;
  assign _EVAL_234 = _EVAL_13 ^ 30'h20000000;
  assign _EVAL_272 = ~_EVAL_82;
  assign _EVAL_98 = ~_EVAL_104;
  assign _EVAL_114 = _EVAL_174 | _EVAL_5;
  assign _EVAL_202 = ~_EVAL_159;
  assign _EVAL_27 = ~_EVAL_204;
  assign _EVAL_251 = _EVAL_271 == 2'h0;
  assign _EVAL_87 = _EVAL_1 == 3'h0;
  assign _EVAL_277 = ~_EVAL_264;
  assign _EVAL_49 = _EVAL_47 >> _EVAL_6;
  assign _EVAL_265 = _EVAL_1 == 3'h1;
  assign _EVAL_170 = 2'h1 << _EVAL_176;
  assign _EVAL_173 = _EVAL_276 & _EVAL_204;
  assign _EVAL_256 = ~_EVAL_146;
  assign _EVAL_245 = _EVAL_9 <= 3'h2;
  assign _EVAL_46 = _EVAL_231 | _EVAL_5;
  assign _EVAL_89 = 8'h1 << _EVAL_2;
  assign _EVAL_218 = ~_EVAL_140;
  assign _EVAL_72 = _EVAL_12 & _EVAL_60;
  assign _EVAL_193 = $signed(_EVAL_78) & -31'sh2000;
  assign _EVAL_243 = _EVAL_274 | _EVAL_20;
  assign _EVAL_21 = _EVAL_73 | _EVAL_5;
  assign _EVAL_141 = _EVAL_120 | _EVAL_17;
  assign _EVAL_100 = _EVAL_235 & _EVAL_90;
  assign _EVAL_160 = _EVAL_262 | _EVAL_5;
  assign _EVAL_169 = _EVAL_171 | _EVAL_5;
  assign _EVAL_198 = ~_EVAL_115;
  assign _EVAL_203 = ~_EVAL_45;
  assign _EVAL_168 = _EVAL_255 | _EVAL_5;
  assign _EVAL_128 = _EVAL_68 | _EVAL_5;
  assign _EVAL_280 = _EVAL_124[0];
  assign _EVAL_90 = _EVAL_13[1];
  assign _EVAL_164 = _EVAL_13 & _EVAL_191;
  assign _EVAL_262 = _EVAL_260 | _EVAL_247;
  assign _EVAL_109 = _EVAL_1 == 3'h5;
  assign _EVAL_124 = _EVAL_97 - 1'h1;
  assign _EVAL_44 = _EVAL_143[0];
  assign _EVAL_205 = _EVAL_228[4:0];
  assign _EVAL_158 = ~_EVAL_128;
  assign _EVAL_215 = _EVAL_1 == 3'h4;
  assign _EVAL_278 = _EVAL_156 & _EVAL_173;
  assign _EVAL_143 = _EVAL_77 >> _EVAL_2;
  assign _EVAL_86 = _EVAL_269 | _EVAL_5;
  assign _EVAL_99 = ~_EVAL_213;
  assign _EVAL_232 = _EVAL_156 & _EVAL_131;
  assign _EVAL_94 = _EVAL_273 | _EVAL_79;
  assign _EVAL_222 = _EVAL_236 & _EVAL_39;
  assign _EVAL_140 = _EVAL_113 | _EVAL_5;
  assign _EVAL_45 = _EVAL_248 | _EVAL_5;
  assign _EVAL_107 = _EVAL_36 | _EVAL_5;
  assign _EVAL_78 = {1'b0,$signed(_EVAL_234)};
  assign _EVAL_73 = _EVAL_10 == _EVAL_144;
  assign _EVAL_253 = _EVAL_235 & _EVAL_276;
  assign _EVAL_41 = ~_EVAL_93;
  assign _EVAL_132 = _EVAL_16 & _EVAL_123;
  assign _EVAL_42 = ~_EVAL_148;
  assign _EVAL_188 = ~_EVAL_184;
  assign _EVAL_138 = _EVAL_1 == 3'h2;
  assign _EVAL_57 = 8'h1 << _EVAL_6;
  assign _EVAL_40 = ~_EVAL_179;
  assign _EVAL_240 = ~_EVAL_21;
  assign _EVAL_211 = _EVAL_43 | _EVAL_251;
  assign _EVAL_101 = _EVAL_161 - 1'h1;
  assign _EVAL_50 = _EVAL_3 == 3'h1;
  assign _EVAL_247 = ~_EVAL_268;
  assign _EVAL_159 = _EVAL_94 | _EVAL_5;
  assign _EVAL_69 = ~_EVAL_62;
  assign _EVAL_24 = _EVAL_0 >= 2'h2;
  assign _EVAL_70 = _EVAL_214 | _EVAL_100;
  assign _EVAL_126 = ~_EVAL_161;
  assign _EVAL_210 = _EVAL_52 | _EVAL_5;
  assign _EVAL_118 = plusarg_reader_out == 32'h0;
  assign _EVAL_177 = _EVAL_16 & _EVAL_65;
  assign _EVAL_259 = _EVAL_9 <= 3'h1;
  assign _EVAL_59 = _EVAL_8 <= 2'h2;
  assign _EVAL_214 = _EVAL_8 >= 2'h2;
  assign _EVAL_135 = ~_EVAL_151;
  assign _EVAL_184 = _EVAL_149 | _EVAL_5;
  assign _EVAL_223 = _EVAL_9 == _EVAL_30;
  assign _EVAL_81 = ~_EVAL_26;
  assign _EVAL_120 = ~_EVAL_10;
  assign _EVAL_281 = _EVAL_91 | _EVAL_5;
  assign _EVAL_102 = ~_EVAL_224;
  assign _EVAL_237 = _EVAL_32 | _EVAL_5;
  assign _EVAL_85 = _EVAL_217 & _EVAL_226;
  assign _EVAL_96 = _EVAL_6[2:1];
  assign _EVAL_192 = _EVAL_11 & _EVAL_119;
  assign _EVAL_196 = _EVAL_164 == 30'h0;
  assign _EVAL_167 = ~_EVAL_168;
  assign _EVAL_230 = _EVAL_24 | _EVAL_5;
  assign _EVAL_229 = _EVAL_96 == 2'h0;
  assign _EVAL_136 = _EVAL_141 | _EVAL_5;
  assign _EVAL_127 = ~_EVAL_281;
  assign _EVAL_56 = _EVAL_101[0];
  assign _EVAL_176 = _EVAL_8[0];
  assign _EVAL_171 = ~_EVAL_14;
  assign _EVAL_220 = _EVAL_16 & _EVAL_187;
  assign _EVAL_266 = _EVAL_163 | _EVAL_5;
  assign _EVAL_182 = $signed(_EVAL_105) == 31'sh0;
  assign _EVAL_123 = _EVAL_3 == 3'h2;
  assign _EVAL_269 = _EVAL_92 == 4'h0;
  assign _EVAL_133 = _EVAL_207[0];
  assign _EVAL_80 = _EVAL_137 | _EVAL_232;
  assign _EVAL_186 = _EVAL_12 & _EVAL_87;
  assign _EVAL_75 = _EVAL_3 == 3'h6;
  assign _EVAL_254 = _EVAL_1 == _EVAL_197;
  assign _EVAL_137 = _EVAL_214 | _EVAL_253;
  assign _EVAL_194 = _EVAL_25 | _EVAL_5;
  assign _EVAL_134 = ~_EVAL_210;
  assign _EVAL_129 = _EVAL_70 | _EVAL_58;
  assign _EVAL_162 = _EVAL_12 & _EVAL_215;
  assign _EVAL_26 = _EVAL_219 | _EVAL_5;
  assign _EVAL_153 = _EVAL_111 | _EVAL_5;
  assign _EVAL_52 = _EVAL_9 <= 3'h3;
  assign _EVAL_48 = _EVAL_29 + 32'h1;
  assign _EVAL_110 = _EVAL_6 == _EVAL_201;
  assign _EVAL_204 = _EVAL_13[0];
  assign _EVAL_166 = _EVAL_214 | _EVAL_5;
  assign _EVAL_231 = _EVAL_192 == 4'h0;
  assign _EVAL_39 = ~_EVAL_270;
  assign _EVAL_225 = _EVAL_90 & _EVAL_204;
  assign _EVAL_68 = _EVAL_8 == _EVAL_227;
  assign _EVAL_261 = _EVAL_3 == 3'h5;
  assign _EVAL_175 = _EVAL_222 ? _EVAL_57 : 8'h0;
  assign _EVAL_217 = _EVAL & _EVAL_12;
  assign _EVAL_255 = _EVAL_0 == _EVAL_155;
  assign _EVAL_257 = _EVAL_12 & _EVAL_270;
  assign _EVAL_146 = _EVAL_77 != 5'h0;
  assign _EVAL_267 = _EVAL_90 & _EVAL_27;
  assign _EVAL_274 = _EVAL_285 | _EVAL_229;
  assign _EVAL_104 = _EVAL_196 | _EVAL_5;
  assign _EVAL_181 = ~_EVAL_160;
  assign _EVAL_38 = _EVAL_59 & _EVAL_182;
  assign _EVAL_51 = _EVAL_211 | _EVAL_157;
  assign _EVAL_35 = ~_EVAL_88;
  assign _EVAL_185 = _EVAL_9 != 3'h0;
  assign _EVAL_111 = _EVAL_4 != 2'h2;
  assign _EVAL_268 = _EVAL_205 != 5'h0;
  assign _EVAL_187 = _EVAL_3 == 3'h0;
  assign _EVAL_55 = _EVAL_16 & _EVAL_106;
  assign _EVAL_249 = ~_EVAL_114;
  assign _EVAL_95 = 5'h3 << _EVAL_8;
  assign _EVAL_106 = _EVAL_3 == 3'h4;
  assign _EVAL_67 = _EVAL_83 | _EVAL_5;
  assign _EVAL_28 = {_EVAL_129,_EVAL_250,_EVAL_53,_EVAL_80};
  assign _EVAL_270 = _EVAL_1 == 3'h6;
  assign _EVAL_82 = _EVAL_259 | _EVAL_5;
  assign _EVAL_250 = _EVAL_70 | _EVAL_64;
  assign _EVAL_63 = ~_EVAL_46;
  assign _EVAL_152 = _EVAL_244 | _EVAL_5;
  assign _EVAL_76 = _EVAL_3 == 3'h3;
  assign _EVAL_148 = _EVAL_185 | _EVAL_5;
  assign _EVAL_117 = ~_EVAL_61;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_29 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_30 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_77 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_97 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_116 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_130 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_144 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_147 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_155 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_161 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_183 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_189 = _RAND_12[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_197 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_201 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_227 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_279 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_15) begin
    if (_EVAL_85) begin
      _EVAL_23 <= _EVAL_18;
    end
    if (_EVAL_5) begin
      _EVAL_29 <= 32'h0;
    end else if (_EVAL_33) begin
      _EVAL_29 <= 32'h0;
    end else begin
      _EVAL_29 <= _EVAL_22;
    end
    if (_EVAL_180) begin
      _EVAL_30 <= _EVAL_9;
    end
    if (_EVAL_5) begin
      _EVAL_77 <= 5'h0;
    end else begin
      _EVAL_77 <= _EVAL_233;
    end
    if (_EVAL_5) begin
      _EVAL_97 <= 1'h0;
    end else if (_EVAL_150) begin
      if (_EVAL_61) begin
        _EVAL_97 <= 1'h0;
      end else begin
        _EVAL_97 <= _EVAL_280;
      end
    end
    if (_EVAL_5) begin
      _EVAL_116 <= 1'h0;
    end else if (_EVAL_150) begin
      if (_EVAL_112) begin
        _EVAL_116 <= 1'h0;
      end else begin
        _EVAL_116 <= _EVAL_66;
      end
    end
    if (_EVAL_5) begin
      _EVAL_130 <= 1'h0;
    end else if (_EVAL_217) begin
      if (_EVAL_226) begin
        _EVAL_130 <= 1'h0;
      end else begin
        _EVAL_130 <= _EVAL_133;
      end
    end
    if (_EVAL_85) begin
      _EVAL_144 <= _EVAL_10;
    end
    if (_EVAL_85) begin
      _EVAL_147 <= _EVAL_4;
    end
    if (_EVAL_85) begin
      _EVAL_155 <= _EVAL_0;
    end
    if (_EVAL_5) begin
      _EVAL_161 <= 1'h0;
    end else if (_EVAL_217) begin
      if (_EVAL_126) begin
        _EVAL_161 <= 1'h0;
      end else begin
        _EVAL_161 <= _EVAL_56;
      end
    end
    if (_EVAL_180) begin
      _EVAL_183 <= _EVAL_3;
    end
    if (_EVAL_180) begin
      _EVAL_189 <= _EVAL_13;
    end
    if (_EVAL_85) begin
      _EVAL_197 <= _EVAL_1;
    end
    if (_EVAL_85) begin
      _EVAL_201 <= _EVAL_6;
    end
    if (_EVAL_180) begin
      _EVAL_227 <= _EVAL_8;
    end
    if (_EVAL_180) begin
      _EVAL_279 <= _EVAL_2;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a219997d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d86af58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1d5f1a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(590bb7d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ed2fe4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5da18dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3490b4cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5946042)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(affc04c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2403d296)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_275) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5aae083d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f1e19cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68c4cb41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89967b03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5438e4c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8f7d3b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19821de5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4636123)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ec0dfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_275) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(888f78f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fafae22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e90a2d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfd182b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(843195cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(914787fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b678d6cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b587bf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ae2289c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bfb7ba4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6f5b029)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64d4e109)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(718f49b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18934298)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9699482e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11c42c7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_275) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(258b1158)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38025dae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9f85e8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c381a7ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a2f2223)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7dc98393)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af548851)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_31) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5dd58177)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(150a644a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85dd8d47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d7381ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_275) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abba8d6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f84e455d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4d2bb3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1356846a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5efab74c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a5edf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b779dd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_284) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3da1149)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39b5627b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b9b066e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dec3c92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe37cd3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56696367)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5244e582)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1f9d6d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bb9c118)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_31) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed3a95ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acc598bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c92c8c4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a1c53ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d99851b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(496acfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15185c62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5f76373)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4367091a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da660764)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89ebfc64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e392ce7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45e0894)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6603b2fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_284) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(728d8a14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d614e5d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10f8eb3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(659c7995)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bffcb25d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(838057cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9ff4cc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(496c40de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50ae2cbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dad53424)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bec8c2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(affd3034)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1d26a0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68a92bf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9407c91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7383f7fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69acf6a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
