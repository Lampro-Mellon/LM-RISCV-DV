//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_23_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [1:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [30:0] _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input  [3:0]  _EVAL_15,
  input  [2:0]  _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18
);
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire [5:0] _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  reg [2:0] _EVAL_28;
  reg [31:0] _RAND_0;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire [4:0] _EVAL_33;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire [5:0] _EVAL_37;
  wire  _EVAL_38;
  wire [1:0] _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_48;
  wire [5:0] _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire [1:0] _EVAL_52;
  wire  _EVAL_53;
  reg [4:0] _EVAL_54;
  reg [31:0] _RAND_1;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire [12:0] _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire [12:0] _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire [31:0] _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_76;
  wire [3:0] _EVAL_77;
  wire [3:0] _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire [31:0] _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire [4:0] _EVAL_92;
  wire [4:0] _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire [4:0] _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  reg [2:0] _EVAL_105;
  reg [31:0] _RAND_2;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire [30:0] _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire [3:0] _EVAL_122;
  wire [30:0] _EVAL_123;
  reg [2:0] _EVAL_124;
  reg [31:0] _RAND_3;
  wire  _EVAL_125;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire [3:0] _EVAL_129;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_131;
  wire  _EVAL_132;
  reg [2:0] _EVAL_133;
  reg [31:0] _RAND_4;
  wire  _EVAL_134;
  reg [2:0] _EVAL_135;
  reg [31:0] _RAND_5;
  wire [4:0] _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire [4:0] _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  reg  _EVAL_144;
  reg [31:0] _RAND_6;
  wire  _EVAL_145;
  reg [3:0] _EVAL_146;
  reg [31:0] _RAND_7;
  wire  _EVAL_147;
  wire [7:0] _EVAL_148;
  wire  _EVAL_149;
  wire [3:0] _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire [4:0] _EVAL_158;
  wire [4:0] _EVAL_159;
  wire  _EVAL_160;
  reg [31:0] _EVAL_161;
  reg [31:0] _RAND_8;
  wire  _EVAL_162;
  wire [31:0] _EVAL_163;
  wire  _EVAL_164;
  wire [3:0] _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire [3:0] _EVAL_170;
  wire  _EVAL_171;
  wire [4:0] _EVAL_172;
  wire  _EVAL_173;
  wire [7:0] _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire [5:0] _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire [4:0] _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire [31:0] _EVAL_199;
  wire  _EVAL_200;
  wire [7:0] _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  reg [3:0] _EVAL_211;
  reg [31:0] _RAND_9;
  wire [3:0] _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  reg [30:0] _EVAL_215;
  reg [31:0] _RAND_10;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  reg [2:0] _EVAL_224;
  reg [31:0] _RAND_11;
  wire [4:0] _EVAL_225;
  wire  _EVAL_227;
  wire  _EVAL_228;
  reg [3:0] _EVAL_229;
  reg [31:0] _RAND_12;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire [7:0] _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire [1:0] _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire [1:0] _EVAL_249;
  wire  _EVAL_250;
  wire [4:0] _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  reg [1:0] _EVAL_260;
  reg [31:0] _RAND_13;
  wire [30:0] _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire [3:0] _EVAL_270;
  wire  _EVAL_271;
  reg  _EVAL_272;
  reg [31:0] _RAND_14;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire [32:0] _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire [3:0] _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  reg [2:0] _EVAL_291;
  reg [31:0] _RAND_15;
  reg [3:0] _EVAL_292;
  reg [31:0] _RAND_16;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_171 = _EVAL_236 & _EVAL_69;
  assign _EVAL_280 = _EVAL_191 | _EVAL_8;
  assign _EVAL_222 = _EVAL_244 == 2'h0;
  assign _EVAL_116 = ~_EVAL_180;
  assign _EVAL_219 = ~_EVAL_70;
  assign _EVAL_281 = _EVAL_12 <= 3'h3;
  assign _EVAL_253 = _EVAL_0 == _EVAL_28;
  assign _EVAL_290 = _EVAL_14 & _EVAL_32;
  assign _EVAL_207 = _EVAL_12 <= 3'h2;
  assign _EVAL_42 = _EVAL_76 & _EVAL_258;
  assign _EVAL_63 = ~_EVAL_153;
  assign _EVAL_230 = _EVAL_137 | _EVAL_8;
  assign _EVAL_108 = _EVAL_253 | _EVAL_8;
  assign _EVAL_284 = _EVAL_15 & _EVAL_122;
  assign _EVAL_85 = _EVAL_9 & _EVAL_14;
  assign _EVAL_134 = _EVAL_12 != 3'h0;
  assign _EVAL_196 = _EVAL_1 == 3'h0;
  assign _EVAL_181 = _EVAL_1 == 3'h5;
  assign _EVAL_131 = _EVAL_106 | _EVAL_8;
  assign _EVAL_237 = ~_EVAL_5;
  assign _EVAL_39 = _EVAL_16[2:1];
  assign _EVAL_19 = _EVAL_236 & _EVAL_71;
  assign _EVAL_78 = _EVAL_93[3:0];
  assign _EVAL_30 = _EVAL_15 == _EVAL_212;
  assign _EVAL_113 = _EVAL_12 == _EVAL_224;
  assign _EVAL_264 = _EVAL_237 | _EVAL;
  assign _EVAL_118 = _EVAL_48 | _EVAL_8;
  assign _EVAL_156 = ~_EVAL_97;
  assign _EVAL_59 = ~_EVAL_206;
  assign _EVAL_227 = _EVAL_2 == 2'h0;
  assign _EVAL_238 = _EVAL_85 & _EVAL_79;
  assign _EVAL_141 = _EVAL_6 & _EVAL_125;
  assign _EVAL_267 = ~_EVAL_72;
  assign _EVAL_185 = _EVAL_7 == _EVAL_215;
  assign _EVAL_21 = _EVAL_61[5:0];
  assign _EVAL_162 = _EVAL_7[1];
  assign _EVAL_149 = _EVAL_4 == _EVAL_124;
  assign _EVAL_86 = _EVAL_0 >= 3'h2;
  assign _EVAL_294 = _EVAL_0 <= 3'h6;
  assign _EVAL_73 = $signed(_EVAL_199) & -32'sh2000;
  assign _EVAL_177 = _EVAL_292 == 4'h0;
  assign _EVAL_293 = _EVAL_92[0];
  assign _EVAL_48 = _EVAL_5 == _EVAL_144;
  assign _EVAL_112 = _EVAL_16 == 3'h4;
  assign _EVAL_132 = _EVAL_295 | _EVAL_8;
  assign _EVAL_236 = _EVAL_52[0];
  assign _EVAL_50 = ~_EVAL_68;
  assign _EVAL_254 = _EVAL_39 == 2'h1;
  assign _EVAL_129 = _EVAL_195[3:0];
  assign _EVAL_107 = ~_EVAL_205;
  assign _EVAL_255 = ~_EVAL_132;
  assign _EVAL_178 = _EVAL_53 | _EVAL_8;
  assign _EVAL_125 = _EVAL_1 == 3'h2;
  assign _EVAL_102 = _EVAL_52[1];
  assign _EVAL_183 = _EVAL_1 == 3'h1;
  assign _EVAL_200 = _EVAL_56 | _EVAL_8;
  assign _EVAL_288 = _EVAL_86 | _EVAL_216;
  assign _EVAL_175 = ~_EVAL_8;
  assign _EVAL_70 = _EVAL_66 | _EVAL_8;
  assign _EVAL_221 = _EVAL_257 | _EVAL_8;
  assign _EVAL_208 = _EVAL_3 == 3'h4;
  assign _EVAL_169 = ~_EVAL_230;
  assign _EVAL_246 = ~_EVAL_74;
  assign _EVAL_186 = _EVAL_6 & _EVAL_181;
  assign _EVAL_287 = _EVAL_256 | _EVAL_8;
  assign _EVAL_258 = _EVAL_211 == 4'h0;
  assign _EVAL_217 = _EVAL_185 | _EVAL_8;
  assign _EVAL_68 = _EVAL_1 == 3'h6;
  assign _EVAL_235 = _EVAL_3 == 3'h1;
  assign _EVAL_275 = _EVAL_3 == 3'h5;
  assign _EVAL_286 = _EVAL_14 & _EVAL_275;
  assign _EVAL_69 = _EVAL_162 & _EVAL_59;
  assign _EVAL_182 = _EVAL_264 | _EVAL_8;
  assign _EVAL_256 = _EVAL_2 == _EVAL_260;
  assign _EVAL_206 = _EVAL_7[0];
  assign _EVAL_101 = _EVAL_155 | _EVAL_8;
  assign _EVAL_120 = _EVAL_3 == 3'h2;
  assign _EVAL_283 = _EVAL_121 | _EVAL_8;
  assign _EVAL_277 = _EVAL_85 & _EVAL_177;
  assign _EVAL_153 = _EVAL_149 | _EVAL_8;
  assign _EVAL_249 = 2'h1 << _EVAL_147;
  assign _EVAL_81 = _EVAL_162 & _EVAL_206;
  assign _EVAL_61 = 13'h3f << _EVAL_0;
  assign _EVAL_184 = _EVAL_17 == _EVAL_272;
  assign _EVAL_104 = _EVAL_3[2];
  assign _EVAL_142 = _EVAL_1 <= 3'h6;
  assign _EVAL_38 = _EVAL_225 != _EVAL_99;
  assign _EVAL_55 = ~_EVAL_209;
  assign _EVAL_210 = plusarg_reader_out == 32'h0;
  assign _EVAL_167 = ~_EVAL_96;
  assign _EVAL_232 = ~_EVAL_80;
  assign _EVAL_119 = $signed(_EVAL_163) == 32'sh0;
  assign _EVAL_79 = _EVAL_146 == 4'h0;
  assign _EVAL_170 = _EVAL_37[5:2];
  assign _EVAL_137 = ~_EVAL_18;
  assign _EVAL_35 = ~_EVAL_109;
  assign _EVAL_31 = _EVAL_42 & _EVAL_50;
  assign _EVAL_192 = ~_EVAL_21;
  assign _EVAL_121 = _EVAL_16 == _EVAL_135;
  assign _EVAL_76 = _EVAL_13 & _EVAL_6;
  assign _EVAL_53 = _EVAL_94 | _EVAL_259;
  assign _EVAL_122 = ~_EVAL_212;
  assign _EVAL_201 = _EVAL_238 ? _EVAL_148 : 8'h0;
  assign _EVAL_268 = _EVAL_236 & _EVAL_285;
  assign _EVAL_214 = _EVAL_254 | _EVAL_282;
  assign _EVAL_123 = _EVAL_7 ^ 31'h40000000;
  assign _EVAL_174 = 8'h1 << _EVAL_16;
  assign _EVAL_228 = _EVAL_214 | _EVAL_112;
  assign _EVAL_44 = _EVAL_134 | _EVAL_8;
  assign _EVAL_49 = _EVAL_57[5:0];
  assign _EVAL_33 = _EVAL_159 & _EVAL_172;
  assign _EVAL_244 = _EVAL_4[2:1];
  assign _EVAL_58 = _EVAL_2 != 2'h2;
  assign _EVAL_191 = ~_EVAL_293;
  assign _EVAL_88 = _EVAL_6 & _EVAL_68;
  assign _EVAL_43 = _EVAL_6 & _EVAL_183;
  assign _EVAL_289 = ~_EVAL_287;
  assign _EVAL_278 = _EVAL_4 == 3'h4;
  assign _EVAL_51 = _EVAL_229 == 4'h0;
  assign _EVAL_245 = ~_EVAL_84;
  assign _EVAL_98 = ~_EVAL_91;
  assign _EVAL_25 = _EVAL_102 & _EVAL_36;
  assign _EVAL_56 = _EVAL_2 <= 2'h2;
  assign _EVAL_193 = ~_EVAL_108;
  assign _EVAL_180 = _EVAL_90 | _EVAL_8;
  assign _EVAL_143 = _EVAL_14 & _EVAL_114;
  assign _EVAL_168 = ~_EVAL_177;
  assign _EVAL_204 = ~_EVAL_51;
  assign _EVAL_173 = _EVAL_86 | _EVAL_25;
  assign _EVAL_248 = _EVAL_225 != 5'h0;
  assign _EVAL_195 = _EVAL_229 - 4'h1;
  assign _EVAL_60 = ~_EVAL_104;
  assign _EVAL_251 = _EVAL_211 - 4'h1;
  assign _EVAL_242 = ~_EVAL_217;
  assign _EVAL_80 = _EVAL_228 | _EVAL_8;
  assign _EVAL_209 = _EVAL_54 != 5'h0;
  assign _EVAL_259 = _EVAL_161 < plusarg_reader_out;
  assign _EVAL_285 = _EVAL_36 & _EVAL_206;
  assign _EVAL_197 = ~_EVAL_118;
  assign _EVAL_295 = _EVAL_1 == _EVAL_133;
  assign _EVAL_198 = _EVAL_76 & _EVAL_51;
  assign _EVAL_250 = _EVAL_14 & _EVAL_67;
  assign _EVAL_82 = _EVAL_213 | _EVAL_8;
  assign _EVAL_32 = _EVAL_3 == 3'h3;
  assign _EVAL_52 = _EVAL_249 | 2'h1;
  assign _EVAL_270 = _EVAL_192[5:2];
  assign _EVAL_67 = _EVAL_3 == 3'h6;
  assign _EVAL_22 = _EVAL_30 | _EVAL_8;
  assign _EVAL_166 = _EVAL_284 == 4'h0;
  assign _EVAL_24 = _EVAL_288 | _EVAL_171;
  assign _EVAL_100 = ~_EVAL_103;
  assign _EVAL_27 = _EVAL_1 == 3'h4;
  assign _EVAL_151 = ~_EVAL_127;
  assign _EVAL_265 = _EVAL_288 | _EVAL_29;
  assign _EVAL_66 = _EVAL_12 == 3'h0;
  assign _EVAL_92 = _EVAL_54 >> _EVAL_4;
  assign _EVAL_220 = ~_EVAL;
  assign _EVAL_205 = _EVAL_271 | _EVAL_8;
  assign _EVAL_91 = _EVAL_58 | _EVAL_8;
  assign _EVAL_233 = _EVAL_14 & _EVAL_154;
  assign _EVAL_243 = _EVAL_1[0];
  assign _EVAL_83 = _EVAL_276[31:0];
  assign _EVAL_94 = _EVAL_55 | _EVAL_210;
  assign _EVAL_194 = _EVAL_14 & _EVAL_208;
  assign _EVAL_89 = _EVAL_261 == 31'h0;
  assign _EVAL_158 = _EVAL_146 - 4'h1;
  assign _EVAL_72 = _EVAL_207 | _EVAL_8;
  assign _EVAL_179 = ~_EVAL_164;
  assign _EVAL_276 = _EVAL_161 + 32'h1;
  assign _EVAL_203 = ~_EVAL_101;
  assign _EVAL_145 = _EVAL_85 | _EVAL_76;
  assign _EVAL_247 = _EVAL_294 & _EVAL_119;
  assign _EVAL_64 = ~_EVAL_187;
  assign _EVAL_136 = _EVAL_225 | _EVAL_54;
  assign _EVAL_223 = ~_EVAL_248;
  assign _EVAL_269 = ~_EVAL_200;
  assign _EVAL_172 = ~_EVAL_99;
  assign _EVAL_282 = _EVAL_39 == 2'h0;
  assign _EVAL_240 = _EVAL_31 ? _EVAL_174 : 8'h0;
  assign _EVAL_147 = _EVAL_0[0];
  assign _EVAL_261 = _EVAL_7 & _EVAL_110;
  assign _EVAL_160 = _EVAL_14 & _EVAL_168;
  assign _EVAL_140 = _EVAL_136 >> _EVAL_16;
  assign _EVAL_239 = _EVAL_188 | _EVAL_222;
  assign _EVAL_77 = _EVAL_251[3:0];
  assign _EVAL_45 = ~_EVAL_263;
  assign _EVAL_71 = _EVAL_36 & _EVAL_59;
  assign _EVAL_202 = _EVAL_227 | _EVAL_8;
  assign _EVAL_36 = ~_EVAL_162;
  assign _EVAL_273 = _EVAL_173 | _EVAL_19;
  assign _EVAL_154 = _EVAL_3 == 3'h0;
  assign _EVAL_150 = ~_EVAL_15;
  assign _EVAL_20 = _EVAL_6 & _EVAL_27;
  assign _EVAL_155 = _EVAL_38 | _EVAL_223;
  assign _EVAL_199 = {1'b0,$signed(_EVAL_123)};
  assign _EVAL_188 = _EVAL_244 == 2'h1;
  assign _EVAL_97 = _EVAL_139 | _EVAL_8;
  assign _EVAL_110 = {{25'd0}, _EVAL_192};
  assign _EVAL_216 = _EVAL_102 & _EVAL_162;
  assign _EVAL_252 = ~_EVAL_280;
  assign _EVAL_213 = _EVAL_11 >= 3'h2;
  assign _EVAL_138 = ~_EVAL_178;
  assign _EVAL_128 = _EVAL_6 & _EVAL_204;
  assign _EVAL_111 = ~_EVAL_234;
  assign _EVAL_95 = _EVAL_237 | _EVAL_8;
  assign _EVAL_189 = _EVAL_14 & _EVAL_120;
  assign _EVAL_37 = ~_EVAL_49;
  assign _EVAL_103 = _EVAL_86 | _EVAL_8;
  assign _EVAL_127 = _EVAL_113 | _EVAL_8;
  assign _EVAL_62 = _EVAL_6 & _EVAL_196;
  assign _EVAL_218 = _EVAL_3 == _EVAL_291;
  assign _EVAL_234 = _EVAL_247 | _EVAL_8;
  assign _EVAL_257 = _EVAL_150 == 4'h0;
  assign _EVAL_190 = ~_EVAL_22;
  assign _EVAL_152 = ~_EVAL_44;
  assign _EVAL_109 = _EVAL_40 | _EVAL_8;
  assign _EVAL_57 = 13'h3f << _EVAL_11;
  assign _EVAL_225 = _EVAL_201[4:0];
  assign _EVAL_74 = _EVAL_184 | _EVAL_8;
  assign _EVAL_271 = _EVAL_11 == _EVAL_105;
  assign _EVAL_96 = _EVAL_281 | _EVAL_8;
  assign _EVAL_87 = ~_EVAL_266;
  assign _EVAL_263 = _EVAL_218 | _EVAL_8;
  assign _EVAL_266 = _EVAL_166 | _EVAL_8;
  assign _EVAL_41 = ~_EVAL_95;
  assign _EVAL_114 = _EVAL_3 == 3'h7;
  assign _EVAL_29 = _EVAL_236 & _EVAL_81;
  assign _EVAL_262 = ~_EVAL_202;
  assign _EVAL_90 = _EVAL_239 | _EVAL_278;
  assign _EVAL_212 = {_EVAL_265,_EVAL_24,_EVAL_115,_EVAL_273};
  assign _EVAL_84 = _EVAL_220 | _EVAL_8;
  assign _EVAL_176 = ~_EVAL_131;
  assign _EVAL_164 = _EVAL_89 | _EVAL_8;
  assign _EVAL_165 = _EVAL_158[3:0];
  assign _EVAL_148 = 8'h1 << _EVAL_4;
  assign _EVAL_159 = _EVAL_54 | _EVAL_225;
  assign _EVAL_40 = _EVAL_12 <= 3'h4;
  assign _EVAL_187 = _EVAL_142 | _EVAL_8;
  assign _EVAL_139 = _EVAL_140[0];
  assign _EVAL_163 = _EVAL_73;
  assign _EVAL_106 = _EVAL_12 <= 3'h1;
  assign _EVAL_99 = _EVAL_240[4:0];
  assign _EVAL_274 = ~_EVAL_182;
  assign _EVAL_23 = ~_EVAL_221;
  assign _EVAL_93 = _EVAL_292 - 4'h1;
  assign _EVAL_26 = _EVAL_14 & _EVAL_235;
  assign _EVAL_115 = _EVAL_173 | _EVAL_268;
  assign _EVAL_231 = ~_EVAL_283;
  assign _EVAL_241 = ~_EVAL_82;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_28 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_54 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_105 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_124 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_133 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_135 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_144 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_146 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_161 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_211 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_215 = _RAND_10[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_224 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_229 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_260 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_272 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_291 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_292 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_10) begin
    if (_EVAL_277) begin
      _EVAL_28 <= _EVAL_0;
    end
    if (_EVAL_8) begin
      _EVAL_54 <= 5'h0;
    end else begin
      _EVAL_54 <= _EVAL_33;
    end
    if (_EVAL_198) begin
      _EVAL_105 <= _EVAL_11;
    end
    if (_EVAL_277) begin
      _EVAL_124 <= _EVAL_4;
    end
    if (_EVAL_198) begin
      _EVAL_133 <= _EVAL_1;
    end
    if (_EVAL_198) begin
      _EVAL_135 <= _EVAL_16;
    end
    if (_EVAL_198) begin
      _EVAL_144 <= _EVAL_5;
    end
    if (_EVAL_8) begin
      _EVAL_146 <= 4'h0;
    end else if (_EVAL_85) begin
      if (_EVAL_79) begin
        if (_EVAL_60) begin
          _EVAL_146 <= _EVAL_270;
        end else begin
          _EVAL_146 <= 4'h0;
        end
      end else begin
        _EVAL_146 <= _EVAL_165;
      end
    end
    if (_EVAL_8) begin
      _EVAL_161 <= 32'h0;
    end else if (_EVAL_145) begin
      _EVAL_161 <= 32'h0;
    end else begin
      _EVAL_161 <= _EVAL_83;
    end
    if (_EVAL_8) begin
      _EVAL_211 <= 4'h0;
    end else if (_EVAL_76) begin
      if (_EVAL_258) begin
        if (_EVAL_243) begin
          _EVAL_211 <= _EVAL_170;
        end else begin
          _EVAL_211 <= 4'h0;
        end
      end else begin
        _EVAL_211 <= _EVAL_77;
      end
    end
    if (_EVAL_277) begin
      _EVAL_215 <= _EVAL_7;
    end
    if (_EVAL_277) begin
      _EVAL_224 <= _EVAL_12;
    end
    if (_EVAL_8) begin
      _EVAL_229 <= 4'h0;
    end else if (_EVAL_76) begin
      if (_EVAL_51) begin
        if (_EVAL_243) begin
          _EVAL_229 <= _EVAL_170;
        end else begin
          _EVAL_229 <= 4'h0;
        end
      end else begin
        _EVAL_229 <= _EVAL_129;
      end
    end
    if (_EVAL_198) begin
      _EVAL_260 <= _EVAL_2;
    end
    if (_EVAL_198) begin
      _EVAL_272 <= _EVAL_17;
    end
    if (_EVAL_277) begin
      _EVAL_291 <= _EVAL_3;
    end
    if (_EVAL_8) begin
      _EVAL_292 <= 4'h0;
    end else if (_EVAL_85) begin
      if (_EVAL_177) begin
        if (_EVAL_60) begin
          _EVAL_292 <= _EVAL_270;
        end else begin
          _EVAL_292 <= 4'h0;
        end
      end else begin
        _EVAL_292 <= _EVAL_78;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c453e93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bb966f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55c64379)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6f1616e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b76f52d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d30fdbc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ce68870)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cb87bf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87f6c1f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3db870d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de4f7044)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46855bab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(348edefe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cc790d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f721f2da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(132eb8c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8de6ccab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11e6a41c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8511dbfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23f0d0eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d3aaa50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2cdd3e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a33c2750)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95abb7c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f87b9ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(838b8227)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d18cc9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf652462)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18d04357)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e355979)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33e580e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27ec16e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4baab8bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea6a2753)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4128b46b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d79b5a8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d6cd263)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb10b563)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f352c46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b57e530c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31e8f82c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_255) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19a37425)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5260c9e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1292e2e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1341f9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6270016)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48ae5507)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db496915)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(898026bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6ae0142)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94a100ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c2c28a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bab55e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc87850f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cd4908a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_274) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89b6e733)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7949eb65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8aaf0a84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69292c9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10a1a41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8697490)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60d9a538)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2cf342a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17066053)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7c3d417)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d7b8b6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce55d102)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aeea1a27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b52c267)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(392c1af7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e9aa495)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b9b61bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12a519c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46e987a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df7289e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_274) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb9f1138)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0569570)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce421ddf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_255) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27b0a6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e93557b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b49aef20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d439edd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78a4af06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16e39e0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab779d75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f43c5305)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_143 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d98f173f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd081c58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df3751d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13061bc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35e993da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(310af077)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72f091b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
