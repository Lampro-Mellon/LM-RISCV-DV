//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_169(
  input  [31:0] _EVAL,
  input         _EVAL_0,
  output        _EVAL_1,
  input  [1:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  output [2:0]  _EVAL_4,
  input         _EVAL_5,
  output [2:0]  _EVAL_6,
  output        _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  output [2:0]  _EVAL_11,
  output [1:0]  _EVAL_12,
  input         _EVAL_13,
  output [1:0]  _EVAL_14,
  output [3:0]  _EVAL_15,
  output [31:0] _EVAL_16,
  output [31:0] _EVAL_17,
  input         _EVAL_18,
  input  [1:0]  _EVAL_19,
  output        _EVAL_20,
  output        _EVAL_21,
  input  [31:0] _EVAL_22,
  input  [31:0] _EVAL_23,
  output        _EVAL_24,
  input  [2:0]  _EVAL_25,
  output [31:0] _EVAL_26,
  input  [3:0]  _EVAL_27,
  output [2:0]  _EVAL_28,
  input  [2:0]  _EVAL_29,
  input         _EVAL_30,
  input  [2:0]  _EVAL_31,
  output [2:0]  _EVAL_32
);
  assign _EVAL_6 = _EVAL_31;
  assign _EVAL_12 = _EVAL_2;
  assign _EVAL_4 = _EVAL_9;
  assign _EVAL_26 = _EVAL;
  assign _EVAL_1 = _EVAL_18;
  assign _EVAL_7 = _EVAL_30;
  assign _EVAL_20 = _EVAL_0;
  assign _EVAL_17 = _EVAL_23;
  assign _EVAL_21 = _EVAL_13;
  assign _EVAL_16 = _EVAL_22;
  assign _EVAL_32 = _EVAL_29;
  assign _EVAL_11 = _EVAL_25;
  assign _EVAL_15 = _EVAL_27;
  assign _EVAL_24 = _EVAL_8;
  assign _EVAL_28 = _EVAL_3;
  assign _EVAL_14 = _EVAL_19;
endmodule
