//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_98_assert(
  input         _EVAL,
  input  [1:0]  _EVAL_0,
  input  [1:0]  _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [14:0] _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [2:0]  _EVAL_13,
  input  [3:0]  _EVAL_14
);
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire [3:0] _EVAL_23;
  reg [2:0] _EVAL_24;
  reg [31:0] _RAND_0;
  reg [14:0] _EVAL_25;
  reg [31:0] _RAND_1;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire [4:0] _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire [15:0] _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire [4:0] _EVAL_53;
  wire  _EVAL_55;
  wire [3:0] _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire [1:0] _EVAL_63;
  wire [14:0] _EVAL_64;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire [15:0] _EVAL_76;
  wire [31:0] _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire [4:0] _EVAL_80;
  wire  _EVAL_81;
  wire [4:0] _EVAL_82;
  reg [2:0] _EVAL_83;
  reg [31:0] _RAND_2;
  wire  _EVAL_84;
  wire [15:0] _EVAL_85;
  wire  _EVAL_86;
  wire [4:0] _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire [1:0] _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire [1:0] _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire [3:0] _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  reg [1:0] _EVAL_103;
  reg [31:0] _RAND_3;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire [7:0] _EVAL_111;
  reg [2:0] _EVAL_112;
  reg [31:0] _RAND_4;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire [1:0] _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  reg [2:0] _EVAL_129;
  reg [31:0] _RAND_5;
  wire [31:0] plusarg_reader_out;
  wire [7:0] _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire [14:0] _EVAL_138;
  wire  _EVAL_139;
  wire [1:0] _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire [4:0] _EVAL_145;
  wire  _EVAL_147;
  wire  _EVAL_149;
  reg [1:0] _EVAL_150;
  reg [31:0] _RAND_6;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  reg  _EVAL_175;
  reg [31:0] _RAND_7;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire [3:0] _EVAL_181;
  wire [1:0] _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  reg [4:0] _EVAL_189;
  reg [31:0] _RAND_8;
  wire  _EVAL_190;
  wire  _EVAL_192;
  wire [32:0] _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire [14:0] _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  reg  _EVAL_209;
  reg [31:0] _RAND_9;
  wire [4:0] _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  reg  _EVAL_214;
  reg [31:0] _RAND_10;
  wire [1:0] _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire [1:0] _EVAL_218;
  wire [7:0] _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire [1:0] _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire [1:0] _EVAL_230;
  wire  _EVAL_231;
  reg [31:0] _EVAL_232;
  reg [31:0] _RAND_11;
  wire [4:0] _EVAL_233;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire [7:0] _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  reg  _EVAL_243;
  reg [31:0] _RAND_12;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  reg [2:0] _EVAL_249;
  reg [31:0] _RAND_13;
  wire [4:0] _EVAL_250;
  wire  _EVAL_251;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_231 = _EVAL_170 | _EVAL_10;
  assign _EVAL_241 = _EVAL_5 & _EVAL_206;
  assign _EVAL_40 = ~_EVAL_153;
  assign _EVAL_233 = 5'h3 << _EVAL_0;
  assign _EVAL_50 = {1'b0,$signed(_EVAL_64)};
  assign _EVAL_187 = _EVAL_3 == 3'h7;
  assign _EVAL_217 = ~_EVAL_137;
  assign _EVAL_48 = _EVAL_13 != 3'h0;
  assign _EVAL_104 = ~_EVAL_160;
  assign _EVAL_247 = _EVAL_93 | _EVAL_242;
  assign _EVAL_204 = _EVAL_8 & _EVAL_138;
  assign _EVAL_250 = _EVAL_189 | _EVAL_53;
  assign _EVAL_124 = _EVAL_243 - 1'h1;
  assign _EVAL_96 = ~_EVAL_156;
  assign _EVAL_88 = ~_EVAL_227;
  assign _EVAL_113 = _EVAL_6 & _EVAL_15;
  assign _EVAL_97 = ~_EVAL_78;
  assign _EVAL_46 = _EVAL_171 & _EVAL_225;
  assign _EVAL_105 = _EVAL_90[0];
  assign _EVAL_99 = ~_EVAL_243;
  assign _EVAL_120 = _EVAL_124[0];
  assign _EVAL_108 = _EVAL_171 & _EVAL_99;
  assign _EVAL_125 = _EVAL_39 & _EVAL_47;
  assign _EVAL_183 = _EVAL_5 & _EVAL_186;
  assign _EVAL_248 = _EVAL_30 | _EVAL_10;
  assign _EVAL_57 = $signed(_EVAL_85) == 16'sh0;
  assign _EVAL_21 = _EVAL_43 | _EVAL_10;
  assign _EVAL_210 = _EVAL_250 & _EVAL_80;
  assign _EVAL_134 = _EVAL_161 | _EVAL_79;
  assign _EVAL_196 = _EVAL_179 | _EVAL_10;
  assign _EVAL_123 = ~_EVAL_236;
  assign _EVAL_121 = _EVAL_12 == 3'h4;
  assign _EVAL_176 = _EVAL_134 | _EVAL_121;
  assign _EVAL_61 = _EVAL_102 & _EVAL_229;
  assign _EVAL_140 = _EVAL_214 - 1'h1;
  assign _EVAL_159 = ~_EVAL_35;
  assign _EVAL_67 = _EVAL_16 | _EVAL_235;
  assign _EVAL_76 = $signed(_EVAL_50) & -16'sh1000;
  assign _EVAL_147 = _EVAL_5 & _EVAL_69;
  assign _EVAL_143 = _EVAL_7 == 3'h4;
  assign _EVAL_185 = _EVAL_32 & _EVAL_122;
  assign _EVAL_190 = _EVAL_247 | _EVAL_10;
  assign _EVAL_84 = _EVAL_0 >= 2'h2;
  assign _EVAL_144 = _EVAL_173 | _EVAL_10;
  assign _EVAL_137 = _EVAL_116 | _EVAL_10;
  assign _EVAL_145 = _EVAL_219[4:0];
  assign _EVAL_227 = _EVAL_51 | _EVAL_10;
  assign _EVAL_153 = _EVAL_117 | _EVAL_10;
  assign _EVAL_27 = _EVAL_84 | _EVAL_125;
  assign _EVAL_188 = _EVAL_12 == _EVAL_129;
  assign _EVAL_19 = ~_EVAL_34;
  assign _EVAL_95 = _EVAL_4 == 3'h5;
  assign _EVAL_205 = _EVAL_208 | _EVAL_92;
  assign _EVAL_149 = _EVAL_3 == 3'h4;
  assign _EVAL_128 = ~_EVAL_62;
  assign _EVAL_164 = _EVAL_94[0];
  assign _EVAL_163 = _EVAL_6 & _EVAL_95;
  assign _EVAL_63 = _EVAL_233[1:0];
  assign _EVAL_117 = _EVAL_38 & _EVAL_57;
  assign _EVAL_82 = _EVAL_37 >> _EVAL_7;
  assign _EVAL_162 = _EVAL_3 == 3'h3;
  assign _EVAL_44 = _EVAL_5 & _EVAL_187;
  assign _EVAL_38 = _EVAL_0 <= 2'h2;
  assign _EVAL_79 = _EVAL_182 == 2'h0;
  assign _EVAL_166 = _EVAL_3 == 3'h5;
  assign _EVAL_220 = _EVAL_1 == _EVAL_150;
  assign _EVAL_180 = _EVAL_3 == 3'h2;
  assign _EVAL_15 = _EVAL_4 == 3'h6;
  assign _EVAL_17 = ~_EVAL_66;
  assign _EVAL_100 = _EVAL_6 & _EVAL_224;
  assign _EVAL_56 = ~_EVAL_98;
  assign _EVAL_240 = ~_EVAL_10;
  assign _EVAL_109 = _EVAL_39 & _EVAL_154;
  assign _EVAL_75 = _EVAL_0[0];
  assign _EVAL_91 = _EVAL_5 & _EVAL_166;
  assign _EVAL_181 = _EVAL_14 & _EVAL_56;
  assign _EVAL_111 = 8'h1 << _EVAL_12;
  assign _EVAL_167 = _EVAL_6 & _EVAL_31;
  assign _EVAL_225 = ~_EVAL_214;
  assign _EVAL_141 = _EVAL_154 & _EVAL_128;
  assign _EVAL_59 = ~_EVAL_245;
  assign _EVAL_223 = _EVAL_32 & _EVAL_68;
  assign _EVAL_35 = _EVAL_70 | _EVAL_10;
  assign _EVAL_192 = _EVAL_97 | _EVAL_10;
  assign _EVAL_26 = _EVAL_3 == _EVAL_112;
  assign _EVAL_130 = _EVAL_108 ? _EVAL_111 : 8'h0;
  assign _EVAL_62 = _EVAL_8[0];
  assign _EVAL_224 = _EVAL_4 == 3'h1;
  assign _EVAL_160 = _EVAL_48 | _EVAL_10;
  assign _EVAL_107 = _EVAL_4 == _EVAL_83;
  assign _EVAL_156 = _EVAL_176 | _EVAL_10;
  assign _EVAL_218 = _EVAL_226 | 2'h1;
  assign _EVAL_80 = ~_EVAL_145;
  assign _EVAL_242 = ~_EVAL_244;
  assign _EVAL_221 = ~_EVAL_172;
  assign _EVAL_16 = _EVAL_84 | _EVAL_109;
  assign _EVAL_81 = _EVAL_13 <= 3'h1;
  assign _EVAL_215 = ~_EVAL_63;
  assign _EVAL_216 = ~_EVAL_213;
  assign _EVAL_161 = _EVAL_182 == 2'h1;
  assign _EVAL_133 = _EVAL_211 | _EVAL_10;
  assign _EVAL_246 = _EVAL_26 | _EVAL_10;
  assign _EVAL_238 = 8'h1 << _EVAL_7;
  assign _EVAL_135 = _EVAL_0 == _EVAL_103;
  assign _EVAL_90 = _EVAL_175 - 1'h1;
  assign _EVAL_139 = ~_EVAL_22;
  assign _EVAL_229 = ~_EVAL_15;
  assign _EVAL_142 = _EVAL_4 == 3'h0;
  assign _EVAL_235 = _EVAL_32 & _EVAL_141;
  assign _EVAL_171 = _EVAL & _EVAL_5;
  assign _EVAL_102 = _EVAL_222 & _EVAL_178;
  assign _EVAL_55 = plusarg_reader_out == 32'h0;
  assign _EVAL_118 = _EVAL_32 & _EVAL_152;
  assign _EVAL_169 = ~_EVAL_144;
  assign _EVAL_33 = _EVAL_4 <= 3'h6;
  assign _EVAL_211 = _EVAL_181 == 4'h0;
  assign _EVAL_195 = ~_EVAL_60;
  assign _EVAL_47 = ~_EVAL_154;
  assign _EVAL_58 = ~_EVAL_197;
  assign _EVAL_228 = ~_EVAL_190;
  assign _EVAL_86 = _EVAL_131 | _EVAL_55;
  assign _EVAL_70 = _EVAL_1 >= 2'h2;
  assign _EVAL_49 = _EVAL_232 < plusarg_reader_out;
  assign _EVAL_36 = _EVAL_33 | _EVAL_10;
  assign _EVAL_94 = _EVAL_209 - 1'h1;
  assign _EVAL_194 = _EVAL_232 + 32'h1;
  assign _EVAL_98 = {_EVAL_132,_EVAL_67,_EVAL_203,_EVAL_71};
  assign _EVAL_154 = _EVAL_8[1];
  assign _EVAL_101 = _EVAL_6 & _EVAL_202;
  assign _EVAL_52 = _EVAL_171 | _EVAL_222;
  assign _EVAL_23 = ~_EVAL_14;
  assign _EVAL_201 = _EVAL_13 <= 3'h4;
  assign _EVAL_92 = _EVAL_230 == 2'h0;
  assign _EVAL_89 = ~_EVAL_175;
  assign _EVAL_244 = _EVAL_53 != 5'h0;
  assign _EVAL_68 = _EVAL_47 & _EVAL_62;
  assign _EVAL_78 = _EVAL_87[0];
  assign _EVAL_32 = _EVAL_218[0];
  assign _EVAL_173 = _EVAL_8 == _EVAL_25;
  assign _EVAL_186 = _EVAL_3 == 3'h0;
  assign _EVAL_251 = ~_EVAL_36;
  assign _EVAL_69 = _EVAL_3 == 3'h1;
  assign _EVAL_213 = _EVAL_119 | _EVAL_10;
  assign _EVAL_177 = _EVAL_157 | _EVAL_10;
  assign _EVAL_60 = _EVAL_188 | _EVAL_10;
  assign _EVAL_178 = ~_EVAL_209;
  assign _EVAL_198 = _EVAL_5 & _EVAL_149;
  assign _EVAL_239 = ~_EVAL_246;
  assign _EVAL_174 = _EVAL_5 & _EVAL_110;
  assign _EVAL_53 = _EVAL_130[4:0];
  assign _EVAL_222 = _EVAL_2 & _EVAL_6;
  assign _EVAL_170 = _EVAL_7 == _EVAL_24;
  assign _EVAL_197 = _EVAL_41 | _EVAL_10;
  assign _EVAL_152 = _EVAL_47 & _EVAL_128;
  assign _EVAL_93 = _EVAL_53 != _EVAL_145;
  assign _EVAL_39 = _EVAL_218[1];
  assign _EVAL_236 = _EVAL_220 | _EVAL_10;
  assign _EVAL_29 = _EVAL_5 & _EVAL_180;
  assign _EVAL_203 = _EVAL_27 | _EVAL_223;
  assign _EVAL_212 = ~_EVAL_21;
  assign _EVAL_74 = _EVAL_86 | _EVAL_49;
  assign _EVAL_41 = _EVAL_13 <= 3'h3;
  assign _EVAL_200 = ~_EVAL_199;
  assign _EVAL_71 = _EVAL_27 | _EVAL_118;
  assign _EVAL_155 = _EVAL_140[0];
  assign _EVAL_106 = ~_EVAL_192;
  assign _EVAL_85 = _EVAL_76;
  assign _EVAL_158 = _EVAL_81 | _EVAL_10;
  assign _EVAL_87 = _EVAL_189 >> _EVAL_12;
  assign _EVAL_114 = _EVAL_4 == 3'h4;
  assign _EVAL_179 = _EVAL_14 == _EVAL_98;
  assign _EVAL_28 = _EVAL_42 | _EVAL_10;
  assign _EVAL_157 = _EVAL_13 == _EVAL_249;
  assign _EVAL_136 = ~_EVAL_158;
  assign _EVAL_22 = _EVAL_201 | _EVAL_10;
  assign _EVAL_199 = _EVAL_107 | _EVAL_10;
  assign _EVAL_226 = 2'h1 << _EVAL_75;
  assign _EVAL_165 = _EVAL_6 & _EVAL_114;
  assign _EVAL_73 = _EVAL_13 <= 3'h2;
  assign _EVAL_30 = _EVAL_205 | _EVAL_143;
  assign _EVAL_119 = _EVAL_204 == 15'h0;
  assign _EVAL_151 = _EVAL_189 != 5'h0;
  assign _EVAL_208 = _EVAL_230 == 2'h1;
  assign _EVAL_64 = _EVAL_8 ^ 15'h4000;
  assign _EVAL_34 = _EVAL_73 | _EVAL_10;
  assign _EVAL_66 = _EVAL_135 | _EVAL_10;
  assign _EVAL_245 = _EVAL_74 | _EVAL_10;
  assign _EVAL_110 = _EVAL_3 == 3'h6;
  assign _EVAL_184 = ~_EVAL_133;
  assign _EVAL_42 = _EVAL_82[0];
  assign _EVAL_43 = ~_EVAL_9;
  assign _EVAL_219 = _EVAL_61 ? _EVAL_238 : 8'h0;
  assign _EVAL_207 = _EVAL_6 & _EVAL_142;
  assign _EVAL_138 = {{13'd0}, _EVAL_215};
  assign _EVAL_115 = ~_EVAL_248;
  assign _EVAL_31 = ~_EVAL_89;
  assign _EVAL_230 = _EVAL_7[2:1];
  assign _EVAL_18 = _EVAL_222 & _EVAL_89;
  assign _EVAL_45 = _EVAL_5 & _EVAL_162;
  assign _EVAL_206 = ~_EVAL_225;
  assign _EVAL_77 = _EVAL_194[31:0];
  assign _EVAL_37 = _EVAL_53 | _EVAL_189;
  assign _EVAL_168 = ~_EVAL_231;
  assign _EVAL_51 = _EVAL_13 == 3'h0;
  assign _EVAL_72 = ~_EVAL_177;
  assign _EVAL_122 = _EVAL_154 & _EVAL_62;
  assign _EVAL_131 = ~_EVAL_151;
  assign _EVAL_127 = ~_EVAL_196;
  assign _EVAL_132 = _EVAL_16 | _EVAL_185;
  assign _EVAL_202 = _EVAL_4 == 3'h2;
  assign _EVAL_126 = ~_EVAL_28;
  assign _EVAL_172 = _EVAL_84 | _EVAL_10;
  assign _EVAL_182 = _EVAL_12[2:1];
  assign _EVAL_116 = _EVAL_23 == 4'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_24 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_25 = _RAND_1[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_83 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_103 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_112 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_129 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_150 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_175 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_189 = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_209 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_214 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_232 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_243 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_249 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_11) begin
    if (_EVAL_18) begin
      _EVAL_24 <= _EVAL_7;
    end
    if (_EVAL_46) begin
      _EVAL_25 <= _EVAL_8;
    end
    if (_EVAL_18) begin
      _EVAL_83 <= _EVAL_4;
    end
    if (_EVAL_46) begin
      _EVAL_103 <= _EVAL_0;
    end
    if (_EVAL_46) begin
      _EVAL_112 <= _EVAL_3;
    end
    if (_EVAL_46) begin
      _EVAL_129 <= _EVAL_12;
    end
    if (_EVAL_18) begin
      _EVAL_150 <= _EVAL_1;
    end
    if (_EVAL_10) begin
      _EVAL_175 <= 1'h0;
    end else if (_EVAL_222) begin
      if (_EVAL_89) begin
        _EVAL_175 <= 1'h0;
      end else begin
        _EVAL_175 <= _EVAL_105;
      end
    end
    if (_EVAL_10) begin
      _EVAL_189 <= 5'h0;
    end else begin
      _EVAL_189 <= _EVAL_210;
    end
    if (_EVAL_10) begin
      _EVAL_209 <= 1'h0;
    end else if (_EVAL_222) begin
      if (_EVAL_178) begin
        _EVAL_209 <= 1'h0;
      end else begin
        _EVAL_209 <= _EVAL_164;
      end
    end
    if (_EVAL_10) begin
      _EVAL_214 <= 1'h0;
    end else if (_EVAL_171) begin
      if (_EVAL_225) begin
        _EVAL_214 <= 1'h0;
      end else begin
        _EVAL_214 <= _EVAL_155;
      end
    end
    if (_EVAL_10) begin
      _EVAL_232 <= 32'h0;
    end else if (_EVAL_52) begin
      _EVAL_232 <= 32'h0;
    end else begin
      _EVAL_232 <= _EVAL_77;
    end
    if (_EVAL_10) begin
      _EVAL_243 <= 1'h0;
    end else if (_EVAL_171) begin
      if (_EVAL_99) begin
        _EVAL_243 <= 1'h0;
      end else begin
        _EVAL_243 <= _EVAL_120;
      end
    end
    if (_EVAL_46) begin
      _EVAL_249 <= _EVAL_13;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dce3fa47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1597a73d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28a1f551)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ba0c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd83c825)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e8ced2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b19cbcd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ef0e486)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(541501c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(482570cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a6b53b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cf44291)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74d399c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1c68bc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac4746f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f2c7feb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f347e44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6dbac69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2307f04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae7c4b69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(439e3ce2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c655fc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eac7984a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d675a887)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d23d2c37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29ce1843)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(729b6116)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(656a0143)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7db784b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85359f97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1de931e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15c6a9f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abfa3cfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa059851)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_19) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28659f3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4636637c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4786bfe5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eaad4a86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aadfbd72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d50ea0dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15a45e7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59cdf34a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_19) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2b3ce73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de73467d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b14225da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56a92e6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a9a5121)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5907d71b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30c51e4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b18bc29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d99c2bac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d63302da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce32dbba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb3e36f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1dc8ed2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d5d2597)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7052f2fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19dc2154)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f69c2fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a7b72f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32711a50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8257548a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ae49839)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f114c20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c64bbb10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f9d79dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e538377)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7d8d315)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9d2b318)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6821be89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bb2f119)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed5ebbbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cada22aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
