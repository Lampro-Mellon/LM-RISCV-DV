//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_150(
  output [4:0]  _EVAL,
  output [4:0]  _EVAL_0,
  output        _EVAL_1,
  output [31:0] _EVAL_2,
  output [4:0]  _EVAL_3,
  input  [31:0] _EVAL_4
);
  wire [2:0] _EVAL_5;
  wire [31:0] _EVAL_6;
  wire [4:0] _EVAL_7;
  wire [31:0] _EVAL_8;
  wire [27:0] _EVAL_9;
  wire [4:0] _EVAL_10;
  wire  _EVAL_11;
  wire [4:0] _EVAL_12;
  wire  _EVAL_13;
  wire  _EVAL_14;
  wire [4:0] _EVAL_15;
  wire [4:0] _EVAL_16;
  wire  _EVAL_17;
  wire [2:0] _EVAL_18;
  wire [4:0] _EVAL_19;
  wire [4:0] _EVAL_20;
  wire [31:0] _EVAL_21;
  wire [4:0] _EVAL_22;
  wire [31:0] _EVAL_23;
  wire [1:0] _EVAL_24;
  wire [3:0] _EVAL_25;
  wire [4:0] _EVAL_26;
  wire [2:0] _EVAL_27;
  wire [27:0] _EVAL_28;
  wire [4:0] _EVAL_29;
  wire [27:0] _EVAL_30;
  wire [1:0] _EVAL_31;
  wire [4:0] _EVAL_32;
  wire [4:0] _EVAL_33;
  wire [31:0] _EVAL_34;
  wire [2:0] _EVAL_35;
  wire [2:0] _EVAL_36;
  wire [26:0] _EVAL_37;
  wire  _EVAL_38;
  wire [24:0] _EVAL_39;
  wire [4:0] _EVAL_40;
  wire [31:0] _EVAL_41;
  wire [4:0] _EVAL_42;
  wire  _EVAL_43;
  wire [2:0] _EVAL_44;
  wire [4:0] _EVAL_45;
  wire [4:0] _EVAL_46;
  wire [9:0] _EVAL_47;
  wire [31:0] _EVAL_48;
  wire [4:0] _EVAL_49;
  wire [24:0] _EVAL_50;
  wire  _EVAL_51;
  wire [4:0] _EVAL_52;
  wire [4:0] _EVAL_53;
  wire [4:0] _EVAL_54;
  wire [4:0] _EVAL_55;
  wire [4:0] _EVAL_56;
  wire [4:0] _EVAL_57;
  wire [14:0] _EVAL_58;
  wire [4:0] _EVAL_59;
  wire [31:0] _EVAL_60;
  wire [27:0] _EVAL_61;
  wire [3:0] _EVAL_62;
  wire [7:0] _EVAL_63;
  wire  _EVAL_64;
  wire [31:0] _EVAL_65;
  wire [4:0] _EVAL_66;
  wire [1:0] _EVAL_67;
  wire [30:0] _EVAL_68;
  wire [31:0] _EVAL_69;
  wire [31:0] _EVAL_70;
  wire [4:0] _EVAL_71;
  wire  _EVAL_72;
  wire [4:0] _EVAL_73;
  wire [31:0] _EVAL_74;
  wire [6:0] _EVAL_75;
  wire [31:0] _EVAL_76;
  wire [4:0] _EVAL_77;
  wire  _EVAL_78;
  wire [8:0] _EVAL_79;
  wire  _EVAL_80;
  wire [31:0] _EVAL_81;
  wire [31:0] _EVAL_82;
  wire [4:0] _EVAL_83;
  wire [31:0] _EVAL_84;
  wire [4:0] _EVAL_85;
  wire [31:0] _EVAL_86;
  wire [4:0] _EVAL_87;
  wire  _EVAL_88;
  wire [4:0] _EVAL_89;
  wire [2:0] _EVAL_90;
  wire [4:0] _EVAL_91;
  wire [4:0] _EVAL_92;
  wire [2:0] _EVAL_93;
  wire  _EVAL_94;
  wire [31:0] _EVAL_95;
  wire [31:0] _EVAL_96;
  wire [4:0] _EVAL_97;
  wire  _EVAL_98;
  wire [4:0] _EVAL_99;
  wire [2:0] _EVAL_100;
  wire [31:0] _EVAL_101;
  wire [4:0] _EVAL_102;
  wire [4:0] _EVAL_103;
  wire [2:0] _EVAL_104;
  wire  _EVAL_105;
  wire [4:0] _EVAL_106;
  wire  _EVAL_107;
  wire [31:0] _EVAL_108;
  wire [31:0] _EVAL_109;
  wire [24:0] _EVAL_110;
  wire [3:0] _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire [31:0] _EVAL_114;
  wire [4:0] _EVAL_115;
  wire [31:0] _EVAL_116;
  wire [4:0] _EVAL_117;
  wire [31:0] _EVAL_118;
  wire [4:0] _EVAL_119;
  wire [31:0] _EVAL_120;
  wire [4:0] _EVAL_121;
  wire [4:0] _EVAL_122;
  wire [24:0] _EVAL_123;
  wire [5:0] _EVAL_124;
  wire [19:0] _EVAL_125;
  wire [11:0] _EVAL_126;
  wire [4:0] _EVAL_127;
  wire  _EVAL_128;
  wire [4:0] _EVAL_129;
  wire  _EVAL_130;
  wire [31:0] _EVAL_131;
  wire [31:0] _EVAL_132;
  wire [31:0] _EVAL_133;
  wire [31:0] _EVAL_134;
  wire [30:0] _EVAL_135;
  wire [4:0] _EVAL_136;
  wire [31:0] _EVAL_137;
  wire [4:0] _EVAL_138;
  wire [4:0] _EVAL_139;
  wire [31:0] _EVAL_140;
  wire  _EVAL_141;
  wire [31:0] _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire [31:0] _EVAL_145;
  wire [6:0] _EVAL_146;
  wire [31:0] _EVAL_147;
  wire [4:0] _EVAL_148;
  wire [4:0] _EVAL_149;
  wire  _EVAL_150;
  wire [24:0] _EVAL_151;
  wire  _EVAL_152;
  wire [4:0] _EVAL_153;
  wire  _EVAL_154;
  wire [24:0] _EVAL_155;
  wire [30:0] _EVAL_156;
  wire [31:0] _EVAL_157;
  wire [2:0] _EVAL_158;
  wire [4:0] _EVAL_159;
  wire [31:0] _EVAL_160;
  wire [4:0] _EVAL_161;
  wire [4:0] _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire [4:0] _EVAL_165;
  wire [4:0] _EVAL_166;
  wire  _EVAL_167;
  wire [4:0] _EVAL_168;
  wire [4:0] _EVAL_169;
  wire [2:0] _EVAL_170;
  wire [4:0] _EVAL_171;
  wire [1:0] _EVAL_172;
  wire [31:0] _EVAL_173;
  wire [31:0] _EVAL_174;
  wire [4:0] _EVAL_175;
  wire [4:0] _EVAL_176;
  wire [4:0] _EVAL_177;
  wire [2:0] _EVAL_178;
  wire [4:0] _EVAL_179;
  wire [4:0] _EVAL_180;
  wire  _EVAL_181;
  wire [4:0] _EVAL_182;
  wire  _EVAL_183;
  wire [6:0] _EVAL_184;
  wire  _EVAL_185;
  wire [4:0] _EVAL_186;
  wire  _EVAL_187;
  wire [24:0] _EVAL_188;
  wire [4:0] _EVAL_189;
  wire  _EVAL_190;
  wire [31:0] _EVAL_191;
  wire [4:0] _EVAL_192;
  wire [27:0] _EVAL_193;
  wire  _EVAL_194;
  wire [26:0] _EVAL_195;
  wire  _EVAL_196;
  wire [31:0] _EVAL_197;
  wire  _EVAL_198;
  wire [4:0] _EVAL_199;
  wire [7:0] _EVAL_200;
  wire [31:0] _EVAL_201;
  wire [4:0] _EVAL_202;
  wire [4:0] _EVAL_203;
  wire  _EVAL_204;
  wire [31:0] _EVAL_205;
  wire [31:0] _EVAL_206;
  wire  _EVAL_207;
  wire [4:0] _EVAL_208;
  wire [31:0] _EVAL_209;
  wire [31:0] _EVAL_210;
  wire [4:0] _EVAL_211;
  wire [4:0] _EVAL_212;
  wire  _EVAL_213;
  wire [31:0] _EVAL_214;
  wire [4:0] _EVAL_215;
  wire [4:0] _EVAL_216;
  wire [31:0] _EVAL_217;
  wire [4:0] _EVAL_218;
  wire [4:0] _EVAL_219;
  wire  _EVAL_220;
  wire [31:0] _EVAL_221;
  wire [4:0] _EVAL_222;
  wire [31:0] _EVAL_223;
  wire [7:0] _EVAL_224;
  wire [31:0] _EVAL_225;
  wire  _EVAL_226;
  wire [4:0] _EVAL_227;
  wire [30:0] _EVAL_228;
  wire [31:0] _EVAL_229;
  wire  _EVAL_230;
  wire [2:0] _EVAL_231;
  wire [31:0] _EVAL_232;
  wire [4:0] _EVAL_233;
  wire [31:0] _EVAL_234;
  wire [31:0] _EVAL_235;
  wire [31:0] _EVAL_236;
  wire [31:0] _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire [31:0] _EVAL_241;
  wire [4:0] _EVAL_242;
  wire [31:0] _EVAL_243;
  wire  _EVAL_244;
  wire [4:0] _EVAL_245;
  wire [6:0] _EVAL_246;
  wire [4:0] _EVAL_247;
  wire [4:0] _EVAL_248;
  wire [4:0] _EVAL_249;
  wire [20:0] _EVAL_250;
  wire [6:0] _EVAL_251;
  wire [1:0] _EVAL_252;
  wire [4:0] _EVAL_253;
  wire [4:0] _EVAL_254;
  wire [4:0] _EVAL_255;
  wire [30:0] _EVAL_256;
  wire [24:0] _EVAL_257;
  wire [4:0] _EVAL_258;
  wire [4:0] _EVAL_259;
  wire [31:0] _EVAL_260;
  wire [6:0] _EVAL_261;
  wire [28:0] _EVAL_262;
  wire [17:0] _EVAL_263;
  wire [27:0] _EVAL_264;
  wire [4:0] _EVAL_265;
  wire [26:0] _EVAL_266;
  wire [4:0] _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire [25:0] _EVAL_270;
  wire [4:0] _EVAL_271;
  wire [31:0] _EVAL_272;
  wire  _EVAL_273;
  wire [7:0] _EVAL_274;
  wire [1:0] _EVAL_275;
  wire [4:0] _EVAL_276;
  wire [31:0] _EVAL_277;
  wire [4:0] _EVAL_278;
  wire [4:0] _EVAL_279;
  wire [31:0] _EVAL_280;
  wire  _EVAL_281;
  wire [9:0] _EVAL_282;
  wire [24:0] _EVAL_283;
  wire [3:0] _EVAL_284;
  wire [2:0] _EVAL_285;
  wire [31:0] _EVAL_286;
  wire [1:0] _EVAL_287;
  wire [4:0] _EVAL_288;
  wire  _EVAL_289;
  wire [25:0] _EVAL_290;
  wire [4:0] _EVAL_291;
  wire [4:0] _EVAL_292;
  wire [4:0] _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire [24:0] _EVAL_296;
  wire [29:0] _EVAL_297;
  wire [4:0] _EVAL_298;
  wire [2:0] _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire [2:0] _EVAL_303;
  wire [12:0] _EVAL_304;
  wire [4:0] _EVAL_305;
  wire [26:0] _EVAL_306;
  wire [1:0] _EVAL_307;
  wire [6:0] _EVAL_308;
  wire [1:0] _EVAL_309;
  wire [28:0] _EVAL_310;
  wire [31:0] _EVAL_311;
  wire [26:0] _EVAL_312;
  wire [30:0] _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire [4:0] _EVAL_316;
  wire  _EVAL_317;
  assign _EVAL_146 = _EVAL_17 ? 7'h37 : 7'h3f;
  assign _EVAL_157 = _EVAL_167 ? _EVAL_4 : _EVAL_241;
  assign _EVAL_317 = _EVAL_36 == 3'h6;
  assign _EVAL_108 = {{7'd0}, _EVAL_257};
  assign _EVAL_57 = _EVAL_164 ? _EVAL_73 : _EVAL_32;
  assign _EVAL_180 = _EVAL_113 ? _EVAL_278 : _EVAL_85;
  assign _EVAL_106 = _EVAL_72 ? _EVAL_129 : _EVAL_215;
  assign _EVAL_311 = _EVAL_213 ? {{1'd0}, _EVAL_313} : _EVAL_147;
  assign _EVAL_9 = {_EVAL_252,_EVAL_80,_EVAL_231,2'h0,5'h2,3'h2,_EVAL_278,7'h7};
  assign _EVAL_291 = _EVAL_315 ? _EVAL_10 : _EVAL_136;
  assign _EVAL_256 = {{6'd0}, _EVAL_155};
  assign _EVAL_95 = {_EVAL_308,_EVAL_54,5'h0,3'h0,_EVAL_278,7'h13};
  assign _EVAL_228 = {{5'd0}, _EVAL_290};
  assign _EVAL_133 = _EVAL_315 ? _EVAL_280 : _EVAL_6;
  assign _EVAL_144 = _EVAL_216 == 5'h1e;
  assign _EVAL_150 = _EVAL_216 == 5'h2;
  assign _EVAL_107 = _EVAL_216 == 5'h1c;
  assign _EVAL_74 = _EVAL_163 ? _EVAL_4 : _EVAL_34;
  assign _EVAL_221 = _EVAL_113 ? _EVAL_101 : _EVAL_197;
  assign _EVAL_90 = _EVAL_4[15:13];
  assign _EVAL_222 = _EVAL_152 ? _EVAL_42 : _EVAL_233;
  assign _EVAL_117 = _EVAL_51 ? _EVAL_119 : _EVAL_305;
  assign _EVAL_18 = _EVAL_274[7:5];
  assign _EVAL_25 = _EVAL_79[8:5];
  assign _EVAL_19 = _EVAL_154 ? _EVAL_54 : _EVAL_20;
  assign _EVAL_267 = _EVAL_167 ? _EVAL_186 : _EVAL_171;
  assign _EVAL_262 = {_EVAL_104,_EVAL_80,_EVAL_24,3'h0,5'h2,3'h3,_EVAL_278,7'h7};
  assign _EVAL_253 = _EVAL_183 ? _EVAL_73 : _EVAL_40;
  assign _EVAL_207 = _EVAL_278 == 5'h2;
  assign _EVAL_79 = {_EVAL_27,_EVAL_158,3'h0};
  assign _EVAL_123 = {_EVAL_54,_EVAL_278,3'h0,12'he7};
  assign _EVAL_197 = _EVAL_94 ? _EVAL_174 : _EVAL_21;
  assign _EVAL_159 = _EVAL_63[4:0];
  assign _EVAL_13 = _EVAL_304[12];
  assign _EVAL_86 = {{2'd0}, _EVAL_297};
  assign _EVAL_139 = _EVAL_98 ? _EVAL_73 : _EVAL_259;
  assign _EVAL_23 = _EVAL_295 ? _EVAL_70 : _EVAL_145;
  assign _EVAL_110 = {_EVAL_54,_EVAL_278,3'h0,12'h67};
  assign _EVAL_289 = _EVAL_216 == 5'h5;
  assign _EVAL_191 = {{4'd0}, _EVAL_28};
  assign _EVAL_84 = {{7'd0}, _EVAL_188};
  assign _EVAL_293 = _EVAL_51 ? _EVAL_219 : _EVAL_57;
  assign _EVAL_48 = {_EVAL_268,_EVAL_47,_EVAL_244,_EVAL_200,5'h0,7'h6f};
  assign _EVAL_265 = _EVAL_269 ? _EVAL_54 : _EVAL_77;
  assign _EVAL_315 = _EVAL_216 == 5'h14;
  assign _EVAL_21 = _EVAL_98 ? _EVAL_137 : _EVAL_131;
  assign _EVAL_234 = _EVAL_152 ? _EVAL_311 : _EVAL_8;
  assign _EVAL_29 = _EVAL_315 ? _EVAL_71 : _EVAL_179;
  assign _EVAL_240 = _EVAL_36 == 3'h5;
  assign _EVAL_129 = _EVAL_4[24:20];
  assign _EVAL_116 = _EVAL_185 ? _EVAL_286 : _EVAL_229;
  assign _EVAL_114 = _EVAL_269 ? _EVAL_235 : _EVAL_217;
  assign _EVAL_38 = _EVAL_278 == 5'h0;
  assign _EVAL_270 = {_EVAL_80,_EVAL_54,_EVAL_278,3'h1,_EVAL_278,7'h13};
  assign _EVAL_232 = {{5'd0}, _EVAL_312};
  assign _EVAL_40 = _EVAL_185 ? _EVAL_73 : _EVAL_249;
  assign _EVAL_51 = _EVAL_216 == 5'hb;
  assign _EVAL_115 = _EVAL_141 ? _EVAL_54 : _EVAL_291;
  assign _EVAL_306 = {_EVAL_309,2'h1,_EVAL_104,2'h1,_EVAL_27,3'h2,_EVAL_22,7'h23};
  assign _EVAL_141 = _EVAL_216 == 5'h15;
  assign _EVAL_119 = _EVAL_194 ? _EVAL_278 : _EVAL_278;
  assign _EVAL_36 = {_EVAL_80,_EVAL_24};
  assign _EVAL_82 = _EVAL_239 ? _EVAL_48 : _EVAL_234;
  assign _EVAL_202 = _EVAL_107 ? _EVAL_278 : _EVAL_149;
  assign _EVAL_277 = {_EVAL_13,_EVAL_124,5'h0,2'h1,_EVAL_27,3'h1,_EVAL_111,_EVAL_204,7'h63};
  assign _EVAL_269 = _EVAL_216 == 5'h10;
  assign _EVAL_105 = _EVAL_36 == 3'h4;
  assign _EVAL_268 = _EVAL_250[20];
  assign _EVAL_211 = _EVAL_196 ? _EVAL_129 : _EVAL_106;
  assign _EVAL_53 = _EVAL_113 ? _EVAL_278 : _EVAL_15;
  assign _EVAL_254 = _EVAL_295 ? 5'h2 : _EVAL_166;
  assign _EVAL_188 = {_EVAL_54,5'h0,3'h0,_EVAL_278,7'h33};
  assign _EVAL_283 = _EVAL_281 ? _EVAL_123 : _EVAL_151;
  assign _EVAL_160 = {_EVAL_268,_EVAL_47,_EVAL_244,_EVAL_200,5'h1,7'h6f};
  assign _EVAL_242 = _EVAL_43 ? 5'h0 : _EVAL_278;
  assign _EVAL_109 = {_EVAL_5,_EVAL_307,_EVAL_301,_EVAL_190,_EVAL_300,4'h0,_EVAL_278,3'h0,_EVAL_278,_EVAL_251};
  assign _EVAL_226 = _EVAL_216 == 5'hf;
  assign _EVAL_33 = _EVAL_198 ? _EVAL_278 : _EVAL_92;
  assign _EVAL_2 = _EVAL_14 ? _EVAL_4 : _EVAL_120;
  assign _EVAL_280 = _EVAL_80 ? _EVAL_65 : _EVAL_206;
  assign _EVAL_210 = {_EVAL_125,_EVAL_278,_EVAL_146};
  assign _EVAL_239 = _EVAL_216 == 5'hd;
  assign _EVAL_11 = _EVAL_216 == 5'h11;
  assign _EVAL_229 = _EVAL_150 ? _EVAL_232 : _EVAL_140;
  assign _EVAL_67 = _EVAL_4[10:9];
  assign _EVAL_274 = {_EVAL_31,_EVAL_284,2'h0};
  assign _EVAL_113 = _EVAL_216 == 5'h8;
  assign _EVAL_70 = {{4'd0}, _EVAL_61};
  assign _EVAL_92 = _EVAL_154 ? _EVAL_278 : _EVAL_247;
  assign _EVAL_174 = {{5'd0}, _EVAL_266};
  assign _EVAL_101 = {_EVAL_308,_EVAL_54,_EVAL_278,3'h0,_EVAL_278,7'h13};
  assign _EVAL_54 = _EVAL_4[6:2];
  assign _EVAL_81 = {{4'd0}, _EVAL_9};
  assign _EVAL_1 = _EVAL_172 != 2'h3;
  assign _EVAL_88 = _EVAL_216 == 5'h17;
  assign _EVAL_216 = {_EVAL_172,_EVAL_90};
  assign _EVAL_248 = _EVAL_185 ? _EVAL_42 : _EVAL_121;
  assign _EVAL_285 = _EVAL_4[5:3];
  assign _EVAL_190 = _EVAL_4[2];
  assign _EVAL_0 = _EVAL_14 ? _EVAL_278 : _EVAL_192;
  assign _EVAL_279 = _EVAL_274[4:0];
  assign _EVAL_56 = _EVAL_163 ? _EVAL_129 : _EVAL_161;
  assign _EVAL_3 = _EVAL_14 ? _EVAL_186 : _EVAL_203;
  assign _EVAL_173 = {_EVAL_58,_EVAL_54,12'h0};
  assign _EVAL_121 = _EVAL_150 ? _EVAL_42 : _EVAL_99;
  assign _EVAL_245 = _EVAL_269 ? _EVAL_278 : _EVAL_49;
  assign _EVAL_30 = {_EVAL_252,_EVAL_80,_EVAL_231,2'h0,5'h2,3'h2,_EVAL_278,_EVAL_246};
  assign _EVAL_60 = _EVAL_88 ? _EVAL_237 : _EVAL_23;
  assign _EVAL_206 = _EVAL_43 ? _EVAL_84 : _EVAL_260;
  assign _EVAL_198 = _EVAL_216 == 5'h13;
  assign _EVAL_16 = _EVAL_112 ? _EVAL_42 : _EVAL_208;
  assign _EVAL_65 = _EVAL_43 ? _EVAL_108 : _EVAL_41;
  assign _EVAL_205 = _EVAL_11 ? _EVAL_209 : _EVAL_114;
  assign _EVAL_179 = _EVAL_198 ? 5'h2 : _EVAL_87;
  assign _EVAL_177 = _EVAL_113 ? _EVAL_73 : _EVAL_85;
  assign _EVAL_213 = _EVAL_275 == 2'h3;
  assign _EVAL_132 = _EVAL_112 ? _EVAL_223 : _EVAL_82;
  assign _EVAL_299 = _EVAL_105 ? 3'h0 : _EVAL_178;
  assign _EVAL_125 = _EVAL_173[31:12];
  assign _EVAL_272 = {{5'd0}, _EVAL_37};
  assign _EVAL_224 = _EVAL_4[12:5];
  assign _EVAL_122 = _EVAL_80 ? _EVAL_91 : _EVAL_168;
  assign _EVAL_260 = {{7'd0}, _EVAL_296};
  assign _EVAL_127 = _EVAL_239 ? _EVAL_73 : _EVAL_148;
  assign _EVAL_183 = _EVAL_216 == 5'h4;
  assign _EVAL_288 = _EVAL_181 ? 5'h1 : _EVAL_180;
  assign _EVAL_52 = _EVAL_72 ? _EVAL_186 : _EVAL_66;
  assign _EVAL_68 = _EVAL_228 | 31'h40000000;
  assign _EVAL_103 = _EVAL_112 ? _EVAL_42 : _EVAL_46;
  assign _EVAL_305 = _EVAL_164 ? _EVAL_278 : _EVAL_288;
  assign _EVAL_27 = _EVAL_4[9:7];
  assign _EVAL_175 = _EVAL_43 ? _EVAL_54 : _EVAL_54;
  assign _EVAL_58 = _EVAL_80 ? 15'h7fff : 15'h0;
  assign _EVAL_124 = _EVAL_304[10:5];
  assign _EVAL_39 = {_EVAL_263,7'h73};
  assign _EVAL_241 = _EVAL_107 ? _EVAL_4 : _EVAL_74;
  assign _EVAL_243 = _EVAL_72 ? _EVAL_4 : _EVAL_60;
  assign _EVAL_73 = {2'h1,_EVAL_104};
  assign _EVAL_199 = _EVAL_164 ? 5'h0 : _EVAL_218;
  assign _EVAL_278 = _EVAL_4[11:7];
  assign _EVAL_307 = _EVAL_4[4:3];
  assign _EVAL_111 = _EVAL_304[4:1];
  assign _EVAL_257 = {_EVAL_54,_EVAL_278,3'h0,_EVAL_278,7'h33};
  assign _EVAL_99 = _EVAL_273 ? _EVAL_42 : 5'h2;
  assign _EVAL_246 = _EVAL_281 ? 7'h3 : 7'h1f;
  assign _EVAL_223 = {_EVAL_13,_EVAL_124,5'h0,2'h1,_EVAL_27,3'h0,_EVAL_111,_EVAL_204,7'h63};
  assign _EVAL_32 = _EVAL_181 ? _EVAL_73 : _EVAL_177;
  assign _EVAL_273 = _EVAL_216 == 5'h1;
  assign _EVAL_59 = _EVAL_295 ? _EVAL_278 : _EVAL_138;
  assign _EVAL_194 = _EVAL_38 | _EVAL_207;
  assign _EVAL_314 = _EVAL_216 == 5'h1a;
  assign _EVAL_263 = _EVAL_110[24:7];
  assign _EVAL_50 = {_EVAL_263,7'h1f};
  assign _EVAL_218 = _EVAL_181 ? _EVAL_278 : _EVAL_53;
  assign _EVAL_252 = _EVAL_4[3:2];
  assign _EVAL_182 = _EVAL_112 ? 5'h0 : _EVAL_127;
  assign _EVAL_76 = {_EVAL_308,_EVAL_54,2'h1,_EVAL_27,3'h7,2'h1,_EVAL_27,7'h13};
  assign _EVAL_151 = _EVAL_39 | 25'h100000;
  assign _EVAL_313 = _EVAL_256 | _EVAL_156;
  assign _EVAL_287 = _EVAL_4[12:11];
  assign _EVAL_192 = _EVAL_144 ? _EVAL_278 : _EVAL_162;
  assign _EVAL_301 = _EVAL_4[5];
  assign _EVAL_212 = _EVAL_314 ? _EVAL_186 : _EVAL_271;
  assign _EVAL_15 = _EVAL_94 ? _EVAL_42 : _EVAL_55;
  assign _EVAL_181 = _EVAL_216 == 5'h9;
  assign _EVAL_49 = _EVAL_226 ? 5'h0 : _EVAL_16;
  assign _EVAL_184 = _EVAL_80 ? 7'h3b : 7'h33;
  assign _EVAL_43 = _EVAL_54 != 5'h0;
  assign _EVAL_156 = _EVAL_143 ? 31'h40000000 : 31'h0;
  assign _EVAL_292 = _EVAL_196 ? _EVAL_278 : _EVAL_189;
  assign _EVAL_217 = _EVAL_226 ? _EVAL_277 : _EVAL_132;
  assign _EVAL_5 = _EVAL_80 ? 3'h7 : 3'h0;
  assign _EVAL_130 = _EVAL_275 == 2'h2;
  assign _EVAL_230 = _EVAL_4[7];
  assign _EVAL_131 = _EVAL_289 ? _EVAL_191 : _EVAL_236;
  assign _EVAL_154 = _EVAL_216 == 5'h12;
  assign _EVAL_304 = {_EVAL_12,_EVAL_24,_EVAL_190,_EVAL_275,_EVAL_307,1'h0};
  assign _EVAL_186 = _EVAL_4[19:15];
  assign _EVAL_204 = _EVAL_304[11];
  assign _EVAL_37 = {_EVAL_309,2'h1,_EVAL_104,2'h1,_EVAL_27,3'h2,_EVAL_22,7'h3f};
  assign _EVAL_275 = _EVAL_4[11:10];
  assign _EVAL_281 = _EVAL_278 != 5'h0;
  assign _EVAL_12 = _EVAL_80 ? 5'h1f : 5'h0;
  assign _EVAL_7 = _EVAL_269 ? _EVAL_278 : _EVAL_102;
  assign _EVAL_64 = _EVAL_36 == 3'h1;
  assign _EVAL_296 = _EVAL_281 ? _EVAL_110 : _EVAL_50;
  assign _EVAL_298 = _EVAL_315 ? _EVAL_122 : _EVAL_33;
  assign _EVAL_46 = _EVAL_239 ? _EVAL_42 : _EVAL_222;
  assign _EVAL_143 = _EVAL_24 == 2'h0;
  assign _EVAL_55 = _EVAL_98 ? _EVAL_42 : _EVAL_258;
  assign _EVAL_31 = _EVAL_4[8:7];
  assign _EVAL_168 = _EVAL_43 ? _EVAL_278 : 5'h0;
  assign _EVAL_91 = _EVAL_43 ? _EVAL_278 : 5'h1;
  assign _EVAL_135 = _EVAL_220 ? _EVAL_68 : {{5'd0}, _EVAL_290};
  assign _EVAL_66 = _EVAL_88 ? 5'h2 : _EVAL_254;
  assign _EVAL_34 = _EVAL_314 ? _EVAL_4 : _EVAL_225;
  assign _EVAL_155 = {2'h1,_EVAL_104,2'h1,_EVAL_27,_EVAL_100,2'h1,_EVAL_27,_EVAL_184};
  assign _EVAL_297 = {_EVAL_62,_EVAL_287,_EVAL_301,_EVAL_300,2'h0,5'h2,3'h0,2'h1,_EVAL_104,_EVAL_261};
  assign _EVAL_303 = _EVAL_64 ? 3'h4 : 3'h0;
  assign _EVAL_266 = {_EVAL_309,2'h1,_EVAL_104,2'h1,_EVAL_27,3'h2,_EVAL_22,7'h27};
  assign _EVAL_20 = _EVAL_11 ? _EVAL_54 : _EVAL_265;
  assign _EVAL_148 = _EVAL_152 ? _EVAL_73 : _EVAL_293;
  assign _EVAL_284 = _EVAL_4[12:9];
  assign _EVAL_94 = _EVAL_216 == 5'h7;
  assign _EVAL_35 = _EVAL_63[7:5];
  assign _EVAL_215 = _EVAL_88 ? _EVAL_54 : _EVAL_89;
  assign _EVAL_78 = _EVAL_36 == 3'h2;
  assign _EVAL_8 = _EVAL_51 ? _EVAL_134 : _EVAL_69;
  assign _EVAL_147 = _EVAL_130 ? _EVAL_76 : {{1'd0}, _EVAL_135};
  assign _EVAL_83 = _EVAL_88 ? _EVAL_278 : _EVAL_59;
  assign _EVAL_14 = _EVAL_216 == 5'h1f;
  assign _EVAL_137 = {{5'd0}, _EVAL_306};
  assign _EVAL_61 = {_EVAL_18,_EVAL_54,5'h2,3'h2,_EVAL_279,7'h23};
  assign _EVAL_220 = _EVAL_275 == 2'h1;
  assign _EVAL_309 = _EVAL_75[6:5];
  assign _EVAL_112 = _EVAL_216 == 5'he;
  assign _EVAL_316 = _EVAL_107 ? _EVAL_129 : _EVAL_56;
  assign _EVAL_290 = {_EVAL_80,_EVAL_54,2'h1,_EVAL_27,3'h5,2'h1,_EVAL_27,7'h13};
  assign _EVAL_187 = _EVAL_4[11];
  assign _EVAL_178 = _EVAL_238 ? 3'h7 : _EVAL_170;
  assign _EVAL_104 = _EVAL_4[4:2];
  assign _EVAL_126 = {_EVAL_308,_EVAL_54};
  assign _EVAL = _EVAL_14 ? _EVAL_129 : _EVAL_169;
  assign _EVAL_140 = _EVAL_273 ? _EVAL_118 : _EVAL_86;
  assign _EVAL_195 = {_EVAL_301,_EVAL_158,_EVAL_300,2'h0,2'h1,_EVAL_27,3'h2,2'h1,_EVAL_104,7'h7};
  assign _EVAL_225 = _EVAL_196 ? _EVAL_4 : _EVAL_243;
  assign _EVAL_165 = _EVAL_163 ? _EVAL_186 : _EVAL_212;
  assign _EVAL_244 = _EVAL_250[11];
  assign _EVAL_72 = _EVAL_216 == 5'h18;
  assign _EVAL_97 = _EVAL_79[4:0];
  assign _EVAL_196 = _EVAL_216 == 5'h19;
  assign _EVAL_77 = _EVAL_226 ? 5'h0 : _EVAL_182;
  assign _EVAL_136 = _EVAL_198 ? _EVAL_54 : _EVAL_19;
  assign _EVAL_233 = _EVAL_51 ? _EVAL_119 : _EVAL_199;
  assign _EVAL_152 = _EVAL_216 == 5'hc;
  assign _EVAL_22 = _EVAL_75[4:0];
  assign _EVAL_250 = {_EVAL_282,_EVAL_302,_EVAL_67,_EVAL_300,_EVAL_230,_EVAL_190,_EVAL_187,_EVAL_285,1'h0};
  assign _EVAL_96 = {{4'd0}, _EVAL_30};
  assign _EVAL_45 = _EVAL_273 ? _EVAL_73 : _EVAL_73;
  assign _EVAL_153 = _EVAL_152 ? _EVAL_42 : _EVAL_117;
  assign _EVAL_201 = {{3'd0}, _EVAL_310};
  assign _EVAL_145 = _EVAL_141 ? _EVAL_201 : _EVAL_133;
  assign _EVAL_10 = _EVAL_80 ? _EVAL_175 : _EVAL_175;
  assign _EVAL_26 = _EVAL_183 ? _EVAL_42 : _EVAL_248;
  assign _EVAL_62 = _EVAL_4[10:7];
  assign _EVAL_98 = _EVAL_216 == 5'h6;
  assign _EVAL_308 = _EVAL_80 ? 7'h7f : 7'h0;
  assign _EVAL_142 = _EVAL_181 ? _EVAL_160 : _EVAL_221;
  assign _EVAL_71 = _EVAL_80 ? _EVAL_176 : _EVAL_242;
  assign _EVAL_235 = {{6'd0}, _EVAL_270};
  assign _EVAL_128 = _EVAL_36 == 3'h7;
  assign _EVAL_163 = _EVAL_216 == 5'h1b;
  assign _EVAL_162 = _EVAL_167 ? _EVAL_278 : _EVAL_202;
  assign _EVAL_169 = _EVAL_144 ? _EVAL_129 : _EVAL_255;
  assign _EVAL_44 = _EVAL_317 ? 3'h2 : _EVAL_93;
  assign _EVAL_42 = {2'h1,_EVAL_27};
  assign _EVAL_259 = _EVAL_289 ? _EVAL_73 : _EVAL_253;
  assign _EVAL_87 = _EVAL_154 ? 5'h2 : _EVAL_227;
  assign _EVAL_41 = {{7'd0}, _EVAL_283};
  assign _EVAL_149 = _EVAL_163 ? _EVAL_278 : _EVAL_276;
  assign _EVAL_189 = _EVAL_72 ? _EVAL_278 : _EVAL_83;
  assign _EVAL_310 = {_EVAL_25,_EVAL_54,5'h2,3'h3,_EVAL_97,7'h27};
  assign _EVAL_214 = _EVAL_154 ? _EVAL_96 : _EVAL_205;
  assign _EVAL_17 = _EVAL_126 != 12'h0;
  assign _EVAL_100 = _EVAL_128 ? 3'h3 : _EVAL_44;
  assign _EVAL_89 = _EVAL_295 ? _EVAL_54 : _EVAL_115;
  assign _EVAL_172 = _EVAL_4[1:0];
  assign _EVAL_238 = _EVAL_36 == 3'h3;
  assign _EVAL_102 = _EVAL_226 ? _EVAL_42 : _EVAL_103;
  assign _EVAL_295 = _EVAL_216 == 5'h16;
  assign _EVAL_282 = _EVAL_80 ? 10'h3ff : 10'h0;
  assign _EVAL_118 = {{4'd0}, _EVAL_193};
  assign _EVAL_249 = _EVAL_150 ? _EVAL_73 : _EVAL_45;
  assign _EVAL_193 = {_EVAL_24,_EVAL_158,3'h0,2'h1,_EVAL_27,3'h3,2'h1,_EVAL_104,7'h7};
  assign _EVAL_200 = _EVAL_250[19:12];
  assign _EVAL_75 = {_EVAL_301,_EVAL_158,_EVAL_300,2'h0};
  assign _EVAL_164 = _EVAL_216 == 5'ha;
  assign _EVAL_203 = _EVAL_144 ? _EVAL_186 : _EVAL_267;
  assign _EVAL_236 = _EVAL_183 ? _EVAL_272 : _EVAL_116;
  assign _EVAL_176 = _EVAL_43 ? _EVAL_278 : _EVAL_278;
  assign _EVAL_167 = _EVAL_216 == 5'h1d;
  assign _EVAL_28 = {_EVAL_35,2'h1,_EVAL_104,2'h1,_EVAL_27,3'h3,_EVAL_159,7'h27};
  assign _EVAL_286 = {{5'd0}, _EVAL_195};
  assign _EVAL_24 = _EVAL_4[6:5];
  assign _EVAL_158 = _EVAL_4[12:10];
  assign _EVAL_209 = {{3'd0}, _EVAL_262};
  assign _EVAL_264 = {_EVAL_18,_EVAL_54,5'h2,3'h2,_EVAL_279,7'h27};
  assign _EVAL_134 = _EVAL_194 ? _EVAL_109 : _EVAL_210;
  assign _EVAL_6 = _EVAL_198 ? _EVAL_81 : _EVAL_214;
  assign _EVAL_120 = _EVAL_144 ? _EVAL_4 : _EVAL_157;
  assign _EVAL_251 = _EVAL_17 ? 7'h13 : 7'h1f;
  assign _EVAL_231 = _EVAL_4[6:4];
  assign _EVAL_69 = _EVAL_164 ? _EVAL_95 : _EVAL_142;
  assign _EVAL_258 = _EVAL_289 ? _EVAL_42 : _EVAL_26;
  assign _EVAL_276 = _EVAL_314 ? _EVAL_278 : _EVAL_292;
  assign _EVAL_166 = _EVAL_141 ? 5'h2 : _EVAL_29;
  assign _EVAL_138 = _EVAL_141 ? _EVAL_278 : _EVAL_298;
  assign _EVAL_47 = _EVAL_250[10:1];
  assign _EVAL_294 = _EVAL_224 != 8'h0;
  assign _EVAL_185 = _EVAL_216 == 5'h3;
  assign _EVAL_271 = _EVAL_196 ? _EVAL_186 : _EVAL_52;
  assign _EVAL_300 = _EVAL_4[6];
  assign _EVAL_261 = _EVAL_294 ? 7'h13 : 7'h1f;
  assign _EVAL_255 = _EVAL_167 ? _EVAL_129 : _EVAL_316;
  assign _EVAL_208 = _EVAL_239 ? 5'h0 : _EVAL_153;
  assign _EVAL_312 = {_EVAL_301,_EVAL_158,_EVAL_300,2'h0,2'h1,_EVAL_27,3'h2,2'h1,_EVAL_104,7'h3};
  assign _EVAL_302 = _EVAL_4[8];
  assign _EVAL_171 = _EVAL_107 ? _EVAL_186 : _EVAL_165;
  assign _EVAL_93 = _EVAL_240 ? 3'h0 : _EVAL_299;
  assign _EVAL_63 = {_EVAL_24,_EVAL_158,3'h0};
  assign _EVAL_85 = _EVAL_94 ? _EVAL_73 : _EVAL_139;
  assign _EVAL_227 = _EVAL_11 ? 5'h2 : _EVAL_7;
  assign _EVAL_237 = {{4'd0}, _EVAL_264};
  assign _EVAL_80 = _EVAL_4[12];
  assign _EVAL_161 = _EVAL_314 ? _EVAL_129 : _EVAL_211;
  assign _EVAL_219 = _EVAL_194 ? _EVAL_73 : _EVAL_73;
  assign _EVAL_170 = _EVAL_78 ? 3'h6 : _EVAL_303;
  assign _EVAL_247 = _EVAL_11 ? _EVAL_278 : _EVAL_245;
endmodule
