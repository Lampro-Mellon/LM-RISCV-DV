//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_183_assert(
  input        _EVAL,
  input        _EVAL_0,
  input        _EVAL_1,
  input  [3:0] _EVAL_24
);
  wire  _EVAL_3;
  wire  _EVAL_6;
  wire  _EVAL_8;
  wire  _EVAL_9;
  wire  _EVAL_10;
  wire  _EVAL_11;
  wire  _EVAL_12;
  wire  _EVAL_14;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_53;
  wire  _EVAL_56;
  wire  _EVAL_58;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_71;
  wire  _EVAL_73;
  wire  _EVAL_76;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_88;
  wire  _EVAL_90;
  wire  _EVAL_92;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_104;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  assign _EVAL_42 = _EVAL_95 & _EVAL_99;
  assign _EVAL_58 = _EVAL_11 & _EVAL;
  assign _EVAL_108 = _EVAL_39 & _EVAL_53;
  assign _EVAL_34 = _EVAL_104 & _EVAL;
  assign _EVAL_110 = _EVAL_102 & _EVAL_53;
  assign _EVAL_68 = _EVAL_84 & _EVAL_53;
  assign _EVAL_84 = _EVAL_24 == 4'h2;
  assign _EVAL_25 = _EVAL_84 & _EVAL;
  assign _EVAL_38 = _EVAL_14 & _EVAL_53;
  assign _EVAL_79 = _EVAL_43 & _EVAL;
  assign _EVAL_17 = _EVAL_36 & _EVAL_53;
  assign _EVAL_50 = _EVAL_112 & _EVAL_99;
  assign _EVAL_90 = _EVAL_39 & _EVAL_99;
  assign _EVAL_35 = _EVAL_71 & _EVAL_99;
  assign _EVAL_12 = _EVAL_43 & _EVAL_99;
  assign _EVAL_3 = _EVAL_109 & _EVAL;
  assign _EVAL_21 = _EVAL_112 & _EVAL;
  assign _EVAL_26 = ~_EVAL_99;
  assign _EVAL_14 = _EVAL_24 == 4'hf;
  assign _EVAL_113 = _EVAL_11 & _EVAL_99;
  assign _EVAL_36 = _EVAL_24 == 4'h3;
  assign _EVAL_102 = _EVAL_24 == 4'h1;
  assign _EVAL_99 = _EVAL_0;
  assign _EVAL_9 = _EVAL_24 == 4'hb;
  assign _EVAL_64 = _EVAL_18 & _EVAL_53;
  assign _EVAL_65 = _EVAL_104 & _EVAL_53;
  assign _EVAL_112 = _EVAL_24 == 4'h5;
  assign _EVAL_69 = _EVAL_111 & _EVAL_53;
  assign _EVAL_39 = _EVAL_24 == 4'h9;
  assign _EVAL_97 = _EVAL_43 & _EVAL_53;
  assign _EVAL_18 = _EVAL_24 == 4'hd;
  assign _EVAL_6 = _EVAL_18 & _EVAL_99;
  assign _EVAL_95 = _EVAL_24 == 4'hc;
  assign _EVAL_73 = _EVAL_36 & _EVAL_99;
  assign _EVAL_19 = _EVAL_71 & _EVAL_53;
  assign _EVAL_8 = _EVAL_9 & _EVAL_99;
  assign _EVAL_85 = _EVAL_102 & _EVAL;
  assign _EVAL_86 = _EVAL_11 & _EVAL_53;
  assign _EVAL_10 = _EVAL_9 & _EVAL_53;
  assign _EVAL_98 = _EVAL_24 == 4'h6;
  assign _EVAL_106 = _EVAL_95 & _EVAL;
  assign _EVAL_78 = _EVAL_98 & _EVAL_53;
  assign _EVAL_96 = _EVAL_84 & _EVAL_99;
  assign _EVAL_20 = _EVAL_112 & _EVAL_53;
  assign _EVAL_63 = _EVAL_111 & _EVAL_99;
  assign _EVAL_82 = _EVAL_102 & _EVAL_99;
  assign _EVAL_101 = _EVAL_104 & _EVAL_99;
  assign _EVAL_107 = _EVAL_9 & _EVAL;
  assign _EVAL_30 = _EVAL_98 & _EVAL_99;
  assign _EVAL_31 = _EVAL_98 & _EVAL;
  assign _EVAL_88 = _EVAL_14 & _EVAL;
  assign _EVAL_92 = _EVAL_18 & _EVAL;
  assign _EVAL_51 = _EVAL_39 & _EVAL;
  assign _EVAL_41 = _EVAL_109 & _EVAL_53;
  assign _EVAL_83 = _EVAL_71 & _EVAL;
  assign _EVAL_71 = _EVAL_24 == 4'ha;
  assign _EVAL_111 = _EVAL_24 == 4'h7;
  assign _EVAL_104 = _EVAL_24 == 4'h8;
  assign _EVAL_49 = _EVAL_95 & _EVAL_53;
  assign _EVAL_56 = _EVAL_36 & _EVAL;
  assign _EVAL_109 = _EVAL_24 == 4'he;
  assign _EVAL_53 = ~_EVAL;
  assign _EVAL_11 = _EVAL_24 == 4'h4;
  assign _EVAL_43 = _EVAL_24 == 4'h0;
  assign _EVAL_76 = _EVAL_109 & _EVAL_99;
  assign _EVAL_29 = _EVAL_111 & _EVAL;
  assign _EVAL_27 = _EVAL_14 & _EVAL_99;
  always @(posedge _EVAL_1) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23209941)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbd14242)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4063409c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9354c8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_10 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cec7298a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(564e0447)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(240b2c8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56d5add3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(762d94a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fd1fc89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95776544)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f34e1981)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72ea99fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19cccdf8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6c7c3d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b1b230c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb95267)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c93f6fcb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54eb487c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa49f817)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d494e55a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6f7736d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8282d629)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61d6fb31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1889f32b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f1bba4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b978e73b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d256f12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c456feb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e84c7f70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a16adac5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_8 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bc134fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5f0a6b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d997b4fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44a67fee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8362fc97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6551f21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2f6e18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0a4a287)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f39bb7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6fec0b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdbf35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af7edd20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a49a7b2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6e8c898)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(397043f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b3d24d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(658e600b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
