//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_104(
  output        _EVAL,
  output        _EVAL_0,
  input         _EVAL_1,
  output        _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [3:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  input  [2:0]  _EVAL_7,
  output [3:0]  _EVAL_8,
  input         _EVAL_9,
  output        _EVAL_10,
  input  [29:0] _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  output [31:0] _EVAL_14,
  output        _EVAL_15,
  input  [2:0]  _EVAL_16,
  output        _EVAL_17,
  input         _EVAL_18,
  output        _EVAL_19,
  output [3:0]  _EVAL_20,
  input         _EVAL_21,
  input         _EVAL_22,
  output [29:0] _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  output        _EVAL_26,
  output [2:0]  _EVAL_27,
  output [2:0]  _EVAL_28,
  output        _EVAL_29,
  output [2:0]  _EVAL_30,
  output        _EVAL_31,
  input         _EVAL_32,
  input  [3:0]  _EVAL_33,
  input  [31:0] _EVAL_34
);
  reg  _EVAL_35 [0:0];
  reg [31:0] _RAND_0;
  wire  _EVAL_35__EVAL_36_data;
  wire  _EVAL_35__EVAL_36_addr;
  wire  _EVAL_35__EVAL_37_data;
  wire  _EVAL_35__EVAL_37_addr;
  wire  _EVAL_35__EVAL_37_mask;
  wire  _EVAL_35__EVAL_37_en;
  reg [3:0] _EVAL_38 [0:0];
  reg [31:0] _RAND_1;
  wire [3:0] _EVAL_38__EVAL_39_data;
  wire  _EVAL_38__EVAL_39_addr;
  wire [3:0] _EVAL_38__EVAL_40_data;
  wire  _EVAL_38__EVAL_40_addr;
  wire  _EVAL_38__EVAL_40_mask;
  wire  _EVAL_38__EVAL_40_en;
  wire  _EVAL_41;
  reg  _EVAL_42 [0:0];
  reg [31:0] _RAND_2;
  wire  _EVAL_42__EVAL_43_data;
  wire  _EVAL_42__EVAL_43_addr;
  wire  _EVAL_42__EVAL_44_data;
  wire  _EVAL_42__EVAL_44_addr;
  wire  _EVAL_42__EVAL_44_mask;
  wire  _EVAL_42__EVAL_44_en;
  reg  _EVAL_45 [0:0];
  reg [31:0] _RAND_3;
  wire  _EVAL_45__EVAL_46_data;
  wire  _EVAL_45__EVAL_46_addr;
  wire  _EVAL_45__EVAL_47_data;
  wire  _EVAL_45__EVAL_47_addr;
  wire  _EVAL_45__EVAL_47_mask;
  wire  _EVAL_45__EVAL_47_en;
  reg  _EVAL_49 [0:0];
  reg [31:0] _RAND_4;
  wire  _EVAL_49__EVAL_50_data;
  wire  _EVAL_49__EVAL_50_addr;
  wire  _EVAL_49__EVAL_51_data;
  wire  _EVAL_49__EVAL_51_addr;
  wire  _EVAL_49__EVAL_51_mask;
  wire  _EVAL_49__EVAL_51_en;
  reg  _EVAL_52 [0:0];
  reg [31:0] _RAND_5;
  wire  _EVAL_52__EVAL_53_data;
  wire  _EVAL_52__EVAL_53_addr;
  wire  _EVAL_52__EVAL_54_data;
  wire  _EVAL_52__EVAL_54_addr;
  wire  _EVAL_52__EVAL_54_mask;
  wire  _EVAL_52__EVAL_54_en;
  wire  _EVAL_55;
  wire  _EVAL_56;
  reg [29:0] _EVAL_57 [0:0];
  reg [31:0] _RAND_6;
  wire [29:0] _EVAL_57__EVAL_58_data;
  wire  _EVAL_57__EVAL_58_addr;
  wire [29:0] _EVAL_57__EVAL_59_data;
  wire  _EVAL_57__EVAL_59_addr;
  wire  _EVAL_57__EVAL_59_mask;
  wire  _EVAL_57__EVAL_59_en;
  reg  _EVAL_60 [0:0];
  reg [31:0] _RAND_7;
  wire  _EVAL_60__EVAL_61_data;
  wire  _EVAL_60__EVAL_61_addr;
  wire  _EVAL_60__EVAL_62_data;
  wire  _EVAL_60__EVAL_62_addr;
  wire  _EVAL_60__EVAL_62_mask;
  wire  _EVAL_60__EVAL_62_en;
  reg [2:0] _EVAL_63 [0:0];
  reg [31:0] _RAND_8;
  wire [2:0] _EVAL_63__EVAL_64_data;
  wire  _EVAL_63__EVAL_64_addr;
  wire [2:0] _EVAL_63__EVAL_65_data;
  wire  _EVAL_63__EVAL_65_addr;
  wire  _EVAL_63__EVAL_65_mask;
  wire  _EVAL_63__EVAL_65_en;
  reg  _EVAL_66;
  reg [31:0] _RAND_9;
  reg  _EVAL_67 [0:0];
  reg [31:0] _RAND_10;
  wire  _EVAL_67__EVAL_68_data;
  wire  _EVAL_67__EVAL_68_addr;
  wire  _EVAL_67__EVAL_69_data;
  wire  _EVAL_67__EVAL_69_addr;
  wire  _EVAL_67__EVAL_69_mask;
  wire  _EVAL_67__EVAL_69_en;
  reg [31:0] _EVAL_70 [0:0];
  reg [31:0] _RAND_11;
  wire [31:0] _EVAL_70__EVAL_71_data;
  wire  _EVAL_70__EVAL_71_addr;
  wire [31:0] _EVAL_70__EVAL_72_data;
  wire  _EVAL_70__EVAL_72_addr;
  wire  _EVAL_70__EVAL_72_mask;
  wire  _EVAL_70__EVAL_72_en;
  reg [3:0] _EVAL_73 [0:0];
  reg [31:0] _RAND_12;
  wire [3:0] _EVAL_73__EVAL_74_data;
  wire  _EVAL_73__EVAL_74_addr;
  wire [3:0] _EVAL_73__EVAL_75_data;
  wire  _EVAL_73__EVAL_75_addr;
  wire  _EVAL_73__EVAL_75_mask;
  wire  _EVAL_73__EVAL_75_en;
  reg [2:0] _EVAL_76 [0:0];
  reg [31:0] _RAND_13;
  wire [2:0] _EVAL_76__EVAL_77_data;
  wire  _EVAL_76__EVAL_77_addr;
  wire [2:0] _EVAL_76__EVAL_78_data;
  wire  _EVAL_76__EVAL_78_addr;
  wire  _EVAL_76__EVAL_78_mask;
  wire  _EVAL_76__EVAL_78_en;
  reg [2:0] _EVAL_79 [0:0];
  reg [31:0] _RAND_14;
  wire [2:0] _EVAL_79__EVAL_80_data;
  wire  _EVAL_79__EVAL_80_addr;
  wire [2:0] _EVAL_79__EVAL_81_data;
  wire  _EVAL_79__EVAL_81_addr;
  wire  _EVAL_79__EVAL_81_mask;
  wire  _EVAL_79__EVAL_81_en;
  wire  _EVAL_82;
  reg  _EVAL_83 [0:0];
  reg [31:0] _RAND_15;
  wire  _EVAL_83__EVAL_84_data;
  wire  _EVAL_83__EVAL_84_addr;
  wire  _EVAL_83__EVAL_85_data;
  wire  _EVAL_83__EVAL_85_addr;
  wire  _EVAL_83__EVAL_85_mask;
  wire  _EVAL_83__EVAL_85_en;
  assign _EVAL_35__EVAL_36_addr = 1'h0;
  assign _EVAL_35__EVAL_36_data = _EVAL_35[_EVAL_35__EVAL_36_addr];
  assign _EVAL_35__EVAL_37_data = _EVAL_21;
  assign _EVAL_35__EVAL_37_addr = 1'h0;
  assign _EVAL_35__EVAL_37_mask = 1'h1;
  assign _EVAL_35__EVAL_37_en = _EVAL_17 & _EVAL_22;
  assign _EVAL_38__EVAL_39_addr = 1'h0;
  assign _EVAL_38__EVAL_39_data = _EVAL_38[_EVAL_38__EVAL_39_addr];
  assign _EVAL_38__EVAL_40_data = _EVAL_33;
  assign _EVAL_38__EVAL_40_addr = 1'h0;
  assign _EVAL_38__EVAL_40_mask = 1'h1;
  assign _EVAL_38__EVAL_40_en = _EVAL_17 & _EVAL_22;
  assign _EVAL_42__EVAL_43_addr = 1'h0;
  assign _EVAL_42__EVAL_43_data = _EVAL_42[_EVAL_42__EVAL_43_addr];
  assign _EVAL_42__EVAL_44_data = _EVAL_1;
  assign _EVAL_42__EVAL_44_addr = 1'h0;
  assign _EVAL_42__EVAL_44_mask = 1'h1;
  assign _EVAL_42__EVAL_44_en = _EVAL_17 & _EVAL_22;
  assign _EVAL_45__EVAL_46_addr = 1'h0;
  assign _EVAL_45__EVAL_46_data = _EVAL_45[_EVAL_45__EVAL_46_addr];
  assign _EVAL_45__EVAL_47_data = _EVAL_32;
  assign _EVAL_45__EVAL_47_addr = 1'h0;
  assign _EVAL_45__EVAL_47_mask = 1'h1;
  assign _EVAL_45__EVAL_47_en = _EVAL_17 & _EVAL_22;
  assign _EVAL_49__EVAL_50_addr = 1'h0;
  assign _EVAL_49__EVAL_50_data = _EVAL_49[_EVAL_49__EVAL_50_addr];
  assign _EVAL_49__EVAL_51_data = _EVAL_13;
  assign _EVAL_49__EVAL_51_addr = 1'h0;
  assign _EVAL_49__EVAL_51_mask = 1'h1;
  assign _EVAL_49__EVAL_51_en = _EVAL_17 & _EVAL_22;
  assign _EVAL_52__EVAL_53_addr = 1'h0;
  assign _EVAL_52__EVAL_53_data = _EVAL_52[_EVAL_52__EVAL_53_addr];
  assign _EVAL_52__EVAL_54_data = _EVAL_3;
  assign _EVAL_52__EVAL_54_addr = 1'h0;
  assign _EVAL_52__EVAL_54_mask = 1'h1;
  assign _EVAL_52__EVAL_54_en = _EVAL_17 & _EVAL_22;
  assign _EVAL_57__EVAL_58_addr = 1'h0;
  assign _EVAL_57__EVAL_58_data = _EVAL_57[_EVAL_57__EVAL_58_addr];
  assign _EVAL_57__EVAL_59_data = _EVAL_11;
  assign _EVAL_57__EVAL_59_addr = 1'h0;
  assign _EVAL_57__EVAL_59_mask = 1'h1;
  assign _EVAL_57__EVAL_59_en = _EVAL_17 & _EVAL_22;
  assign _EVAL_60__EVAL_61_addr = 1'h0;
  assign _EVAL_60__EVAL_61_data = _EVAL_60[_EVAL_60__EVAL_61_addr];
  assign _EVAL_60__EVAL_62_data = _EVAL_9;
  assign _EVAL_60__EVAL_62_addr = 1'h0;
  assign _EVAL_60__EVAL_62_mask = 1'h1;
  assign _EVAL_60__EVAL_62_en = _EVAL_17 & _EVAL_22;
  assign _EVAL_63__EVAL_64_addr = 1'h0;
  assign _EVAL_63__EVAL_64_data = _EVAL_63[_EVAL_63__EVAL_64_addr];
  assign _EVAL_63__EVAL_65_data = _EVAL_6;
  assign _EVAL_63__EVAL_65_addr = 1'h0;
  assign _EVAL_63__EVAL_65_mask = 1'h1;
  assign _EVAL_63__EVAL_65_en = _EVAL_17 & _EVAL_22;
  assign _EVAL_67__EVAL_68_addr = 1'h0;
  assign _EVAL_67__EVAL_68_data = _EVAL_67[_EVAL_67__EVAL_68_addr];
  assign _EVAL_67__EVAL_69_data = _EVAL_12;
  assign _EVAL_67__EVAL_69_addr = 1'h0;
  assign _EVAL_67__EVAL_69_mask = 1'h1;
  assign _EVAL_67__EVAL_69_en = _EVAL_17 & _EVAL_22;
  assign _EVAL_70__EVAL_71_addr = 1'h0;
  assign _EVAL_70__EVAL_71_data = _EVAL_70[_EVAL_70__EVAL_71_addr];
  assign _EVAL_70__EVAL_72_data = _EVAL_34;
  assign _EVAL_70__EVAL_72_addr = 1'h0;
  assign _EVAL_70__EVAL_72_mask = 1'h1;
  assign _EVAL_70__EVAL_72_en = _EVAL_17 & _EVAL_22;
  assign _EVAL_73__EVAL_74_addr = 1'h0;
  assign _EVAL_73__EVAL_74_data = _EVAL_73[_EVAL_73__EVAL_74_addr];
  assign _EVAL_73__EVAL_75_data = _EVAL_5;
  assign _EVAL_73__EVAL_75_addr = 1'h0;
  assign _EVAL_73__EVAL_75_mask = 1'h1;
  assign _EVAL_73__EVAL_75_en = _EVAL_17 & _EVAL_22;
  assign _EVAL_76__EVAL_77_addr = 1'h0;
  assign _EVAL_76__EVAL_77_data = _EVAL_76[_EVAL_76__EVAL_77_addr];
  assign _EVAL_76__EVAL_78_data = _EVAL_7;
  assign _EVAL_76__EVAL_78_addr = 1'h0;
  assign _EVAL_76__EVAL_78_mask = 1'h1;
  assign _EVAL_76__EVAL_78_en = _EVAL_17 & _EVAL_22;
  assign _EVAL_79__EVAL_80_addr = 1'h0;
  assign _EVAL_79__EVAL_80_data = _EVAL_79[_EVAL_79__EVAL_80_addr];
  assign _EVAL_79__EVAL_81_data = _EVAL_16;
  assign _EVAL_79__EVAL_81_addr = 1'h0;
  assign _EVAL_79__EVAL_81_mask = 1'h1;
  assign _EVAL_79__EVAL_81_en = _EVAL_17 & _EVAL_22;
  assign _EVAL_83__EVAL_84_addr = 1'h0;
  assign _EVAL_83__EVAL_84_data = _EVAL_83[_EVAL_83__EVAL_84_addr];
  assign _EVAL_83__EVAL_85_data = _EVAL_25;
  assign _EVAL_83__EVAL_85_addr = 1'h0;
  assign _EVAL_83__EVAL_85_mask = 1'h1;
  assign _EVAL_83__EVAL_85_en = _EVAL_17 & _EVAL_22;
  assign _EVAL_56 = ~_EVAL_66;
  assign _EVAL_82 = _EVAL_24 & _EVAL_31;
  assign _EVAL = _EVAL_42__EVAL_43_data;
  assign _EVAL_20 = _EVAL_73__EVAL_74_data;
  assign _EVAL_14 = _EVAL_70__EVAL_71_data;
  assign _EVAL_15 = _EVAL_83__EVAL_84_data;
  assign _EVAL_23 = _EVAL_57__EVAL_58_data;
  assign _EVAL_17 = _EVAL_24 | _EVAL_56;
  assign _EVAL_8 = _EVAL_38__EVAL_39_data;
  assign _EVAL_28 = _EVAL_63__EVAL_64_data;
  assign _EVAL_41 = _EVAL_17 & _EVAL_22;
  assign _EVAL_55 = _EVAL_41 != _EVAL_82;
  assign _EVAL_29 = _EVAL_45__EVAL_46_data;
  assign _EVAL_27 = _EVAL_79__EVAL_80_data;
  assign _EVAL_10 = _EVAL_52__EVAL_53_data;
  assign _EVAL_26 = _EVAL_49__EVAL_50_data;
  assign _EVAL_2 = _EVAL_35__EVAL_36_data;
  assign _EVAL_30 = _EVAL_76__EVAL_77_data;
  assign _EVAL_31 = ~_EVAL_56;
  assign _EVAL_0 = _EVAL_60__EVAL_61_data;
  assign _EVAL_19 = _EVAL_67__EVAL_68_data;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_35[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_38[initvar] = _RAND_1[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_42[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_45[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_49[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_52[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_57[initvar] = _RAND_6[29:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_60[initvar] = _RAND_7[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_63[initvar] = _RAND_8[2:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_66 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_67[initvar] = _RAND_10[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_11 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_70[initvar] = _RAND_11[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_73[initvar] = _RAND_12[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_13 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_76[initvar] = _RAND_13[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_14 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_79[initvar] = _RAND_14[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_15 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_83[initvar] = _RAND_15[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_18) begin
    if(_EVAL_35__EVAL_37_en & _EVAL_35__EVAL_37_mask) begin
      _EVAL_35[_EVAL_35__EVAL_37_addr] <= _EVAL_35__EVAL_37_data;
    end
    if(_EVAL_38__EVAL_40_en & _EVAL_38__EVAL_40_mask) begin
      _EVAL_38[_EVAL_38__EVAL_40_addr] <= _EVAL_38__EVAL_40_data;
    end
    if(_EVAL_42__EVAL_44_en & _EVAL_42__EVAL_44_mask) begin
      _EVAL_42[_EVAL_42__EVAL_44_addr] <= _EVAL_42__EVAL_44_data;
    end
    if(_EVAL_45__EVAL_47_en & _EVAL_45__EVAL_47_mask) begin
      _EVAL_45[_EVAL_45__EVAL_47_addr] <= _EVAL_45__EVAL_47_data;
    end
    if(_EVAL_49__EVAL_51_en & _EVAL_49__EVAL_51_mask) begin
      _EVAL_49[_EVAL_49__EVAL_51_addr] <= _EVAL_49__EVAL_51_data;
    end
    if(_EVAL_52__EVAL_54_en & _EVAL_52__EVAL_54_mask) begin
      _EVAL_52[_EVAL_52__EVAL_54_addr] <= _EVAL_52__EVAL_54_data;
    end
    if(_EVAL_57__EVAL_59_en & _EVAL_57__EVAL_59_mask) begin
      _EVAL_57[_EVAL_57__EVAL_59_addr] <= _EVAL_57__EVAL_59_data;
    end
    if(_EVAL_60__EVAL_62_en & _EVAL_60__EVAL_62_mask) begin
      _EVAL_60[_EVAL_60__EVAL_62_addr] <= _EVAL_60__EVAL_62_data;
    end
    if(_EVAL_63__EVAL_65_en & _EVAL_63__EVAL_65_mask) begin
      _EVAL_63[_EVAL_63__EVAL_65_addr] <= _EVAL_63__EVAL_65_data;
    end
    if (_EVAL_4) begin
      _EVAL_66 <= 1'h0;
    end else if (_EVAL_55) begin
      _EVAL_66 <= _EVAL_41;
    end
    if(_EVAL_67__EVAL_69_en & _EVAL_67__EVAL_69_mask) begin
      _EVAL_67[_EVAL_67__EVAL_69_addr] <= _EVAL_67__EVAL_69_data;
    end
    if(_EVAL_70__EVAL_72_en & _EVAL_70__EVAL_72_mask) begin
      _EVAL_70[_EVAL_70__EVAL_72_addr] <= _EVAL_70__EVAL_72_data;
    end
    if(_EVAL_73__EVAL_75_en & _EVAL_73__EVAL_75_mask) begin
      _EVAL_73[_EVAL_73__EVAL_75_addr] <= _EVAL_73__EVAL_75_data;
    end
    if(_EVAL_76__EVAL_78_en & _EVAL_76__EVAL_78_mask) begin
      _EVAL_76[_EVAL_76__EVAL_78_addr] <= _EVAL_76__EVAL_78_data;
    end
    if(_EVAL_79__EVAL_81_en & _EVAL_79__EVAL_81_mask) begin
      _EVAL_79[_EVAL_79__EVAL_81_addr] <= _EVAL_79__EVAL_81_data;
    end
    if(_EVAL_83__EVAL_85_en & _EVAL_83__EVAL_85_mask) begin
      _EVAL_83[_EVAL_83__EVAL_85_addr] <= _EVAL_83__EVAL_85_data;
    end
  end
endmodule
