//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_127(
  input         _EVAL,
  output [3:0]  _EVAL_0,
  output [2:0]  _EVAL_1,
  output [2:0]  _EVAL_2,
  input  [1:0]  _EVAL_3,
  output        _EVAL_4,
  input  [1:0]  _EVAL_5,
  output        _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  output        _EVAL_10,
  output [1:0]  _EVAL_11,
  output [31:0] _EVAL_12,
  output [31:0] _EVAL_13,
  input  [2:0]  _EVAL_14,
  output        _EVAL_15,
  input  [2:0]  _EVAL_16,
  input  [31:0] _EVAL_17,
  input  [8:0]  _EVAL_18,
  input  [31:0] _EVAL_19,
  output        _EVAL_20,
  output        _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  input         _EVAL_26,
  output [1:0]  _EVAL_27,
  output        _EVAL_28,
  input         _EVAL_29,
  input  [3:0]  _EVAL_30,
  output [8:0]  _EVAL_31,
  input         _EVAL_32,
  output        _EVAL_33
);
  wire  error__EVAL;
  wire  error__EVAL_0;
  wire  error__EVAL_1;
  wire  error__EVAL_2;
  wire [2:0] error__EVAL_3;
  wire [31:0] error__EVAL_4;
  wire  error__EVAL_5;
  wire [3:0] error__EVAL_6;
  wire  error__EVAL_7;
  wire  error__EVAL_8;
  wire [1:0] error__EVAL_9;
  wire [1:0] error__EVAL_10;
  wire  error__EVAL_11;
  wire [2:0] error__EVAL_12;
  wire  error__EVAL_13;
  wire  error__EVAL_14;
  wire [127:0] error__EVAL_15;
  wire  bar__EVAL;
  wire [31:0] bar__EVAL_0;
  wire [1:0] bar__EVAL_1;
  wire  bar__EVAL_2;
  wire [31:0] bar__EVAL_3;
  wire  bar__EVAL_4;
  wire [31:0] bar__EVAL_5;
  wire [2:0] bar__EVAL_6;
  wire [2:0] bar__EVAL_7;
  wire [2:0] bar__EVAL_8;
  wire  bar__EVAL_9;
  wire [8:0] bar__EVAL_10;
  wire [3:0] bar__EVAL_11;
  wire  bar__EVAL_12;
  wire  bar__EVAL_13;
  wire  bar__EVAL_14;
  wire  bar__EVAL_15;
  wire [3:0] bar__EVAL_16;
  wire [31:0] bar__EVAL_17;
  wire  bar__EVAL_18;
  wire [1:0] bar__EVAL_19;
  wire  bar__EVAL_20;
  wire  bar__EVAL_21;
  wire  bar__EVAL_22;
  wire [1:0] bar__EVAL_23;
  wire [2:0] bar__EVAL_24;
  wire [31:0] bar__EVAL_25;
  wire [8:0] bar__EVAL_26;
  wire [2:0] bar__EVAL_27;
  wire  bar__EVAL_28;
  wire [1:0] bar__EVAL_29;
  wire  bar__EVAL_30;
  wire [1:0] bar__EVAL_31;
  wire  bar__EVAL_32;
  wire [1:0] bar__EVAL_33;
  wire [3:0] bar__EVAL_34;
  wire  bar__EVAL_35;
  wire  bar__EVAL_36;
  wire  bar__EVAL_37;
  wire [2:0] bar__EVAL_38;
  wire  bar__EVAL_39;
  wire [127:0] bar__EVAL_40;
  wire  bar__EVAL_41;
  wire  bar__EVAL_42;
  wire  bar__EVAL_43;
  wire  bar__EVAL_44;
  wire  bar__EVAL_45;
  wire  bar__EVAL_46;
  wire  bar__EVAL_47;
  wire  bar__EVAL_48;
  _EVAL_126 error (
    ._EVAL(error__EVAL),
    ._EVAL_0(error__EVAL_0),
    ._EVAL_1(error__EVAL_1),
    ._EVAL_2(error__EVAL_2),
    ._EVAL_3(error__EVAL_3),
    ._EVAL_4(error__EVAL_4),
    ._EVAL_5(error__EVAL_5),
    ._EVAL_6(error__EVAL_6),
    ._EVAL_7(error__EVAL_7),
    ._EVAL_8(error__EVAL_8),
    ._EVAL_9(error__EVAL_9),
    ._EVAL_10(error__EVAL_10),
    ._EVAL_11(error__EVAL_11),
    ._EVAL_12(error__EVAL_12),
    ._EVAL_13(error__EVAL_13),
    ._EVAL_14(error__EVAL_14),
    ._EVAL_15(error__EVAL_15)
  );
  _EVAL_124 bar (
    ._EVAL(bar__EVAL),
    ._EVAL_0(bar__EVAL_0),
    ._EVAL_1(bar__EVAL_1),
    ._EVAL_2(bar__EVAL_2),
    ._EVAL_3(bar__EVAL_3),
    ._EVAL_4(bar__EVAL_4),
    ._EVAL_5(bar__EVAL_5),
    ._EVAL_6(bar__EVAL_6),
    ._EVAL_7(bar__EVAL_7),
    ._EVAL_8(bar__EVAL_8),
    ._EVAL_9(bar__EVAL_9),
    ._EVAL_10(bar__EVAL_10),
    ._EVAL_11(bar__EVAL_11),
    ._EVAL_12(bar__EVAL_12),
    ._EVAL_13(bar__EVAL_13),
    ._EVAL_14(bar__EVAL_14),
    ._EVAL_15(bar__EVAL_15),
    ._EVAL_16(bar__EVAL_16),
    ._EVAL_17(bar__EVAL_17),
    ._EVAL_18(bar__EVAL_18),
    ._EVAL_19(bar__EVAL_19),
    ._EVAL_20(bar__EVAL_20),
    ._EVAL_21(bar__EVAL_21),
    ._EVAL_22(bar__EVAL_22),
    ._EVAL_23(bar__EVAL_23),
    ._EVAL_24(bar__EVAL_24),
    ._EVAL_25(bar__EVAL_25),
    ._EVAL_26(bar__EVAL_26),
    ._EVAL_27(bar__EVAL_27),
    ._EVAL_28(bar__EVAL_28),
    ._EVAL_29(bar__EVAL_29),
    ._EVAL_30(bar__EVAL_30),
    ._EVAL_31(bar__EVAL_31),
    ._EVAL_32(bar__EVAL_32),
    ._EVAL_33(bar__EVAL_33),
    ._EVAL_34(bar__EVAL_34),
    ._EVAL_35(bar__EVAL_35),
    ._EVAL_36(bar__EVAL_36),
    ._EVAL_37(bar__EVAL_37),
    ._EVAL_38(bar__EVAL_38),
    ._EVAL_39(bar__EVAL_39),
    ._EVAL_40(bar__EVAL_40),
    ._EVAL_41(bar__EVAL_41),
    ._EVAL_42(bar__EVAL_42),
    ._EVAL_43(bar__EVAL_43),
    ._EVAL_44(bar__EVAL_44),
    ._EVAL_45(bar__EVAL_45),
    ._EVAL_46(bar__EVAL_46),
    ._EVAL_47(bar__EVAL_47),
    ._EVAL_48(bar__EVAL_48)
  );
  assign bar__EVAL_8 = _EVAL_16;
  assign error__EVAL_5 = _EVAL;
  assign bar__EVAL = _EVAL_7;
  assign _EVAL_1 = bar__EVAL_38;
  assign bar__EVAL_24 = _EVAL_14;
  assign bar__EVAL_47 = _EVAL_8;
  assign _EVAL_11 = bar__EVAL_33;
  assign bar__EVAL_35 = _EVAL_25;
  assign bar__EVAL_23 = error__EVAL_10;
  assign bar__EVAL_28 = error__EVAL_7;
  assign error__EVAL_14 = bar__EVAL_4;
  assign bar__EVAL_48 = _EVAL_26;
  assign error__EVAL_15 = bar__EVAL_40;
  assign bar__EVAL_3 = error__EVAL_4;
  assign error__EVAL_11 = _EVAL_22;
  assign bar__EVAL_18 = error__EVAL_13;
  assign bar__EVAL_37 = error__EVAL_8;
  assign bar__EVAL_42 = _EVAL_32;
  assign bar__EVAL_31 = _EVAL_5;
  assign _EVAL_27 = bar__EVAL_1;
  assign bar__EVAL_12 = _EVAL;
  assign _EVAL_0 = bar__EVAL_11;
  assign _EVAL_20 = bar__EVAL_44;
  assign bar__EVAL_32 = error__EVAL_2;
  assign _EVAL_2 = bar__EVAL_6;
  assign bar__EVAL_41 = _EVAL_24;
  assign _EVAL_15 = bar__EVAL_2;
  assign bar__EVAL_16 = _EVAL_30;
  assign bar__EVAL_15 = _EVAL_9;
  assign bar__EVAL_26 = _EVAL_18;
  assign error__EVAL_6 = bar__EVAL_34;
  assign bar__EVAL_22 = _EVAL_23;
  assign _EVAL_4 = bar__EVAL_39;
  assign error__EVAL_0 = bar__EVAL_45;
  assign _EVAL_33 = bar__EVAL_36;
  assign error__EVAL_12 = bar__EVAL_27;
  assign bar__EVAL_29 = _EVAL_3;
  assign bar__EVAL_7 = error__EVAL_3;
  assign bar__EVAL_25 = _EVAL_19;
  assign _EVAL_31 = bar__EVAL_10;
  assign bar__EVAL_21 = error__EVAL;
  assign _EVAL_12 = bar__EVAL_17;
  assign _EVAL_28 = bar__EVAL_46;
  assign bar__EVAL_5 = _EVAL_17;
  assign bar__EVAL_13 = _EVAL_22;
  assign _EVAL_21 = bar__EVAL_9;
  assign _EVAL_6 = bar__EVAL_30;
  assign bar__EVAL_43 = error__EVAL_1;
  assign _EVAL_13 = bar__EVAL_0;
  assign bar__EVAL_20 = _EVAL_29;
  assign _EVAL_10 = bar__EVAL_14;
  assign bar__EVAL_19 = error__EVAL_9;
endmodule
