//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module CoreIPSubsystemAllPortRAMTestHarness(
  input   clock,
  input   reset,
  output  io_success
);
  wire  system_clock;
  wire  system_reset;
  wire  system_halt_from_tile_0;
  wire  system_wfi_from_tile_0;
  wire  system_cease_from_tile_0;
  wire  system_psd_test_clock_enable;
  wire  system_meip_0;
  wire  system_resetctrl_hartIsInReset_0;
  wire  system_debug_clock;
  wire  system_debug_reset;
  wire  system_debug_systemjtag_jtag_TCK;
  wire  system_debug_systemjtag_jtag_TMS;
  wire  system_debug_systemjtag_jtag_TDI;
  wire  system_debug_systemjtag_jtag_TDO_data;
  wire  system_debug_systemjtag_jtag_TDO_driven;
  wire  system_debug_systemjtag_reset;
  wire [10:0] system_debug_systemjtag_mfr_id;
  wire [15:0] system_debug_systemjtag_part_number;
  wire [3:0] system_debug_systemjtag_version;
  wire  system_debug_ndreset;
  wire  system_debug_dmactive;
  wire  system_debug_dmactiveAck;
  wire [31:0] system_reset_vector_0;
  wire  system_rtc_toggle;
  wire [126:0] system_local_interrupts_0;
  wire  system_sys_port_ahb_0_hmastlock;
  wire  system_sys_port_ahb_0_hready;
  wire [1:0] system_sys_port_ahb_0_htrans;
  wire [2:0] system_sys_port_ahb_0_hsize;
  wire [2:0] system_sys_port_ahb_0_hburst;
  wire  system_sys_port_ahb_0_hwrite;
  wire [3:0] system_sys_port_ahb_0_hprot;
  wire [30:0] system_sys_port_ahb_0_haddr;
  wire [31:0] system_sys_port_ahb_0_hwdata;
  wire  system_sys_port_ahb_0_hresp;
  wire [31:0] system_sys_port_ahb_0_hrdata;
  wire  system_periph_port_ahb_0_hmastlock;
  wire  system_periph_port_ahb_0_hready;
  wire [1:0] system_periph_port_ahb_0_htrans;
  wire [2:0] system_periph_port_ahb_0_hsize;
  wire [2:0] system_periph_port_ahb_0_hburst;
  wire  system_periph_port_ahb_0_hwrite;
  wire [3:0] system_periph_port_ahb_0_hprot;
  wire [29:0] system_periph_port_ahb_0_haddr;
  wire [31:0] system_periph_port_ahb_0_hwdata;
  wire  system_periph_port_ahb_0_hresp;
  wire [31:0] system_periph_port_ahb_0_hrdata;
  wire  system_front_port_ahb_0_hmastlock;
  wire  system_front_port_ahb_0_hsel;
  wire  system_front_port_ahb_0_hready;
  wire  system_front_port_ahb_0_hreadyout;
  wire [1:0] system_front_port_ahb_0_htrans;
  wire [2:0] system_front_port_ahb_0_hsize;
  wire [2:0] system_front_port_ahb_0_hburst;
  wire  system_front_port_ahb_0_hwrite;
  wire [3:0] system_front_port_ahb_0_hprot;
  wire [31:0] system_front_port_ahb_0_haddr;
  wire [31:0] system_front_port_ahb_0_hwdata;
  wire  system_front_port_ahb_0_hresp;
  wire [31:0] system_front_port_ahb_0_hrdata;
  wire  func_clock_clock;
  wire  func_clock_io_clock_out;
  wire  dpiClockGate_clock_in;
  wire  dpiClockGate_clock_out;
  wire  c_core_reset_driver_clock;
  wire  debug_compatibility_clock;
  wire  debug_compatibility_reset;
  wire  debug_compatibility_debug_outer_reset;
  wire  debug_compatibility_debug_clock;
  wire  debug_compatibility_debug_reset;
  wire  debug_compatibility_debug_dmactive;
  wire  debug_compatibility_debug_dmactiveAck;
  wire  debug_compatibility_debug_resetctrl_hartIsInReset_0;
  wire  DataTap_9__0_clock;
  wire  DataTap_9__0_reset;
  wire  DataTap_9__0_excpt;
  wire [2:0] DataTap_9__0_priv_mode;
  wire [31:0] DataTap_9__0_hartid;
  wire [31:0] DataTap_9__0_timer;
  wire  DataTap_9__0_valid;
  wire [31:0] DataTap_9__0_pc;
  wire [4:0] DataTap_9__0_wrdst;
  wire [31:0] DataTap_9__0_wrdata;
  wire  DataTap_9__0_wrenx;
  wire  DataTap_9__0_wrenf;
  wire [4:0] DataTap_9__0_rd0src;
  wire [31:0] DataTap_9__0_rd0val;
  wire [4:0] DataTap_9__0_rd1src;
  wire [31:0] DataTap_9__0_rd1val;
  wire [31:0] DataTap_9__0_inst;
  wire  DataTap_2__10;
  wire  DataTap_2__9;
  wire  DataTap_2__8;
  wire [7:0] DataTap_2__7;
  wire  DataTap_2__6;
  wire  DataTap_2__5;
  wire [31:0] DataTap_2__4;
  wire [31:0] DataTap_2__3;
  wire [31:0] DataTap_2__2;
  wire [142:0] DataTap_2__1;
  wire [15:0] DataTap_2__0;
  wire  testRAM_clock;
  wire  testRAM_reset;
  wire  testRAM_io_ahb_0_hready;
  wire [1:0] testRAM_io_ahb_0_htrans;
  wire [2:0] testRAM_io_ahb_0_hsize;
  wire  testRAM_io_ahb_0_hwrite;
  wire [29:0] testRAM_io_ahb_0_haddr;
  wire [31:0] testRAM_io_ahb_0_hwdata;
  wire  testRAM_io_ahb_0_hresp;
  wire [31:0] testRAM_io_ahb_0_hrdata;
  wire  testRAM_1_clock;
  wire  testRAM_1_reset;
  wire  testRAM_1_io_ahb_0_hready;
  wire [1:0] testRAM_1_io_ahb_0_htrans;
  wire [2:0] testRAM_1_io_ahb_0_hsize;
  wire  testRAM_1_io_ahb_0_hwrite;
  wire [30:0] testRAM_1_io_ahb_0_haddr;
  wire [31:0] testRAM_1_io_ahb_0_hwdata;
  wire  testRAM_1_io_ahb_0_hresp;
  wire [31:0] testRAM_1_io_ahb_0_hrdata;
  wire  WfiChecker_reset;
  wire  WfiChecker_clock;
  wire  WfiChecker_wfi;
  wire  WfiChecker_excpt;
  wire  WfiChecker_bus_err_int;
  wire  WfiChecker_debug_int;
  wire  WfiChecker_clint_int;
  wire  WfiChecker_allow_wfi;
  wire  WfiChecker_debug;
  wire  WfiChecker_singleStep;
  wire [31:0] WfiChecker_reg_mie;
  wire [31:0] WfiChecker_reg_mip;
  wire  WfiChecker_inst_vld_0;
  wire [31:0] WfiChecker_pc_0;
  wire [31:0] WfiChecker_inst_0;
  wire  core_monitor_m_0_clock;
  wire  core_monitor_m_0_reset;
  wire  core_monitor_m_0_excpt;
  wire [2:0] core_monitor_m_0_priv_mode;
  wire [31:0] core_monitor_m_0_hartid;
  wire [31:0] core_monitor_m_0_timer;
  wire  core_monitor_m_0_valid;
  wire [31:0] core_monitor_m_0_pc;
  wire [4:0] core_monitor_m_0_wrdst;
  wire [31:0] core_monitor_m_0_wrdata;
  wire  core_monitor_m_0_wrenx;
  wire  core_monitor_m_0_wrenf;
  wire [4:0] core_monitor_m_0_rd0src;
  wire [31:0] core_monitor_m_0_rd0val;
  wire [4:0] core_monitor_m_0_rd1src;
  wire [31:0] core_monitor_m_0_rd1val;
  wire [31:0] core_monitor_m_0_inst;
  wire  dpitbh_clock;
  wire  dpitbh_reset;
  wire [31:0] plusarg_reader_out;
  wire  GlobalIntDriver_clock;
  wire  GlobalIntDriver_reset;
  wire [31:0] plusarg_reader_1_out;
  wire  NullInterruptDriver_clock;
  wire  NullInterruptDriver_reset;
  wire [126:0] NullInterruptDriver_interrupts;
  reg [4:0] _T_2;
  reg [31:0] _RAND_0;
  reg  _T_3;
  reg [31:0] _RAND_1;
  wire [4:0] _T_5;
  wire  _T_6;
  wire  _T_7;
  wire  _T_13;
  wire [31:0] _T_30;
  wire  _T_34;
  wire  _T_35;
  wire  _T_36;
  wire  _T_37;
  wire  _T_38;
  wire  _T_41;
  reg [6:0] value_1;
  reg [31:0] _RAND_2;
  wire  _T_43;
  wire [6:0] _T_45;
  wire [31:0] _T_42;
  wire  _T_46;
  wire  _T_47;
  wire  _T_49;
  wire  _T_177;
  reg [6:0] value_2;
  reg [31:0] _RAND_3;
  wire  _T_179;
  wire [6:0] _T_181;
  wire [127:0] _T_182;
  wire  _T_183;
  reg [15:0] _T_184;
  reg [31:0] _RAND_4;
  wire  _T_185;
  wire  _T_188;
  wire  _T_190;
  wire  _T_192;
  wire [15:0] _T_194;
  reg [15:0] _T_196;
  reg [31:0] _RAND_5;
  wire  _T_197;
  wire  _T_200;
  wire  _T_202;
  wire  _T_204;
  wire [15:0] _T_206;
  reg [15:0] _T_208;
  reg [31:0] _RAND_6;
  wire  _T_209;
  wire  _T_212;
  wire  _T_214;
  wire  _T_216;
  wire [15:0] _T_218;
  reg [15:0] _T_220;
  reg [31:0] _RAND_7;
  wire  _T_221;
  wire  _T_224;
  wire  _T_226;
  wire  _T_228;
  wire [15:0] _T_230;
  reg [15:0] _T_232;
  reg [31:0] _RAND_8;
  wire  _T_233;
  wire  _T_236;
  wire  _T_238;
  wire  _T_240;
  wire [15:0] _T_242;
  reg [15:0] _T_244;
  reg [31:0] _RAND_9;
  wire  _T_245;
  wire  _T_248;
  wire  _T_250;
  wire  _T_252;
  wire [15:0] _T_254;
  reg [15:0] _T_256;
  reg [31:0] _RAND_10;
  wire  _T_257;
  wire  _T_260;
  wire  _T_262;
  wire  _T_264;
  wire [15:0] _T_266;
  reg [15:0] _T_268;
  reg [31:0] _RAND_11;
  wire  _T_269;
  wire  _T_272;
  wire  _T_274;
  wire  _T_276;
  wire [15:0] _T_278;
  reg [15:0] _T_280;
  reg [31:0] _RAND_12;
  wire  _T_281;
  wire  _T_284;
  wire  _T_286;
  wire  _T_288;
  wire [15:0] _T_290;
  reg [15:0] _T_292;
  reg [31:0] _RAND_13;
  wire  _T_293;
  wire  _T_296;
  wire  _T_298;
  wire  _T_300;
  wire [15:0] _T_302;
  reg [15:0] _T_304;
  reg [31:0] _RAND_14;
  wire  _T_305;
  wire  _T_308;
  wire  _T_310;
  wire  _T_312;
  wire [15:0] _T_314;
  reg [15:0] _T_316;
  reg [31:0] _RAND_15;
  wire  _T_317;
  wire  _T_320;
  wire  _T_322;
  wire  _T_324;
  wire [15:0] _T_326;
  reg [15:0] _T_328;
  reg [31:0] _RAND_16;
  wire  _T_329;
  wire  _T_332;
  wire  _T_334;
  wire  _T_336;
  wire [15:0] _T_338;
  reg [15:0] _T_340;
  reg [31:0] _RAND_17;
  wire  _T_341;
  wire  _T_344;
  wire  _T_346;
  wire  _T_348;
  wire [15:0] _T_350;
  reg [15:0] _T_352;
  reg [31:0] _RAND_18;
  wire  _T_353;
  wire  _T_356;
  wire  _T_358;
  wire  _T_360;
  wire [15:0] _T_362;
  reg [15:0] _T_364;
  reg [31:0] _RAND_19;
  wire  _T_365;
  wire  _T_368;
  wire  _T_370;
  wire  _T_372;
  wire [15:0] _T_374;
  reg [15:0] _T_376;
  reg [31:0] _RAND_20;
  wire  _T_377;
  wire  _T_380;
  wire  _T_382;
  wire  _T_384;
  wire [15:0] _T_386;
  reg [15:0] _T_388;
  reg [31:0] _RAND_21;
  wire  _T_389;
  wire  _T_392;
  wire  _T_394;
  wire  _T_396;
  wire [15:0] _T_398;
  reg [15:0] _T_400;
  reg [31:0] _RAND_22;
  wire  _T_401;
  wire  _T_404;
  wire  _T_406;
  wire  _T_408;
  wire [15:0] _T_410;
  reg [15:0] _T_412;
  reg [31:0] _RAND_23;
  wire  _T_413;
  wire  _T_416;
  wire  _T_418;
  wire  _T_420;
  wire [15:0] _T_422;
  reg [15:0] _T_424;
  reg [31:0] _RAND_24;
  wire  _T_425;
  wire  _T_428;
  wire  _T_430;
  wire  _T_432;
  wire [15:0] _T_434;
  reg [15:0] _T_436;
  reg [31:0] _RAND_25;
  wire  _T_437;
  wire  _T_440;
  wire  _T_442;
  wire  _T_444;
  wire [15:0] _T_446;
  reg [15:0] _T_448;
  reg [31:0] _RAND_26;
  wire  _T_449;
  wire  _T_452;
  wire  _T_454;
  wire  _T_456;
  wire [15:0] _T_458;
  reg [15:0] _T_460;
  reg [31:0] _RAND_27;
  wire  _T_461;
  wire  _T_464;
  wire  _T_466;
  wire  _T_468;
  wire [15:0] _T_470;
  reg [15:0] _T_472;
  reg [31:0] _RAND_28;
  wire  _T_473;
  wire  _T_476;
  wire  _T_478;
  wire  _T_480;
  wire [15:0] _T_482;
  reg [15:0] _T_484;
  reg [31:0] _RAND_29;
  wire  _T_485;
  wire  _T_488;
  wire  _T_490;
  wire  _T_492;
  wire [15:0] _T_494;
  reg [15:0] _T_496;
  reg [31:0] _RAND_30;
  wire  _T_497;
  wire  _T_500;
  wire  _T_502;
  wire  _T_504;
  wire [15:0] _T_506;
  reg [15:0] _T_508;
  reg [31:0] _RAND_31;
  wire  _T_509;
  wire  _T_512;
  wire  _T_514;
  wire  _T_516;
  wire [15:0] _T_518;
  reg [15:0] _T_520;
  reg [31:0] _RAND_32;
  wire  _T_521;
  wire  _T_524;
  wire  _T_526;
  wire  _T_528;
  wire [15:0] _T_530;
  reg [15:0] _T_532;
  reg [31:0] _RAND_33;
  wire  _T_533;
  wire  _T_536;
  wire  _T_538;
  wire  _T_540;
  wire [15:0] _T_542;
  reg [15:0] _T_544;
  reg [31:0] _RAND_34;
  wire  _T_545;
  wire  _T_548;
  wire  _T_550;
  wire  _T_552;
  wire [15:0] _T_554;
  reg [15:0] _T_556;
  reg [31:0] _RAND_35;
  wire  _T_557;
  wire  _T_560;
  wire  _T_562;
  wire  _T_564;
  wire [15:0] _T_566;
  reg [15:0] _T_568;
  reg [31:0] _RAND_36;
  wire  _T_569;
  wire  _T_572;
  wire  _T_574;
  wire  _T_576;
  wire [15:0] _T_578;
  reg [15:0] _T_580;
  reg [31:0] _RAND_37;
  wire  _T_581;
  wire  _T_584;
  wire  _T_586;
  wire  _T_588;
  wire [15:0] _T_590;
  reg [15:0] _T_592;
  reg [31:0] _RAND_38;
  wire  _T_593;
  wire  _T_596;
  wire  _T_598;
  wire  _T_600;
  wire [15:0] _T_602;
  reg [15:0] _T_604;
  reg [31:0] _RAND_39;
  wire  _T_605;
  wire  _T_608;
  wire  _T_610;
  wire  _T_612;
  wire [15:0] _T_614;
  reg [15:0] _T_616;
  reg [31:0] _RAND_40;
  wire  _T_617;
  wire  _T_620;
  wire  _T_622;
  wire  _T_624;
  wire [15:0] _T_626;
  reg [15:0] _T_628;
  reg [31:0] _RAND_41;
  wire  _T_629;
  wire  _T_632;
  wire  _T_634;
  wire  _T_636;
  wire [15:0] _T_638;
  reg [15:0] _T_640;
  reg [31:0] _RAND_42;
  wire  _T_641;
  wire  _T_644;
  wire  _T_646;
  wire  _T_648;
  wire [15:0] _T_650;
  reg [15:0] _T_652;
  reg [31:0] _RAND_43;
  wire  _T_653;
  wire  _T_656;
  wire  _T_658;
  wire  _T_660;
  wire [15:0] _T_662;
  reg [15:0] _T_664;
  reg [31:0] _RAND_44;
  wire  _T_665;
  wire  _T_668;
  wire  _T_670;
  wire  _T_672;
  wire [15:0] _T_674;
  reg [15:0] _T_676;
  reg [31:0] _RAND_45;
  wire  _T_677;
  wire  _T_680;
  wire  _T_682;
  wire  _T_684;
  wire [15:0] _T_686;
  reg [15:0] _T_688;
  reg [31:0] _RAND_46;
  wire  _T_689;
  wire  _T_692;
  wire  _T_694;
  wire  _T_696;
  wire [15:0] _T_698;
  reg [15:0] _T_700;
  reg [31:0] _RAND_47;
  wire  _T_701;
  wire  _T_704;
  wire  _T_706;
  wire  _T_708;
  wire [15:0] _T_710;
  reg [15:0] _T_712;
  reg [31:0] _RAND_48;
  wire  _T_713;
  wire  _T_716;
  wire  _T_718;
  wire  _T_720;
  wire [15:0] _T_722;
  reg [15:0] _T_724;
  reg [31:0] _RAND_49;
  wire  _T_725;
  wire  _T_728;
  wire  _T_730;
  wire  _T_732;
  wire [15:0] _T_734;
  reg [15:0] _T_736;
  reg [31:0] _RAND_50;
  wire  _T_737;
  wire  _T_740;
  wire  _T_742;
  wire  _T_744;
  wire [15:0] _T_746;
  reg [15:0] _T_748;
  reg [31:0] _RAND_51;
  wire  _T_749;
  wire  _T_752;
  wire  _T_754;
  wire  _T_756;
  wire [15:0] _T_758;
  reg [15:0] _T_760;
  reg [31:0] _RAND_52;
  wire  _T_761;
  wire  _T_764;
  wire  _T_766;
  wire  _T_768;
  wire [15:0] _T_770;
  reg [15:0] _T_772;
  reg [31:0] _RAND_53;
  wire  _T_773;
  wire  _T_776;
  wire  _T_778;
  wire  _T_780;
  wire [15:0] _T_782;
  reg [15:0] _T_784;
  reg [31:0] _RAND_54;
  wire  _T_785;
  wire  _T_788;
  wire  _T_790;
  wire  _T_792;
  wire [15:0] _T_794;
  reg [15:0] _T_796;
  reg [31:0] _RAND_55;
  wire  _T_797;
  wire  _T_800;
  wire  _T_802;
  wire  _T_804;
  wire [15:0] _T_806;
  reg [15:0] _T_808;
  reg [31:0] _RAND_56;
  wire  _T_809;
  wire  _T_812;
  wire  _T_814;
  wire  _T_816;
  wire [15:0] _T_818;
  reg [15:0] _T_820;
  reg [31:0] _RAND_57;
  wire  _T_821;
  wire  _T_824;
  wire  _T_826;
  wire  _T_828;
  wire [15:0] _T_830;
  reg [15:0] _T_832;
  reg [31:0] _RAND_58;
  wire  _T_833;
  wire  _T_836;
  wire  _T_838;
  wire  _T_840;
  wire [15:0] _T_842;
  reg [15:0] _T_844;
  reg [31:0] _RAND_59;
  wire  _T_845;
  wire  _T_848;
  wire  _T_850;
  wire  _T_852;
  wire [15:0] _T_854;
  reg [15:0] _T_856;
  reg [31:0] _RAND_60;
  wire  _T_857;
  wire  _T_860;
  wire  _T_862;
  wire  _T_864;
  wire [15:0] _T_866;
  reg [15:0] _T_868;
  reg [31:0] _RAND_61;
  wire  _T_869;
  wire  _T_872;
  wire  _T_874;
  wire  _T_876;
  wire [15:0] _T_878;
  reg [15:0] _T_880;
  reg [31:0] _RAND_62;
  wire  _T_881;
  wire  _T_884;
  wire  _T_886;
  wire  _T_888;
  wire [15:0] _T_890;
  reg [15:0] _T_892;
  reg [31:0] _RAND_63;
  wire  _T_893;
  wire  _T_896;
  wire  _T_898;
  wire  _T_900;
  wire [15:0] _T_902;
  reg [15:0] _T_904;
  reg [31:0] _RAND_64;
  wire  _T_905;
  wire  _T_908;
  wire  _T_910;
  wire  _T_912;
  wire [15:0] _T_914;
  reg [15:0] _T_916;
  reg [31:0] _RAND_65;
  wire  _T_917;
  wire  _T_920;
  wire  _T_922;
  wire  _T_924;
  wire [15:0] _T_926;
  reg [15:0] _T_928;
  reg [31:0] _RAND_66;
  wire  _T_929;
  wire  _T_932;
  wire  _T_934;
  wire  _T_936;
  wire [15:0] _T_938;
  reg [15:0] _T_940;
  reg [31:0] _RAND_67;
  wire  _T_941;
  wire  _T_944;
  wire  _T_946;
  wire  _T_948;
  wire [15:0] _T_950;
  reg [15:0] _T_952;
  reg [31:0] _RAND_68;
  wire  _T_953;
  wire  _T_956;
  wire  _T_958;
  wire  _T_960;
  wire [15:0] _T_962;
  reg [15:0] _T_964;
  reg [31:0] _RAND_69;
  wire  _T_965;
  wire  _T_968;
  wire  _T_970;
  wire  _T_972;
  wire [15:0] _T_974;
  reg [15:0] _T_976;
  reg [31:0] _RAND_70;
  wire  _T_977;
  wire  _T_980;
  wire  _T_982;
  wire  _T_984;
  wire [15:0] _T_986;
  reg [15:0] _T_988;
  reg [31:0] _RAND_71;
  wire  _T_989;
  wire  _T_992;
  wire  _T_994;
  wire  _T_996;
  wire [15:0] _T_998;
  reg [15:0] _T_1000;
  reg [31:0] _RAND_72;
  wire  _T_1001;
  wire  _T_1004;
  wire  _T_1006;
  wire  _T_1008;
  wire [15:0] _T_1010;
  reg [15:0] _T_1012;
  reg [31:0] _RAND_73;
  wire  _T_1013;
  wire  _T_1016;
  wire  _T_1018;
  wire  _T_1020;
  wire [15:0] _T_1022;
  reg [15:0] _T_1024;
  reg [31:0] _RAND_74;
  wire  _T_1025;
  wire  _T_1028;
  wire  _T_1030;
  wire  _T_1032;
  wire [15:0] _T_1034;
  reg [15:0] _T_1036;
  reg [31:0] _RAND_75;
  wire  _T_1037;
  wire  _T_1040;
  wire  _T_1042;
  wire  _T_1044;
  wire [15:0] _T_1046;
  reg [15:0] _T_1048;
  reg [31:0] _RAND_76;
  wire  _T_1049;
  wire  _T_1052;
  wire  _T_1054;
  wire  _T_1056;
  wire [15:0] _T_1058;
  reg [15:0] _T_1060;
  reg [31:0] _RAND_77;
  wire  _T_1061;
  wire  _T_1064;
  wire  _T_1066;
  wire  _T_1068;
  wire [15:0] _T_1070;
  reg [15:0] _T_1072;
  reg [31:0] _RAND_78;
  wire  _T_1073;
  wire  _T_1076;
  wire  _T_1078;
  wire  _T_1080;
  wire [15:0] _T_1082;
  reg [15:0] _T_1084;
  reg [31:0] _RAND_79;
  wire  _T_1085;
  wire  _T_1088;
  wire  _T_1090;
  wire  _T_1092;
  wire [15:0] _T_1094;
  reg [15:0] _T_1096;
  reg [31:0] _RAND_80;
  wire  _T_1097;
  wire  _T_1100;
  wire  _T_1102;
  wire  _T_1104;
  wire [15:0] _T_1106;
  reg [15:0] _T_1108;
  reg [31:0] _RAND_81;
  wire  _T_1109;
  wire  _T_1112;
  wire  _T_1114;
  wire  _T_1116;
  wire [15:0] _T_1118;
  reg [15:0] _T_1120;
  reg [31:0] _RAND_82;
  wire  _T_1121;
  wire  _T_1124;
  wire  _T_1126;
  wire  _T_1128;
  wire [15:0] _T_1130;
  reg [15:0] _T_1132;
  reg [31:0] _RAND_83;
  wire  _T_1133;
  wire  _T_1136;
  wire  _T_1138;
  wire  _T_1140;
  wire [15:0] _T_1142;
  reg [15:0] _T_1144;
  reg [31:0] _RAND_84;
  wire  _T_1145;
  wire  _T_1148;
  wire  _T_1150;
  wire  _T_1152;
  wire [15:0] _T_1154;
  reg [15:0] _T_1156;
  reg [31:0] _RAND_85;
  wire  _T_1157;
  wire  _T_1160;
  wire  _T_1162;
  wire  _T_1164;
  wire [15:0] _T_1166;
  reg [15:0] _T_1168;
  reg [31:0] _RAND_86;
  wire  _T_1169;
  wire  _T_1172;
  wire  _T_1174;
  wire  _T_1176;
  wire [15:0] _T_1178;
  reg [15:0] _T_1180;
  reg [31:0] _RAND_87;
  wire  _T_1181;
  wire  _T_1184;
  wire  _T_1186;
  wire  _T_1188;
  wire [15:0] _T_1190;
  reg [15:0] _T_1192;
  reg [31:0] _RAND_88;
  wire  _T_1193;
  wire  _T_1196;
  wire  _T_1198;
  wire  _T_1200;
  wire [15:0] _T_1202;
  reg [15:0] _T_1204;
  reg [31:0] _RAND_89;
  wire  _T_1205;
  wire  _T_1208;
  wire  _T_1210;
  wire  _T_1212;
  wire [15:0] _T_1214;
  reg [15:0] _T_1216;
  reg [31:0] _RAND_90;
  wire  _T_1217;
  wire  _T_1220;
  wire  _T_1222;
  wire  _T_1224;
  wire [15:0] _T_1226;
  reg [15:0] _T_1228;
  reg [31:0] _RAND_91;
  wire  _T_1229;
  wire  _T_1232;
  wire  _T_1234;
  wire  _T_1236;
  wire [15:0] _T_1238;
  reg [15:0] _T_1240;
  reg [31:0] _RAND_92;
  wire  _T_1241;
  wire  _T_1244;
  wire  _T_1246;
  wire  _T_1248;
  wire [15:0] _T_1250;
  reg [15:0] _T_1252;
  reg [31:0] _RAND_93;
  wire  _T_1253;
  wire  _T_1256;
  wire  _T_1258;
  wire  _T_1260;
  wire [15:0] _T_1262;
  reg [15:0] _T_1264;
  reg [31:0] _RAND_94;
  wire  _T_1265;
  wire  _T_1268;
  wire  _T_1270;
  wire  _T_1272;
  wire [15:0] _T_1274;
  reg [15:0] _T_1276;
  reg [31:0] _RAND_95;
  wire  _T_1277;
  wire  _T_1280;
  wire  _T_1282;
  wire  _T_1284;
  wire [15:0] _T_1286;
  reg [15:0] _T_1288;
  reg [31:0] _RAND_96;
  wire  _T_1289;
  wire  _T_1292;
  wire  _T_1294;
  wire  _T_1296;
  wire [15:0] _T_1298;
  reg [15:0] _T_1300;
  reg [31:0] _RAND_97;
  wire  _T_1301;
  wire  _T_1304;
  wire  _T_1306;
  wire  _T_1308;
  wire [15:0] _T_1310;
  reg [15:0] _T_1312;
  reg [31:0] _RAND_98;
  wire  _T_1313;
  wire  _T_1316;
  wire  _T_1318;
  wire  _T_1320;
  wire [15:0] _T_1322;
  reg [15:0] _T_1324;
  reg [31:0] _RAND_99;
  wire  _T_1325;
  wire  _T_1328;
  wire  _T_1330;
  wire  _T_1332;
  wire [15:0] _T_1334;
  reg [15:0] _T_1336;
  reg [31:0] _RAND_100;
  wire  _T_1337;
  wire  _T_1340;
  wire  _T_1342;
  wire  _T_1344;
  wire [15:0] _T_1346;
  reg [15:0] _T_1348;
  reg [31:0] _RAND_101;
  wire  _T_1349;
  wire  _T_1352;
  wire  _T_1354;
  wire  _T_1356;
  wire [15:0] _T_1358;
  reg [15:0] _T_1360;
  reg [31:0] _RAND_102;
  wire  _T_1361;
  wire  _T_1364;
  wire  _T_1366;
  wire  _T_1368;
  wire [15:0] _T_1370;
  reg [15:0] _T_1372;
  reg [31:0] _RAND_103;
  wire  _T_1373;
  wire  _T_1376;
  wire  _T_1378;
  wire  _T_1380;
  wire [15:0] _T_1382;
  reg [15:0] _T_1384;
  reg [31:0] _RAND_104;
  wire  _T_1385;
  wire  _T_1388;
  wire  _T_1390;
  wire  _T_1392;
  wire [15:0] _T_1394;
  reg [15:0] _T_1396;
  reg [31:0] _RAND_105;
  wire  _T_1397;
  wire  _T_1400;
  wire  _T_1402;
  wire  _T_1404;
  wire [15:0] _T_1406;
  reg [15:0] _T_1408;
  reg [31:0] _RAND_106;
  wire  _T_1409;
  wire  _T_1412;
  wire  _T_1414;
  wire  _T_1416;
  wire [15:0] _T_1418;
  reg [15:0] _T_1420;
  reg [31:0] _RAND_107;
  wire  _T_1421;
  wire  _T_1424;
  wire  _T_1426;
  wire  _T_1428;
  wire [15:0] _T_1430;
  reg [15:0] _T_1432;
  reg [31:0] _RAND_108;
  wire  _T_1433;
  wire  _T_1436;
  wire  _T_1438;
  wire  _T_1440;
  wire [15:0] _T_1442;
  reg [15:0] _T_1444;
  reg [31:0] _RAND_109;
  wire  _T_1445;
  wire  _T_1448;
  wire  _T_1450;
  wire  _T_1452;
  wire [15:0] _T_1454;
  reg [15:0] _T_1456;
  reg [31:0] _RAND_110;
  wire  _T_1457;
  wire  _T_1460;
  wire  _T_1462;
  wire  _T_1464;
  wire [15:0] _T_1466;
  reg [15:0] _T_1468;
  reg [31:0] _RAND_111;
  wire  _T_1469;
  wire  _T_1472;
  wire  _T_1474;
  wire  _T_1476;
  wire [15:0] _T_1478;
  reg [15:0] _T_1480;
  reg [31:0] _RAND_112;
  wire  _T_1481;
  wire  _T_1484;
  wire  _T_1486;
  wire  _T_1488;
  wire [15:0] _T_1490;
  reg [15:0] _T_1492;
  reg [31:0] _RAND_113;
  wire  _T_1493;
  wire  _T_1496;
  wire  _T_1498;
  wire  _T_1500;
  wire [15:0] _T_1502;
  reg [15:0] _T_1504;
  reg [31:0] _RAND_114;
  wire  _T_1505;
  wire  _T_1508;
  wire  _T_1510;
  wire  _T_1512;
  wire [15:0] _T_1514;
  reg [15:0] _T_1516;
  reg [31:0] _RAND_115;
  wire  _T_1517;
  wire  _T_1520;
  wire  _T_1522;
  wire  _T_1524;
  wire [15:0] _T_1526;
  reg [15:0] _T_1528;
  reg [31:0] _RAND_116;
  wire  _T_1529;
  wire  _T_1532;
  wire  _T_1534;
  wire  _T_1536;
  wire [15:0] _T_1538;
  reg [15:0] _T_1540;
  reg [31:0] _RAND_117;
  wire  _T_1541;
  wire  _T_1544;
  wire  _T_1546;
  wire  _T_1548;
  wire [15:0] _T_1550;
  reg [15:0] _T_1552;
  reg [31:0] _RAND_118;
  wire  _T_1553;
  wire  _T_1556;
  wire  _T_1558;
  wire  _T_1560;
  wire [15:0] _T_1562;
  reg [15:0] _T_1564;
  reg [31:0] _RAND_119;
  wire  _T_1565;
  wire  _T_1568;
  wire  _T_1570;
  wire  _T_1572;
  wire [15:0] _T_1574;
  reg [15:0] _T_1576;
  reg [31:0] _RAND_120;
  wire  _T_1577;
  wire  _T_1580;
  wire  _T_1582;
  wire  _T_1584;
  wire [15:0] _T_1586;
  reg [15:0] _T_1588;
  reg [31:0] _RAND_121;
  wire  _T_1589;
  wire  _T_1592;
  wire  _T_1594;
  wire  _T_1596;
  wire [15:0] _T_1598;
  reg [15:0] _T_1600;
  reg [31:0] _RAND_122;
  wire  _T_1601;
  wire  _T_1604;
  wire  _T_1606;
  wire  _T_1608;
  wire [15:0] _T_1610;
  reg [15:0] _T_1612;
  reg [31:0] _RAND_123;
  wire  _T_1613;
  wire  _T_1616;
  wire  _T_1618;
  wire  _T_1620;
  wire [15:0] _T_1622;
  reg [15:0] _T_1624;
  reg [31:0] _RAND_124;
  wire  _T_1625;
  wire  _T_1628;
  wire  _T_1630;
  wire  _T_1632;
  wire [15:0] _T_1634;
  reg [15:0] _T_1636;
  reg [31:0] _RAND_125;
  wire  _T_1637;
  wire  _T_1640;
  wire  _T_1642;
  wire  _T_1644;
  wire [15:0] _T_1646;
  reg [15:0] _T_1648;
  reg [31:0] _RAND_126;
  wire  _T_1649;
  wire  _T_1652;
  wire  _T_1654;
  wire  _T_1656;
  wire [15:0] _T_1658;
  reg [15:0] _T_1660;
  reg [31:0] _RAND_127;
  wire  _T_1661;
  wire  _T_1664;
  wire  _T_1666;
  wire  _T_1668;
  wire [15:0] _T_1670;
  reg [15:0] _T_1672;
  reg [31:0] _RAND_128;
  wire  _T_1673;
  wire  _T_1676;
  wire  _T_1678;
  wire  _T_1680;
  wire [15:0] _T_1682;
  reg [15:0] _T_1684;
  reg [31:0] _RAND_129;
  wire  _T_1685;
  wire  _T_1688;
  wire  _T_1690;
  wire  _T_1692;
  wire [15:0] _T_1694;
  reg [15:0] _T_1696;
  reg [31:0] _RAND_130;
  wire  _T_1697;
  wire  _T_1700;
  wire  _T_1702;
  wire  _T_1704;
  wire [15:0] _T_1706;
  wire [6:0] _T_1715;
  wire [14:0] _T_1723;
  wire [7:0] _T_1730;
  wire [30:0] _T_1739;
  wire [7:0] _T_1746;
  wire [15:0] _T_1754;
  wire [7:0] _T_1761;
  wire [31:0] _T_1770;
  wire [7:0] _T_1778;
  wire [15:0] _T_1786;
  wire [7:0] _T_1793;
  wire [31:0] _T_1802;
  wire [7:0] _T_1809;
  wire [15:0] _T_1817;
  wire [7:0] _T_1824;
  wire [31:0] _T_1833;
  wire [126:0] _T_1835;
  wire  _T_1836;
  wire  _T_1837;
  reg [15:0] _T_1838;
  reg [31:0] _RAND_131;
  wire  _T_1839;
  wire  _T_1842;
  wire  _T_1844;
  wire  _T_1846;
  wire [15:0] _T_1848;
  reg [15:0] _T_1850;
  reg [31:0] _RAND_132;
  wire  _T_1851;
  wire  _T_1854;
  wire  _T_1856;
  wire  _T_1858;
  wire [15:0] _T_1860;
  reg [15:0] _T_1862;
  reg [31:0] _RAND_133;
  wire  _T_1863;
  wire  _T_1866;
  wire  _T_1868;
  wire  _T_1870;
  wire [15:0] _T_1872;
  reg [15:0] _T_1874;
  reg [31:0] _RAND_134;
  wire  _T_1875;
  wire  _T_1878;
  wire  _T_1880;
  wire  _T_1882;
  wire [15:0] _T_1884;
  reg [15:0] _T_1886;
  reg [31:0] _RAND_135;
  wire  _T_1887;
  wire  _T_1890;
  wire  _T_1892;
  wire  _T_1894;
  wire [15:0] _T_1896;
  reg [15:0] _T_1898;
  reg [31:0] _RAND_136;
  wire  _T_1899;
  wire  _T_1902;
  wire  _T_1904;
  wire  _T_1906;
  wire [15:0] _T_1908;
  reg [15:0] _T_1910;
  reg [31:0] _RAND_137;
  wire  _T_1911;
  wire  _T_1914;
  wire  _T_1916;
  wire  _T_1918;
  wire [15:0] _T_1920;
  reg [15:0] _T_1922;
  reg [31:0] _RAND_138;
  wire  _T_1923;
  wire  _T_1926;
  wire  _T_1928;
  wire  _T_1930;
  wire [15:0] _T_1932;
  reg [15:0] _T_1934;
  reg [31:0] _RAND_139;
  wire  _T_1935;
  wire  _T_1938;
  wire  _T_1940;
  wire  _T_1942;
  wire [15:0] _T_1944;
  reg [15:0] _T_1946;
  reg [31:0] _RAND_140;
  wire  _T_1947;
  wire  _T_1950;
  wire  _T_1952;
  wire  _T_1954;
  wire [15:0] _T_1956;
  reg [15:0] _T_1958;
  reg [31:0] _RAND_141;
  wire  _T_1959;
  wire  _T_1962;
  wire  _T_1964;
  wire  _T_1966;
  wire [15:0] _T_1968;
  reg [15:0] _T_1970;
  reg [31:0] _RAND_142;
  wire  _T_1971;
  wire  _T_1974;
  wire  _T_1976;
  wire  _T_1978;
  wire [15:0] _T_1980;
  reg [15:0] _T_1982;
  reg [31:0] _RAND_143;
  wire  _T_1983;
  wire  _T_1986;
  wire  _T_1988;
  wire  _T_1990;
  wire [15:0] _T_1992;
  reg [15:0] _T_1994;
  reg [31:0] _RAND_144;
  wire  _T_1995;
  wire  _T_1998;
  wire  _T_2000;
  wire  _T_2002;
  wire [15:0] _T_2004;
  reg [15:0] _T_2006;
  reg [31:0] _RAND_145;
  wire  _T_2007;
  wire  _T_2010;
  wire  _T_2012;
  wire  _T_2014;
  wire [15:0] _T_2016;
  reg [15:0] _T_2018;
  reg [31:0] _RAND_146;
  wire  _T_2019;
  wire  _T_2022;
  wire  _T_2024;
  wire  _T_2026;
  wire [15:0] _T_2028;
  reg [15:0] _T_2030;
  reg [31:0] _RAND_147;
  wire  _T_2031;
  wire  _T_2034;
  wire  _T_2036;
  wire  _T_2038;
  wire [15:0] _T_2040;
  reg [15:0] _T_2042;
  reg [31:0] _RAND_148;
  wire  _T_2043;
  wire  _T_2046;
  wire  _T_2048;
  wire  _T_2050;
  wire [15:0] _T_2052;
  reg [15:0] _T_2054;
  reg [31:0] _RAND_149;
  wire  _T_2055;
  wire  _T_2058;
  wire  _T_2060;
  wire  _T_2062;
  wire [15:0] _T_2064;
  reg [15:0] _T_2066;
  reg [31:0] _RAND_150;
  wire  _T_2067;
  wire  _T_2070;
  wire  _T_2072;
  wire  _T_2074;
  wire [15:0] _T_2076;
  reg [15:0] _T_2078;
  reg [31:0] _RAND_151;
  wire  _T_2079;
  wire  _T_2082;
  wire  _T_2084;
  wire  _T_2086;
  wire [15:0] _T_2088;
  reg [15:0] _T_2090;
  reg [31:0] _RAND_152;
  wire  _T_2091;
  wire  _T_2094;
  wire  _T_2096;
  wire  _T_2098;
  wire [15:0] _T_2100;
  reg [15:0] _T_2102;
  reg [31:0] _RAND_153;
  wire  _T_2103;
  wire  _T_2106;
  wire  _T_2108;
  wire  _T_2110;
  wire [15:0] _T_2112;
  reg [15:0] _T_2114;
  reg [31:0] _RAND_154;
  wire  _T_2115;
  wire  _T_2118;
  wire  _T_2120;
  wire  _T_2122;
  wire [15:0] _T_2124;
  reg [15:0] _T_2126;
  reg [31:0] _RAND_155;
  wire  _T_2127;
  wire  _T_2130;
  wire  _T_2132;
  wire  _T_2134;
  wire [15:0] _T_2136;
  reg [15:0] _T_2138;
  reg [31:0] _RAND_156;
  wire  _T_2139;
  wire  _T_2142;
  wire  _T_2144;
  wire  _T_2146;
  wire [15:0] _T_2148;
  reg [15:0] _T_2150;
  reg [31:0] _RAND_157;
  wire  _T_2151;
  wire  _T_2154;
  wire  _T_2156;
  wire  _T_2158;
  wire [15:0] _T_2160;
  reg [15:0] _T_2162;
  reg [31:0] _RAND_158;
  wire  _T_2163;
  wire  _T_2166;
  wire  _T_2168;
  wire  _T_2170;
  wire [15:0] _T_2172;
  reg [15:0] _T_2174;
  reg [31:0] _RAND_159;
  wire  _T_2175;
  wire  _T_2178;
  wire  _T_2180;
  wire  _T_2182;
  wire [15:0] _T_2184;
  reg [15:0] _T_2186;
  reg [31:0] _RAND_160;
  wire  _T_2187;
  wire  _T_2190;
  wire  _T_2192;
  wire  _T_2194;
  wire [15:0] _T_2196;
  reg [15:0] _T_2198;
  reg [31:0] _RAND_161;
  wire  _T_2199;
  wire  _T_2202;
  wire  _T_2204;
  wire  _T_2206;
  wire [15:0] _T_2208;
  reg [15:0] _T_2210;
  reg [31:0] _RAND_162;
  wire  _T_2211;
  wire  _T_2214;
  wire  _T_2216;
  wire  _T_2218;
  wire [15:0] _T_2220;
  reg [15:0] _T_2222;
  reg [31:0] _RAND_163;
  wire  _T_2223;
  wire  _T_2226;
  wire  _T_2228;
  wire  _T_2230;
  wire [15:0] _T_2232;
  reg [15:0] _T_2234;
  reg [31:0] _RAND_164;
  wire  _T_2235;
  wire  _T_2238;
  wire  _T_2240;
  wire  _T_2242;
  wire [15:0] _T_2244;
  reg [15:0] _T_2246;
  reg [31:0] _RAND_165;
  wire  _T_2247;
  wire  _T_2250;
  wire  _T_2252;
  wire  _T_2254;
  wire [15:0] _T_2256;
  reg [15:0] _T_2258;
  reg [31:0] _RAND_166;
  wire  _T_2259;
  wire  _T_2262;
  wire  _T_2264;
  wire  _T_2266;
  wire [15:0] _T_2268;
  reg [15:0] _T_2270;
  reg [31:0] _RAND_167;
  wire  _T_2271;
  wire  _T_2274;
  wire  _T_2276;
  wire  _T_2278;
  wire [15:0] _T_2280;
  reg [15:0] _T_2282;
  reg [31:0] _RAND_168;
  wire  _T_2283;
  wire  _T_2286;
  wire  _T_2288;
  wire  _T_2290;
  wire [15:0] _T_2292;
  reg [15:0] _T_2294;
  reg [31:0] _RAND_169;
  wire  _T_2295;
  wire  _T_2298;
  wire  _T_2300;
  wire  _T_2302;
  wire [15:0] _T_2304;
  reg [15:0] _T_2306;
  reg [31:0] _RAND_170;
  wire  _T_2307;
  wire  _T_2310;
  wire  _T_2312;
  wire  _T_2314;
  wire [15:0] _T_2316;
  reg [15:0] _T_2318;
  reg [31:0] _RAND_171;
  wire  _T_2319;
  wire  _T_2322;
  wire  _T_2324;
  wire  _T_2326;
  wire [15:0] _T_2328;
  reg [15:0] _T_2330;
  reg [31:0] _RAND_172;
  wire  _T_2331;
  wire  _T_2334;
  wire  _T_2336;
  wire  _T_2338;
  wire [15:0] _T_2340;
  reg [15:0] _T_2342;
  reg [31:0] _RAND_173;
  wire  _T_2343;
  wire  _T_2346;
  wire  _T_2348;
  wire  _T_2350;
  wire [15:0] _T_2352;
  reg [15:0] _T_2354;
  reg [31:0] _RAND_174;
  wire  _T_2355;
  wire  _T_2358;
  wire  _T_2360;
  wire  _T_2362;
  wire [15:0] _T_2364;
  reg [15:0] _T_2366;
  reg [31:0] _RAND_175;
  wire  _T_2367;
  wire  _T_2370;
  wire  _T_2372;
  wire  _T_2374;
  wire [15:0] _T_2376;
  reg [15:0] _T_2378;
  reg [31:0] _RAND_176;
  wire  _T_2379;
  wire  _T_2382;
  wire  _T_2384;
  wire  _T_2386;
  wire [15:0] _T_2388;
  reg [15:0] _T_2390;
  reg [31:0] _RAND_177;
  wire  _T_2391;
  wire  _T_2394;
  wire  _T_2396;
  wire  _T_2398;
  wire [15:0] _T_2400;
  reg [15:0] _T_2402;
  reg [31:0] _RAND_178;
  wire  _T_2403;
  wire  _T_2406;
  wire  _T_2408;
  wire  _T_2410;
  wire [15:0] _T_2412;
  reg [15:0] _T_2414;
  reg [31:0] _RAND_179;
  wire  _T_2415;
  wire  _T_2418;
  wire  _T_2420;
  wire  _T_2422;
  wire [15:0] _T_2424;
  reg [15:0] _T_2426;
  reg [31:0] _RAND_180;
  wire  _T_2427;
  wire  _T_2430;
  wire  _T_2432;
  wire  _T_2434;
  wire [15:0] _T_2436;
  reg [15:0] _T_2438;
  reg [31:0] _RAND_181;
  wire  _T_2439;
  wire  _T_2442;
  wire  _T_2444;
  wire  _T_2446;
  wire [15:0] _T_2448;
  reg [15:0] _T_2450;
  reg [31:0] _RAND_182;
  wire  _T_2451;
  wire  _T_2454;
  wire  _T_2456;
  wire  _T_2458;
  wire [15:0] _T_2460;
  reg [15:0] _T_2462;
  reg [31:0] _RAND_183;
  wire  _T_2463;
  wire  _T_2466;
  wire  _T_2468;
  wire  _T_2470;
  wire [15:0] _T_2472;
  reg [15:0] _T_2474;
  reg [31:0] _RAND_184;
  wire  _T_2475;
  wire  _T_2478;
  wire  _T_2480;
  wire  _T_2482;
  wire [15:0] _T_2484;
  reg [15:0] _T_2486;
  reg [31:0] _RAND_185;
  wire  _T_2487;
  wire  _T_2490;
  wire  _T_2492;
  wire  _T_2494;
  wire [15:0] _T_2496;
  reg [15:0] _T_2498;
  reg [31:0] _RAND_186;
  wire  _T_2499;
  wire  _T_2502;
  wire  _T_2504;
  wire  _T_2506;
  wire [15:0] _T_2508;
  reg [15:0] _T_2510;
  reg [31:0] _RAND_187;
  wire  _T_2511;
  wire  _T_2514;
  wire  _T_2516;
  wire  _T_2518;
  wire [15:0] _T_2520;
  reg [15:0] _T_2522;
  reg [31:0] _RAND_188;
  wire  _T_2523;
  wire  _T_2526;
  wire  _T_2528;
  wire  _T_2530;
  wire [15:0] _T_2532;
  reg [15:0] _T_2534;
  reg [31:0] _RAND_189;
  wire  _T_2535;
  wire  _T_2538;
  wire  _T_2540;
  wire  _T_2542;
  wire [15:0] _T_2544;
  reg [15:0] _T_2546;
  reg [31:0] _RAND_190;
  wire  _T_2547;
  wire  _T_2550;
  wire  _T_2552;
  wire  _T_2554;
  wire [15:0] _T_2556;
  reg [15:0] _T_2558;
  reg [31:0] _RAND_191;
  wire  _T_2559;
  wire  _T_2562;
  wire  _T_2564;
  wire  _T_2566;
  wire [15:0] _T_2568;
  reg [15:0] _T_2570;
  reg [31:0] _RAND_192;
  wire  _T_2571;
  wire  _T_2574;
  wire  _T_2576;
  wire  _T_2578;
  wire [15:0] _T_2580;
  reg [15:0] _T_2582;
  reg [31:0] _RAND_193;
  wire  _T_2583;
  wire  _T_2586;
  wire  _T_2588;
  wire  _T_2590;
  wire [15:0] _T_2592;
  reg [15:0] _T_2594;
  reg [31:0] _RAND_194;
  wire  _T_2595;
  wire  _T_2598;
  wire  _T_2600;
  wire  _T_2602;
  wire [15:0] _T_2604;
  reg [15:0] _T_2606;
  reg [31:0] _RAND_195;
  wire  _T_2607;
  wire  _T_2610;
  wire  _T_2612;
  wire  _T_2614;
  wire [15:0] _T_2616;
  reg [15:0] _T_2618;
  reg [31:0] _RAND_196;
  wire  _T_2619;
  wire  _T_2622;
  wire  _T_2624;
  wire  _T_2626;
  wire [15:0] _T_2628;
  reg [15:0] _T_2630;
  reg [31:0] _RAND_197;
  wire  _T_2631;
  wire  _T_2634;
  wire  _T_2636;
  wire  _T_2638;
  wire [15:0] _T_2640;
  reg [15:0] _T_2642;
  reg [31:0] _RAND_198;
  wire  _T_2643;
  wire  _T_2646;
  wire  _T_2648;
  wire  _T_2650;
  wire [15:0] _T_2652;
  reg [15:0] _T_2654;
  reg [31:0] _RAND_199;
  wire  _T_2655;
  wire  _T_2658;
  wire  _T_2660;
  wire  _T_2662;
  wire [15:0] _T_2664;
  reg [15:0] _T_2666;
  reg [31:0] _RAND_200;
  wire  _T_2667;
  wire  _T_2670;
  wire  _T_2672;
  wire  _T_2674;
  wire [15:0] _T_2676;
  reg [15:0] _T_2678;
  reg [31:0] _RAND_201;
  wire  _T_2679;
  wire  _T_2682;
  wire  _T_2684;
  wire  _T_2686;
  wire [15:0] _T_2688;
  reg [15:0] _T_2690;
  reg [31:0] _RAND_202;
  wire  _T_2691;
  wire  _T_2694;
  wire  _T_2696;
  wire  _T_2698;
  wire [15:0] _T_2700;
  reg [15:0] _T_2702;
  reg [31:0] _RAND_203;
  wire  _T_2703;
  wire  _T_2706;
  wire  _T_2708;
  wire  _T_2710;
  wire [15:0] _T_2712;
  reg [15:0] _T_2714;
  reg [31:0] _RAND_204;
  wire  _T_2715;
  wire  _T_2718;
  wire  _T_2720;
  wire  _T_2722;
  wire [15:0] _T_2724;
  reg [15:0] _T_2726;
  reg [31:0] _RAND_205;
  wire  _T_2727;
  wire  _T_2730;
  wire  _T_2732;
  wire  _T_2734;
  wire [15:0] _T_2736;
  reg [15:0] _T_2738;
  reg [31:0] _RAND_206;
  wire  _T_2739;
  wire  _T_2742;
  wire  _T_2744;
  wire  _T_2746;
  wire [15:0] _T_2748;
  reg [15:0] _T_2750;
  reg [31:0] _RAND_207;
  wire  _T_2751;
  wire  _T_2754;
  wire  _T_2756;
  wire  _T_2758;
  wire [15:0] _T_2760;
  reg [15:0] _T_2762;
  reg [31:0] _RAND_208;
  wire  _T_2763;
  wire  _T_2766;
  wire  _T_2768;
  wire  _T_2770;
  wire [15:0] _T_2772;
  reg [15:0] _T_2774;
  reg [31:0] _RAND_209;
  wire  _T_2775;
  wire  _T_2778;
  wire  _T_2780;
  wire  _T_2782;
  wire [15:0] _T_2784;
  reg [15:0] _T_2786;
  reg [31:0] _RAND_210;
  wire  _T_2787;
  wire  _T_2790;
  wire  _T_2792;
  wire  _T_2794;
  wire [15:0] _T_2796;
  reg [15:0] _T_2798;
  reg [31:0] _RAND_211;
  wire  _T_2799;
  wire  _T_2802;
  wire  _T_2804;
  wire  _T_2806;
  wire [15:0] _T_2808;
  reg [15:0] _T_2810;
  reg [31:0] _RAND_212;
  wire  _T_2811;
  wire  _T_2814;
  wire  _T_2816;
  wire  _T_2818;
  wire [15:0] _T_2820;
  reg [15:0] _T_2822;
  reg [31:0] _RAND_213;
  wire  _T_2823;
  wire  _T_2826;
  wire  _T_2828;
  wire  _T_2830;
  wire [15:0] _T_2832;
  reg [15:0] _T_2834;
  reg [31:0] _RAND_214;
  wire  _T_2835;
  wire  _T_2838;
  wire  _T_2840;
  wire  _T_2842;
  wire [15:0] _T_2844;
  reg [15:0] _T_2846;
  reg [31:0] _RAND_215;
  wire  _T_2847;
  wire  _T_2850;
  wire  _T_2852;
  wire  _T_2854;
  wire [15:0] _T_2856;
  reg [15:0] _T_2858;
  reg [31:0] _RAND_216;
  wire  _T_2859;
  wire  _T_2862;
  wire  _T_2864;
  wire  _T_2866;
  wire [15:0] _T_2868;
  reg [15:0] _T_2870;
  reg [31:0] _RAND_217;
  wire  _T_2871;
  wire  _T_2874;
  wire  _T_2876;
  wire  _T_2878;
  wire [15:0] _T_2880;
  reg [15:0] _T_2882;
  reg [31:0] _RAND_218;
  wire  _T_2883;
  wire  _T_2886;
  wire  _T_2888;
  wire  _T_2890;
  wire [15:0] _T_2892;
  reg [15:0] _T_2894;
  reg [31:0] _RAND_219;
  wire  _T_2895;
  wire  _T_2898;
  wire  _T_2900;
  wire  _T_2902;
  wire [15:0] _T_2904;
  reg [15:0] _T_2906;
  reg [31:0] _RAND_220;
  wire  _T_2907;
  wire  _T_2910;
  wire  _T_2912;
  wire  _T_2914;
  wire [15:0] _T_2916;
  reg [15:0] _T_2918;
  reg [31:0] _RAND_221;
  wire  _T_2919;
  wire  _T_2922;
  wire  _T_2924;
  wire  _T_2926;
  wire [15:0] _T_2928;
  reg [15:0] _T_2930;
  reg [31:0] _RAND_222;
  wire  _T_2931;
  wire  _T_2934;
  wire  _T_2936;
  wire  _T_2938;
  wire [15:0] _T_2940;
  reg [15:0] _T_2942;
  reg [31:0] _RAND_223;
  wire  _T_2943;
  wire  _T_2946;
  wire  _T_2948;
  wire  _T_2950;
  wire [15:0] _T_2952;
  reg [15:0] _T_2954;
  reg [31:0] _RAND_224;
  wire  _T_2955;
  wire  _T_2958;
  wire  _T_2960;
  wire  _T_2962;
  wire [15:0] _T_2964;
  reg [15:0] _T_2966;
  reg [31:0] _RAND_225;
  wire  _T_2967;
  wire  _T_2970;
  wire  _T_2972;
  wire  _T_2974;
  wire [15:0] _T_2976;
  reg [15:0] _T_2978;
  reg [31:0] _RAND_226;
  wire  _T_2979;
  wire  _T_2982;
  wire  _T_2984;
  wire  _T_2986;
  wire [15:0] _T_2988;
  reg [15:0] _T_2990;
  reg [31:0] _RAND_227;
  wire  _T_2991;
  wire  _T_2994;
  wire  _T_2996;
  wire  _T_2998;
  wire [15:0] _T_3000;
  reg [15:0] _T_3002;
  reg [31:0] _RAND_228;
  wire  _T_3003;
  wire  _T_3006;
  wire  _T_3008;
  wire  _T_3010;
  wire [15:0] _T_3012;
  reg [15:0] _T_3014;
  reg [31:0] _RAND_229;
  wire  _T_3015;
  wire  _T_3018;
  wire  _T_3020;
  wire  _T_3022;
  wire [15:0] _T_3024;
  reg [15:0] _T_3026;
  reg [31:0] _RAND_230;
  wire  _T_3027;
  wire  _T_3030;
  wire  _T_3032;
  wire  _T_3034;
  wire [15:0] _T_3036;
  reg [15:0] _T_3038;
  reg [31:0] _RAND_231;
  wire  _T_3039;
  wire  _T_3042;
  wire  _T_3044;
  wire  _T_3046;
  wire [15:0] _T_3048;
  reg [15:0] _T_3050;
  reg [31:0] _RAND_232;
  wire  _T_3051;
  wire  _T_3054;
  wire  _T_3056;
  wire  _T_3058;
  wire [15:0] _T_3060;
  reg [15:0] _T_3062;
  reg [31:0] _RAND_233;
  wire  _T_3063;
  wire  _T_3066;
  wire  _T_3068;
  wire  _T_3070;
  wire [15:0] _T_3072;
  reg [15:0] _T_3074;
  reg [31:0] _RAND_234;
  wire  _T_3075;
  wire  _T_3078;
  wire  _T_3080;
  wire  _T_3082;
  wire [15:0] _T_3084;
  reg [15:0] _T_3086;
  reg [31:0] _RAND_235;
  wire  _T_3087;
  wire  _T_3090;
  wire  _T_3092;
  wire  _T_3094;
  wire [15:0] _T_3096;
  reg [15:0] _T_3098;
  reg [31:0] _RAND_236;
  wire  _T_3099;
  wire  _T_3102;
  wire  _T_3104;
  wire  _T_3106;
  wire [15:0] _T_3108;
  reg [15:0] _T_3110;
  reg [31:0] _RAND_237;
  wire  _T_3111;
  wire  _T_3114;
  wire  _T_3116;
  wire  _T_3118;
  wire [15:0] _T_3120;
  reg [15:0] _T_3122;
  reg [31:0] _RAND_238;
  wire  _T_3123;
  wire  _T_3126;
  wire  _T_3128;
  wire  _T_3130;
  wire [15:0] _T_3132;
  reg [15:0] _T_3134;
  reg [31:0] _RAND_239;
  wire  _T_3135;
  wire  _T_3138;
  wire  _T_3140;
  wire  _T_3142;
  wire [15:0] _T_3144;
  reg [15:0] _T_3146;
  reg [31:0] _RAND_240;
  wire  _T_3147;
  wire  _T_3150;
  wire  _T_3152;
  wire  _T_3154;
  wire [15:0] _T_3156;
  reg [15:0] _T_3158;
  reg [31:0] _RAND_241;
  wire  _T_3159;
  wire  _T_3162;
  wire  _T_3164;
  wire  _T_3166;
  wire [15:0] _T_3168;
  reg [15:0] _T_3170;
  reg [31:0] _RAND_242;
  wire  _T_3171;
  wire  _T_3174;
  wire  _T_3176;
  wire  _T_3178;
  wire [15:0] _T_3180;
  reg [15:0] _T_3182;
  reg [31:0] _RAND_243;
  wire  _T_3183;
  wire  _T_3186;
  wire  _T_3188;
  wire  _T_3190;
  wire [15:0] _T_3192;
  reg [15:0] _T_3194;
  reg [31:0] _RAND_244;
  wire  _T_3195;
  wire  _T_3198;
  wire  _T_3200;
  wire  _T_3202;
  wire [15:0] _T_3204;
  reg [15:0] _T_3206;
  reg [31:0] _RAND_245;
  wire  _T_3207;
  wire  _T_3210;
  wire  _T_3212;
  wire  _T_3214;
  wire [15:0] _T_3216;
  reg [15:0] _T_3218;
  reg [31:0] _RAND_246;
  wire  _T_3219;
  wire  _T_3222;
  wire  _T_3224;
  wire  _T_3226;
  wire [15:0] _T_3228;
  reg [15:0] _T_3230;
  reg [31:0] _RAND_247;
  wire  _T_3231;
  wire  _T_3234;
  wire  _T_3236;
  wire  _T_3238;
  wire [15:0] _T_3240;
  reg [15:0] _T_3242;
  reg [31:0] _RAND_248;
  wire  _T_3243;
  wire  _T_3246;
  wire  _T_3248;
  wire  _T_3250;
  wire [15:0] _T_3252;
  reg [15:0] _T_3254;
  reg [31:0] _RAND_249;
  wire  _T_3255;
  wire  _T_3258;
  wire  _T_3260;
  wire  _T_3262;
  wire [15:0] _T_3264;
  reg [15:0] _T_3266;
  reg [31:0] _RAND_250;
  wire  _T_3267;
  wire  _T_3270;
  wire  _T_3272;
  wire  _T_3274;
  wire [15:0] _T_3276;
  reg [15:0] _T_3278;
  reg [31:0] _RAND_251;
  wire  _T_3279;
  wire  _T_3282;
  wire  _T_3284;
  wire  _T_3286;
  wire [15:0] _T_3288;
  reg [15:0] _T_3290;
  reg [31:0] _RAND_252;
  wire  _T_3291;
  wire  _T_3294;
  wire  _T_3296;
  wire  _T_3298;
  wire [15:0] _T_3300;
  reg [15:0] _T_3302;
  reg [31:0] _RAND_253;
  wire  _T_3303;
  wire  _T_3306;
  wire  _T_3308;
  wire  _T_3310;
  wire [15:0] _T_3312;
  reg [15:0] _T_3314;
  reg [31:0] _RAND_254;
  wire  _T_3315;
  wire  _T_3318;
  wire  _T_3320;
  wire  _T_3322;
  wire [15:0] _T_3324;
  reg [15:0] _T_3326;
  reg [31:0] _RAND_255;
  wire  _T_3327;
  wire  _T_3330;
  wire  _T_3332;
  wire  _T_3334;
  wire [15:0] _T_3336;
  reg [15:0] _T_3338;
  reg [31:0] _RAND_256;
  wire  _T_3339;
  wire  _T_3342;
  wire  _T_3344;
  wire  _T_3346;
  wire [15:0] _T_3348;
  reg [15:0] _T_3350;
  reg [31:0] _RAND_257;
  wire  _T_3351;
  wire  _T_3354;
  wire  _T_3356;
  wire  _T_3358;
  wire [15:0] _T_3360;
  wire [6:0] _T_3369;
  wire [14:0] _T_3377;
  wire [7:0] _T_3384;
  wire [30:0] _T_3393;
  wire [7:0] _T_3400;
  wire [15:0] _T_3408;
  wire [7:0] _T_3415;
  wire [31:0] _T_3424;
  wire [7:0] _T_3432;
  wire [15:0] _T_3440;
  wire [7:0] _T_3447;
  wire [31:0] _T_3456;
  wire [7:0] _T_3463;
  wire [15:0] _T_3471;
  wire [7:0] _T_3478;
  wire [31:0] _T_3487;
  wire [126:0] _T_3489;
  wire [126:0] _GEN_514;
  wire [126:0] _GEN_515;
  wire [126:0] _GEN_516;
  wire [127:0] _GEN_517;
  wire [127:0] _GEN_518;
  wire [127:0] _GEN_519;
  wire [127:0] _GEN_520;
  wire [15:0] _T_18;
  wire [142:0] _T_19;
  wire [7:0] _T_25;
  wire  _GEN_521;
  wire  _GEN_522;
  wire  _GEN_523;
  wire  _GEN_524;
  wire  _GEN_525;
  wire  _GEN_526;
  wire  _GEN_527;
  wire  _GEN_528;
  wire  _GEN_529;
  wire  _GEN_539;
  wire  _GEN_540;
  wire  _GEN_541;
  wire  _GEN_542;
  wire  _GEN_543;
  wire  _GEN_544;
  wire  _GEN_545;
  wire  _GEN_546;
  wire  _GEN_547;
  wire  _GEN_548;
  wire  _GEN_549;
  SiFive_CoreIPSubsystem system (
    .clock(system_clock),
    .reset(system_reset),
    .halt_from_tile_0(system_halt_from_tile_0),
    .wfi_from_tile_0(system_wfi_from_tile_0),
    .cease_from_tile_0(system_cease_from_tile_0),
    .psd_test_clock_enable(system_psd_test_clock_enable),
    .meip_0(system_meip_0),
    .resetctrl_hartIsInReset_0(system_resetctrl_hartIsInReset_0),
    .debug_clock(system_debug_clock),
    .debug_reset(system_debug_reset),
    .debug_systemjtag_jtag_TCK(system_debug_systemjtag_jtag_TCK),
    .debug_systemjtag_jtag_TMS(system_debug_systemjtag_jtag_TMS),
    .debug_systemjtag_jtag_TDI(system_debug_systemjtag_jtag_TDI),
    .debug_systemjtag_jtag_TDO_data(system_debug_systemjtag_jtag_TDO_data),
    .debug_systemjtag_jtag_TDO_driven(system_debug_systemjtag_jtag_TDO_driven),
    .debug_systemjtag_reset(system_debug_systemjtag_reset),
    .debug_systemjtag_mfr_id(system_debug_systemjtag_mfr_id),
    .debug_systemjtag_part_number(system_debug_systemjtag_part_number),
    .debug_systemjtag_version(system_debug_systemjtag_version),
    .debug_ndreset(system_debug_ndreset),
    .debug_dmactive(system_debug_dmactive),
    .debug_dmactiveAck(system_debug_dmactiveAck),
    .reset_vector_0(system_reset_vector_0),
    .rtc_toggle(system_rtc_toggle),
    .local_interrupts_0(system_local_interrupts_0),
    .sys_port_ahb_0_hmastlock(system_sys_port_ahb_0_hmastlock),
    .sys_port_ahb_0_hready(system_sys_port_ahb_0_hready),
    .sys_port_ahb_0_htrans(system_sys_port_ahb_0_htrans),
    .sys_port_ahb_0_hsize(system_sys_port_ahb_0_hsize),
    .sys_port_ahb_0_hburst(system_sys_port_ahb_0_hburst),
    .sys_port_ahb_0_hwrite(system_sys_port_ahb_0_hwrite),
    .sys_port_ahb_0_hprot(system_sys_port_ahb_0_hprot),
    .sys_port_ahb_0_haddr(system_sys_port_ahb_0_haddr),
    .sys_port_ahb_0_hwdata(system_sys_port_ahb_0_hwdata),
    .sys_port_ahb_0_hresp(system_sys_port_ahb_0_hresp),
    .sys_port_ahb_0_hrdata(system_sys_port_ahb_0_hrdata),
    .periph_port_ahb_0_hmastlock(system_periph_port_ahb_0_hmastlock),
    .periph_port_ahb_0_hready(system_periph_port_ahb_0_hready),
    .periph_port_ahb_0_htrans(system_periph_port_ahb_0_htrans),
    .periph_port_ahb_0_hsize(system_periph_port_ahb_0_hsize),
    .periph_port_ahb_0_hburst(system_periph_port_ahb_0_hburst),
    .periph_port_ahb_0_hwrite(system_periph_port_ahb_0_hwrite),
    .periph_port_ahb_0_hprot(system_periph_port_ahb_0_hprot),
    .periph_port_ahb_0_haddr(system_periph_port_ahb_0_haddr),
    .periph_port_ahb_0_hwdata(system_periph_port_ahb_0_hwdata),
    .periph_port_ahb_0_hresp(system_periph_port_ahb_0_hresp),
    .periph_port_ahb_0_hrdata(system_periph_port_ahb_0_hrdata),
    .front_port_ahb_0_hmastlock(system_front_port_ahb_0_hmastlock),
    .front_port_ahb_0_hsel(system_front_port_ahb_0_hsel),
    .front_port_ahb_0_hready(system_front_port_ahb_0_hready),
    .front_port_ahb_0_hreadyout(system_front_port_ahb_0_hreadyout),
    .front_port_ahb_0_htrans(system_front_port_ahb_0_htrans),
    .front_port_ahb_0_hsize(system_front_port_ahb_0_hsize),
    .front_port_ahb_0_hburst(system_front_port_ahb_0_hburst),
    .front_port_ahb_0_hwrite(system_front_port_ahb_0_hwrite),
    .front_port_ahb_0_hprot(system_front_port_ahb_0_hprot),
    .front_port_ahb_0_haddr(system_front_port_ahb_0_haddr),
    .front_port_ahb_0_hwdata(system_front_port_ahb_0_hwdata),
    .front_port_ahb_0_hresp(system_front_port_ahb_0_hresp),
    .front_port_ahb_0_hrdata(system_front_port_ahb_0_hrdata)
  );
  Pow2ClockDivider func_clock (
    .clock(func_clock_clock),
    .io_clock_out(func_clock_io_clock_out)
  );
  system_clock_en dpiClockGate (
    .clock_in(dpiClockGate_clock_in),
    .clock_out(dpiClockGate_clock_out)
  );
  c_core_reset_driver c_core_reset_driver (
    .clock(c_core_reset_driver_clock)
  );
  SiFive_DebugCompatibility_DebugCompatibility debug_compatibility (
    .clock(debug_compatibility_clock),
    .reset(debug_compatibility_reset),
    .debug_outer_reset(debug_compatibility_debug_outer_reset),
    .debug_clock(debug_compatibility_debug_clock),
    .debug_reset(debug_compatibility_debug_reset),
    .debug_dmactive(debug_compatibility_debug_dmactive),
    .debug_dmactiveAck(debug_compatibility_debug_dmactiveAck),
    .debug_resetctrl_hartIsInReset_0(debug_compatibility_debug_resetctrl_hartIsInReset_0)
  );
  DataTap_9 DataTap_9 (
    ._0_clock(DataTap_9__0_clock),
    ._0_reset(DataTap_9__0_reset),
    ._0_excpt(DataTap_9__0_excpt),
    ._0_priv_mode(DataTap_9__0_priv_mode),
    ._0_hartid(DataTap_9__0_hartid),
    ._0_timer(DataTap_9__0_timer),
    ._0_valid(DataTap_9__0_valid),
    ._0_pc(DataTap_9__0_pc),
    ._0_wrdst(DataTap_9__0_wrdst),
    ._0_wrdata(DataTap_9__0_wrdata),
    ._0_wrenx(DataTap_9__0_wrenx),
    ._0_wrenf(DataTap_9__0_wrenf),
    ._0_rd0src(DataTap_9__0_rd0src),
    ._0_rd0val(DataTap_9__0_rd0val),
    ._0_rd1src(DataTap_9__0_rd1src),
    ._0_rd1val(DataTap_9__0_rd1val),
    ._0_inst(DataTap_9__0_inst)
  );
  DataTap_2 DataTap_2 (
    ._10(DataTap_2__10),
    ._9(DataTap_2__9),
    ._8(DataTap_2__8),
    ._7(DataTap_2__7),
    ._6(DataTap_2__6),
    ._5(DataTap_2__5),
    ._4(DataTap_2__4),
    ._3(DataTap_2__3),
    ._2(DataTap_2__2),
    ._1(DataTap_2__1),
    ._0(DataTap_2__0)
  );
  AHBPortRAMSlave testRAM (
    .clock(testRAM_clock),
    .reset(testRAM_reset),
    .io_ahb_0_hready(testRAM_io_ahb_0_hready),
    .io_ahb_0_htrans(testRAM_io_ahb_0_htrans),
    .io_ahb_0_hsize(testRAM_io_ahb_0_hsize),
    .io_ahb_0_hwrite(testRAM_io_ahb_0_hwrite),
    .io_ahb_0_haddr(testRAM_io_ahb_0_haddr),
    .io_ahb_0_hwdata(testRAM_io_ahb_0_hwdata),
    .io_ahb_0_hresp(testRAM_io_ahb_0_hresp),
    .io_ahb_0_hrdata(testRAM_io_ahb_0_hrdata)
  );
  AHBPortRAMSlave_1 testRAM_1 (
    .clock(testRAM_1_clock),
    .reset(testRAM_1_reset),
    .io_ahb_0_hready(testRAM_1_io_ahb_0_hready),
    .io_ahb_0_htrans(testRAM_1_io_ahb_0_htrans),
    .io_ahb_0_hsize(testRAM_1_io_ahb_0_hsize),
    .io_ahb_0_hwrite(testRAM_1_io_ahb_0_hwrite),
    .io_ahb_0_haddr(testRAM_1_io_ahb_0_haddr),
    .io_ahb_0_hwdata(testRAM_1_io_ahb_0_hwdata),
    .io_ahb_0_hresp(testRAM_1_io_ahb_0_hresp),
    .io_ahb_0_hrdata(testRAM_1_io_ahb_0_hrdata)
  );
  WfiChecker #(.PCWIDTH(32)) WfiChecker (
    .reset(WfiChecker_reset),
    .clock(WfiChecker_clock),
    .wfi(WfiChecker_wfi),
    .excpt(WfiChecker_excpt),
    .bus_err_int(WfiChecker_bus_err_int),
    .debug_int(WfiChecker_debug_int),
    .clint_int(WfiChecker_clint_int),
    .allow_wfi(WfiChecker_allow_wfi),
    .debug(WfiChecker_debug),
    .singleStep(WfiChecker_singleStep),
    .reg_mie(WfiChecker_reg_mie),
    .reg_mip(WfiChecker_reg_mip),
    .inst_vld_0(WfiChecker_inst_vld_0),
    .pc_0(WfiChecker_pc_0),
    .inst_0(WfiChecker_inst_0)
  );
  core_monitor core_monitor (
    .m_0_clock(core_monitor_m_0_clock),
    .m_0_reset(core_monitor_m_0_reset),
    .m_0_excpt(core_monitor_m_0_excpt),
    .m_0_priv_mode(core_monitor_m_0_priv_mode),
    .m_0_hartid(core_monitor_m_0_hartid),
    .m_0_timer(core_monitor_m_0_timer),
    .m_0_valid(core_monitor_m_0_valid),
    .m_0_pc(core_monitor_m_0_pc),
    .m_0_wrdst(core_monitor_m_0_wrdst),
    .m_0_wrdata(core_monitor_m_0_wrdata),
    .m_0_wrenx(core_monitor_m_0_wrenx),
    .m_0_wrenf(core_monitor_m_0_wrenf),
    .m_0_rd0src(core_monitor_m_0_rd0src),
    .m_0_rd0val(core_monitor_m_0_rd0val),
    .m_0_rd1src(core_monitor_m_0_rd1src),
    .m_0_rd1val(core_monitor_m_0_rd1val),
    .m_0_inst(core_monitor_m_0_inst)
  );
  DPITestbenchHooks dpitbh (
    .clock(dpitbh_clock),
    .reset(dpitbh_reset)
  );
  plusarg_reader #(.FORMAT("drive_global_interrupt_type=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  GlobalIntDriver GlobalIntDriver (
    .clock(GlobalIntDriver_clock),
    .reset(GlobalIntDriver_reset)
  );
  plusarg_reader #(.FORMAT("drive_local_interrupt_type=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 (
    .out(plusarg_reader_1_out)
  );
  NullInterruptDriver #(.ID(0), .WIDTH(127)) NullInterruptDriver (
    .clock(NullInterruptDriver_clock),
    .reset(NullInterruptDriver_reset),
    .interrupts(NullInterruptDriver_interrupts)
  );
  assign _T_5 = _T_2 + 5'h1;
  assign _T_6 = _T_2 == 5'h0;
  assign _T_7 = ~_T_3;
  assign _T_13 = system_reset;
  assign _T_30 = plusarg_reader_out;
  assign _T_34 = _T_30 == 32'h0;
  assign _T_35 = _T_30 == 32'h1;
  assign _T_36 = _T_30 == 32'h2;
  assign _T_37 = _T_30 == 32'h3;
  assign _T_38 = _T_30 == 32'h4;
  assign _T_41 = ~reset;
  assign _T_43 = value_1 == 7'h63;
  assign _T_45 = value_1 + 7'h1;
  assign _T_42 = plusarg_reader_1_out;
  assign _T_46 = _T_42 == 32'h0;
  assign _T_47 = _T_42 == 32'h1;
  assign _T_49 = _T_42 == 32'h2;
  assign _T_177 = _T_42 == 32'h3;
  assign _T_179 = value_2 == 7'h7e;
  assign _T_181 = value_2 + 7'h1;
  assign _T_182 = 128'h1 << value_2;
  assign _T_183 = _T_42 == 32'h4;
  assign _T_185 = _T_184 == 16'h0;
  assign _T_188 = _T_184[0] ^ _T_184[2];
  assign _T_190 = _T_188 ^ _T_184[3];
  assign _T_192 = _T_190 ^ _T_184[5];
  assign _T_194 = {_T_192,_T_184[15:1]};
  assign _T_197 = _T_196 == 16'h0;
  assign _T_200 = _T_196[0] ^ _T_196[2];
  assign _T_202 = _T_200 ^ _T_196[3];
  assign _T_204 = _T_202 ^ _T_196[5];
  assign _T_206 = {_T_204,_T_196[15:1]};
  assign _T_209 = _T_208 == 16'h0;
  assign _T_212 = _T_208[0] ^ _T_208[2];
  assign _T_214 = _T_212 ^ _T_208[3];
  assign _T_216 = _T_214 ^ _T_208[5];
  assign _T_218 = {_T_216,_T_208[15:1]};
  assign _T_221 = _T_220 == 16'h0;
  assign _T_224 = _T_220[0] ^ _T_220[2];
  assign _T_226 = _T_224 ^ _T_220[3];
  assign _T_228 = _T_226 ^ _T_220[5];
  assign _T_230 = {_T_228,_T_220[15:1]};
  assign _T_233 = _T_232 == 16'h0;
  assign _T_236 = _T_232[0] ^ _T_232[2];
  assign _T_238 = _T_236 ^ _T_232[3];
  assign _T_240 = _T_238 ^ _T_232[5];
  assign _T_242 = {_T_240,_T_232[15:1]};
  assign _T_245 = _T_244 == 16'h0;
  assign _T_248 = _T_244[0] ^ _T_244[2];
  assign _T_250 = _T_248 ^ _T_244[3];
  assign _T_252 = _T_250 ^ _T_244[5];
  assign _T_254 = {_T_252,_T_244[15:1]};
  assign _T_257 = _T_256 == 16'h0;
  assign _T_260 = _T_256[0] ^ _T_256[2];
  assign _T_262 = _T_260 ^ _T_256[3];
  assign _T_264 = _T_262 ^ _T_256[5];
  assign _T_266 = {_T_264,_T_256[15:1]};
  assign _T_269 = _T_268 == 16'h0;
  assign _T_272 = _T_268[0] ^ _T_268[2];
  assign _T_274 = _T_272 ^ _T_268[3];
  assign _T_276 = _T_274 ^ _T_268[5];
  assign _T_278 = {_T_276,_T_268[15:1]};
  assign _T_281 = _T_280 == 16'h0;
  assign _T_284 = _T_280[0] ^ _T_280[2];
  assign _T_286 = _T_284 ^ _T_280[3];
  assign _T_288 = _T_286 ^ _T_280[5];
  assign _T_290 = {_T_288,_T_280[15:1]};
  assign _T_293 = _T_292 == 16'h0;
  assign _T_296 = _T_292[0] ^ _T_292[2];
  assign _T_298 = _T_296 ^ _T_292[3];
  assign _T_300 = _T_298 ^ _T_292[5];
  assign _T_302 = {_T_300,_T_292[15:1]};
  assign _T_305 = _T_304 == 16'h0;
  assign _T_308 = _T_304[0] ^ _T_304[2];
  assign _T_310 = _T_308 ^ _T_304[3];
  assign _T_312 = _T_310 ^ _T_304[5];
  assign _T_314 = {_T_312,_T_304[15:1]};
  assign _T_317 = _T_316 == 16'h0;
  assign _T_320 = _T_316[0] ^ _T_316[2];
  assign _T_322 = _T_320 ^ _T_316[3];
  assign _T_324 = _T_322 ^ _T_316[5];
  assign _T_326 = {_T_324,_T_316[15:1]};
  assign _T_329 = _T_328 == 16'h0;
  assign _T_332 = _T_328[0] ^ _T_328[2];
  assign _T_334 = _T_332 ^ _T_328[3];
  assign _T_336 = _T_334 ^ _T_328[5];
  assign _T_338 = {_T_336,_T_328[15:1]};
  assign _T_341 = _T_340 == 16'h0;
  assign _T_344 = _T_340[0] ^ _T_340[2];
  assign _T_346 = _T_344 ^ _T_340[3];
  assign _T_348 = _T_346 ^ _T_340[5];
  assign _T_350 = {_T_348,_T_340[15:1]};
  assign _T_353 = _T_352 == 16'h0;
  assign _T_356 = _T_352[0] ^ _T_352[2];
  assign _T_358 = _T_356 ^ _T_352[3];
  assign _T_360 = _T_358 ^ _T_352[5];
  assign _T_362 = {_T_360,_T_352[15:1]};
  assign _T_365 = _T_364 == 16'h0;
  assign _T_368 = _T_364[0] ^ _T_364[2];
  assign _T_370 = _T_368 ^ _T_364[3];
  assign _T_372 = _T_370 ^ _T_364[5];
  assign _T_374 = {_T_372,_T_364[15:1]};
  assign _T_377 = _T_376 == 16'h0;
  assign _T_380 = _T_376[0] ^ _T_376[2];
  assign _T_382 = _T_380 ^ _T_376[3];
  assign _T_384 = _T_382 ^ _T_376[5];
  assign _T_386 = {_T_384,_T_376[15:1]};
  assign _T_389 = _T_388 == 16'h0;
  assign _T_392 = _T_388[0] ^ _T_388[2];
  assign _T_394 = _T_392 ^ _T_388[3];
  assign _T_396 = _T_394 ^ _T_388[5];
  assign _T_398 = {_T_396,_T_388[15:1]};
  assign _T_401 = _T_400 == 16'h0;
  assign _T_404 = _T_400[0] ^ _T_400[2];
  assign _T_406 = _T_404 ^ _T_400[3];
  assign _T_408 = _T_406 ^ _T_400[5];
  assign _T_410 = {_T_408,_T_400[15:1]};
  assign _T_413 = _T_412 == 16'h0;
  assign _T_416 = _T_412[0] ^ _T_412[2];
  assign _T_418 = _T_416 ^ _T_412[3];
  assign _T_420 = _T_418 ^ _T_412[5];
  assign _T_422 = {_T_420,_T_412[15:1]};
  assign _T_425 = _T_424 == 16'h0;
  assign _T_428 = _T_424[0] ^ _T_424[2];
  assign _T_430 = _T_428 ^ _T_424[3];
  assign _T_432 = _T_430 ^ _T_424[5];
  assign _T_434 = {_T_432,_T_424[15:1]};
  assign _T_437 = _T_436 == 16'h0;
  assign _T_440 = _T_436[0] ^ _T_436[2];
  assign _T_442 = _T_440 ^ _T_436[3];
  assign _T_444 = _T_442 ^ _T_436[5];
  assign _T_446 = {_T_444,_T_436[15:1]};
  assign _T_449 = _T_448 == 16'h0;
  assign _T_452 = _T_448[0] ^ _T_448[2];
  assign _T_454 = _T_452 ^ _T_448[3];
  assign _T_456 = _T_454 ^ _T_448[5];
  assign _T_458 = {_T_456,_T_448[15:1]};
  assign _T_461 = _T_460 == 16'h0;
  assign _T_464 = _T_460[0] ^ _T_460[2];
  assign _T_466 = _T_464 ^ _T_460[3];
  assign _T_468 = _T_466 ^ _T_460[5];
  assign _T_470 = {_T_468,_T_460[15:1]};
  assign _T_473 = _T_472 == 16'h0;
  assign _T_476 = _T_472[0] ^ _T_472[2];
  assign _T_478 = _T_476 ^ _T_472[3];
  assign _T_480 = _T_478 ^ _T_472[5];
  assign _T_482 = {_T_480,_T_472[15:1]};
  assign _T_485 = _T_484 == 16'h0;
  assign _T_488 = _T_484[0] ^ _T_484[2];
  assign _T_490 = _T_488 ^ _T_484[3];
  assign _T_492 = _T_490 ^ _T_484[5];
  assign _T_494 = {_T_492,_T_484[15:1]};
  assign _T_497 = _T_496 == 16'h0;
  assign _T_500 = _T_496[0] ^ _T_496[2];
  assign _T_502 = _T_500 ^ _T_496[3];
  assign _T_504 = _T_502 ^ _T_496[5];
  assign _T_506 = {_T_504,_T_496[15:1]};
  assign _T_509 = _T_508 == 16'h0;
  assign _T_512 = _T_508[0] ^ _T_508[2];
  assign _T_514 = _T_512 ^ _T_508[3];
  assign _T_516 = _T_514 ^ _T_508[5];
  assign _T_518 = {_T_516,_T_508[15:1]};
  assign _T_521 = _T_520 == 16'h0;
  assign _T_524 = _T_520[0] ^ _T_520[2];
  assign _T_526 = _T_524 ^ _T_520[3];
  assign _T_528 = _T_526 ^ _T_520[5];
  assign _T_530 = {_T_528,_T_520[15:1]};
  assign _T_533 = _T_532 == 16'h0;
  assign _T_536 = _T_532[0] ^ _T_532[2];
  assign _T_538 = _T_536 ^ _T_532[3];
  assign _T_540 = _T_538 ^ _T_532[5];
  assign _T_542 = {_T_540,_T_532[15:1]};
  assign _T_545 = _T_544 == 16'h0;
  assign _T_548 = _T_544[0] ^ _T_544[2];
  assign _T_550 = _T_548 ^ _T_544[3];
  assign _T_552 = _T_550 ^ _T_544[5];
  assign _T_554 = {_T_552,_T_544[15:1]};
  assign _T_557 = _T_556 == 16'h0;
  assign _T_560 = _T_556[0] ^ _T_556[2];
  assign _T_562 = _T_560 ^ _T_556[3];
  assign _T_564 = _T_562 ^ _T_556[5];
  assign _T_566 = {_T_564,_T_556[15:1]};
  assign _T_569 = _T_568 == 16'h0;
  assign _T_572 = _T_568[0] ^ _T_568[2];
  assign _T_574 = _T_572 ^ _T_568[3];
  assign _T_576 = _T_574 ^ _T_568[5];
  assign _T_578 = {_T_576,_T_568[15:1]};
  assign _T_581 = _T_580 == 16'h0;
  assign _T_584 = _T_580[0] ^ _T_580[2];
  assign _T_586 = _T_584 ^ _T_580[3];
  assign _T_588 = _T_586 ^ _T_580[5];
  assign _T_590 = {_T_588,_T_580[15:1]};
  assign _T_593 = _T_592 == 16'h0;
  assign _T_596 = _T_592[0] ^ _T_592[2];
  assign _T_598 = _T_596 ^ _T_592[3];
  assign _T_600 = _T_598 ^ _T_592[5];
  assign _T_602 = {_T_600,_T_592[15:1]};
  assign _T_605 = _T_604 == 16'h0;
  assign _T_608 = _T_604[0] ^ _T_604[2];
  assign _T_610 = _T_608 ^ _T_604[3];
  assign _T_612 = _T_610 ^ _T_604[5];
  assign _T_614 = {_T_612,_T_604[15:1]};
  assign _T_617 = _T_616 == 16'h0;
  assign _T_620 = _T_616[0] ^ _T_616[2];
  assign _T_622 = _T_620 ^ _T_616[3];
  assign _T_624 = _T_622 ^ _T_616[5];
  assign _T_626 = {_T_624,_T_616[15:1]};
  assign _T_629 = _T_628 == 16'h0;
  assign _T_632 = _T_628[0] ^ _T_628[2];
  assign _T_634 = _T_632 ^ _T_628[3];
  assign _T_636 = _T_634 ^ _T_628[5];
  assign _T_638 = {_T_636,_T_628[15:1]};
  assign _T_641 = _T_640 == 16'h0;
  assign _T_644 = _T_640[0] ^ _T_640[2];
  assign _T_646 = _T_644 ^ _T_640[3];
  assign _T_648 = _T_646 ^ _T_640[5];
  assign _T_650 = {_T_648,_T_640[15:1]};
  assign _T_653 = _T_652 == 16'h0;
  assign _T_656 = _T_652[0] ^ _T_652[2];
  assign _T_658 = _T_656 ^ _T_652[3];
  assign _T_660 = _T_658 ^ _T_652[5];
  assign _T_662 = {_T_660,_T_652[15:1]};
  assign _T_665 = _T_664 == 16'h0;
  assign _T_668 = _T_664[0] ^ _T_664[2];
  assign _T_670 = _T_668 ^ _T_664[3];
  assign _T_672 = _T_670 ^ _T_664[5];
  assign _T_674 = {_T_672,_T_664[15:1]};
  assign _T_677 = _T_676 == 16'h0;
  assign _T_680 = _T_676[0] ^ _T_676[2];
  assign _T_682 = _T_680 ^ _T_676[3];
  assign _T_684 = _T_682 ^ _T_676[5];
  assign _T_686 = {_T_684,_T_676[15:1]};
  assign _T_689 = _T_688 == 16'h0;
  assign _T_692 = _T_688[0] ^ _T_688[2];
  assign _T_694 = _T_692 ^ _T_688[3];
  assign _T_696 = _T_694 ^ _T_688[5];
  assign _T_698 = {_T_696,_T_688[15:1]};
  assign _T_701 = _T_700 == 16'h0;
  assign _T_704 = _T_700[0] ^ _T_700[2];
  assign _T_706 = _T_704 ^ _T_700[3];
  assign _T_708 = _T_706 ^ _T_700[5];
  assign _T_710 = {_T_708,_T_700[15:1]};
  assign _T_713 = _T_712 == 16'h0;
  assign _T_716 = _T_712[0] ^ _T_712[2];
  assign _T_718 = _T_716 ^ _T_712[3];
  assign _T_720 = _T_718 ^ _T_712[5];
  assign _T_722 = {_T_720,_T_712[15:1]};
  assign _T_725 = _T_724 == 16'h0;
  assign _T_728 = _T_724[0] ^ _T_724[2];
  assign _T_730 = _T_728 ^ _T_724[3];
  assign _T_732 = _T_730 ^ _T_724[5];
  assign _T_734 = {_T_732,_T_724[15:1]};
  assign _T_737 = _T_736 == 16'h0;
  assign _T_740 = _T_736[0] ^ _T_736[2];
  assign _T_742 = _T_740 ^ _T_736[3];
  assign _T_744 = _T_742 ^ _T_736[5];
  assign _T_746 = {_T_744,_T_736[15:1]};
  assign _T_749 = _T_748 == 16'h0;
  assign _T_752 = _T_748[0] ^ _T_748[2];
  assign _T_754 = _T_752 ^ _T_748[3];
  assign _T_756 = _T_754 ^ _T_748[5];
  assign _T_758 = {_T_756,_T_748[15:1]};
  assign _T_761 = _T_760 == 16'h0;
  assign _T_764 = _T_760[0] ^ _T_760[2];
  assign _T_766 = _T_764 ^ _T_760[3];
  assign _T_768 = _T_766 ^ _T_760[5];
  assign _T_770 = {_T_768,_T_760[15:1]};
  assign _T_773 = _T_772 == 16'h0;
  assign _T_776 = _T_772[0] ^ _T_772[2];
  assign _T_778 = _T_776 ^ _T_772[3];
  assign _T_780 = _T_778 ^ _T_772[5];
  assign _T_782 = {_T_780,_T_772[15:1]};
  assign _T_785 = _T_784 == 16'h0;
  assign _T_788 = _T_784[0] ^ _T_784[2];
  assign _T_790 = _T_788 ^ _T_784[3];
  assign _T_792 = _T_790 ^ _T_784[5];
  assign _T_794 = {_T_792,_T_784[15:1]};
  assign _T_797 = _T_796 == 16'h0;
  assign _T_800 = _T_796[0] ^ _T_796[2];
  assign _T_802 = _T_800 ^ _T_796[3];
  assign _T_804 = _T_802 ^ _T_796[5];
  assign _T_806 = {_T_804,_T_796[15:1]};
  assign _T_809 = _T_808 == 16'h0;
  assign _T_812 = _T_808[0] ^ _T_808[2];
  assign _T_814 = _T_812 ^ _T_808[3];
  assign _T_816 = _T_814 ^ _T_808[5];
  assign _T_818 = {_T_816,_T_808[15:1]};
  assign _T_821 = _T_820 == 16'h0;
  assign _T_824 = _T_820[0] ^ _T_820[2];
  assign _T_826 = _T_824 ^ _T_820[3];
  assign _T_828 = _T_826 ^ _T_820[5];
  assign _T_830 = {_T_828,_T_820[15:1]};
  assign _T_833 = _T_832 == 16'h0;
  assign _T_836 = _T_832[0] ^ _T_832[2];
  assign _T_838 = _T_836 ^ _T_832[3];
  assign _T_840 = _T_838 ^ _T_832[5];
  assign _T_842 = {_T_840,_T_832[15:1]};
  assign _T_845 = _T_844 == 16'h0;
  assign _T_848 = _T_844[0] ^ _T_844[2];
  assign _T_850 = _T_848 ^ _T_844[3];
  assign _T_852 = _T_850 ^ _T_844[5];
  assign _T_854 = {_T_852,_T_844[15:1]};
  assign _T_857 = _T_856 == 16'h0;
  assign _T_860 = _T_856[0] ^ _T_856[2];
  assign _T_862 = _T_860 ^ _T_856[3];
  assign _T_864 = _T_862 ^ _T_856[5];
  assign _T_866 = {_T_864,_T_856[15:1]};
  assign _T_869 = _T_868 == 16'h0;
  assign _T_872 = _T_868[0] ^ _T_868[2];
  assign _T_874 = _T_872 ^ _T_868[3];
  assign _T_876 = _T_874 ^ _T_868[5];
  assign _T_878 = {_T_876,_T_868[15:1]};
  assign _T_881 = _T_880 == 16'h0;
  assign _T_884 = _T_880[0] ^ _T_880[2];
  assign _T_886 = _T_884 ^ _T_880[3];
  assign _T_888 = _T_886 ^ _T_880[5];
  assign _T_890 = {_T_888,_T_880[15:1]};
  assign _T_893 = _T_892 == 16'h0;
  assign _T_896 = _T_892[0] ^ _T_892[2];
  assign _T_898 = _T_896 ^ _T_892[3];
  assign _T_900 = _T_898 ^ _T_892[5];
  assign _T_902 = {_T_900,_T_892[15:1]};
  assign _T_905 = _T_904 == 16'h0;
  assign _T_908 = _T_904[0] ^ _T_904[2];
  assign _T_910 = _T_908 ^ _T_904[3];
  assign _T_912 = _T_910 ^ _T_904[5];
  assign _T_914 = {_T_912,_T_904[15:1]};
  assign _T_917 = _T_916 == 16'h0;
  assign _T_920 = _T_916[0] ^ _T_916[2];
  assign _T_922 = _T_920 ^ _T_916[3];
  assign _T_924 = _T_922 ^ _T_916[5];
  assign _T_926 = {_T_924,_T_916[15:1]};
  assign _T_929 = _T_928 == 16'h0;
  assign _T_932 = _T_928[0] ^ _T_928[2];
  assign _T_934 = _T_932 ^ _T_928[3];
  assign _T_936 = _T_934 ^ _T_928[5];
  assign _T_938 = {_T_936,_T_928[15:1]};
  assign _T_941 = _T_940 == 16'h0;
  assign _T_944 = _T_940[0] ^ _T_940[2];
  assign _T_946 = _T_944 ^ _T_940[3];
  assign _T_948 = _T_946 ^ _T_940[5];
  assign _T_950 = {_T_948,_T_940[15:1]};
  assign _T_953 = _T_952 == 16'h0;
  assign _T_956 = _T_952[0] ^ _T_952[2];
  assign _T_958 = _T_956 ^ _T_952[3];
  assign _T_960 = _T_958 ^ _T_952[5];
  assign _T_962 = {_T_960,_T_952[15:1]};
  assign _T_965 = _T_964 == 16'h0;
  assign _T_968 = _T_964[0] ^ _T_964[2];
  assign _T_970 = _T_968 ^ _T_964[3];
  assign _T_972 = _T_970 ^ _T_964[5];
  assign _T_974 = {_T_972,_T_964[15:1]};
  assign _T_977 = _T_976 == 16'h0;
  assign _T_980 = _T_976[0] ^ _T_976[2];
  assign _T_982 = _T_980 ^ _T_976[3];
  assign _T_984 = _T_982 ^ _T_976[5];
  assign _T_986 = {_T_984,_T_976[15:1]};
  assign _T_989 = _T_988 == 16'h0;
  assign _T_992 = _T_988[0] ^ _T_988[2];
  assign _T_994 = _T_992 ^ _T_988[3];
  assign _T_996 = _T_994 ^ _T_988[5];
  assign _T_998 = {_T_996,_T_988[15:1]};
  assign _T_1001 = _T_1000 == 16'h0;
  assign _T_1004 = _T_1000[0] ^ _T_1000[2];
  assign _T_1006 = _T_1004 ^ _T_1000[3];
  assign _T_1008 = _T_1006 ^ _T_1000[5];
  assign _T_1010 = {_T_1008,_T_1000[15:1]};
  assign _T_1013 = _T_1012 == 16'h0;
  assign _T_1016 = _T_1012[0] ^ _T_1012[2];
  assign _T_1018 = _T_1016 ^ _T_1012[3];
  assign _T_1020 = _T_1018 ^ _T_1012[5];
  assign _T_1022 = {_T_1020,_T_1012[15:1]};
  assign _T_1025 = _T_1024 == 16'h0;
  assign _T_1028 = _T_1024[0] ^ _T_1024[2];
  assign _T_1030 = _T_1028 ^ _T_1024[3];
  assign _T_1032 = _T_1030 ^ _T_1024[5];
  assign _T_1034 = {_T_1032,_T_1024[15:1]};
  assign _T_1037 = _T_1036 == 16'h0;
  assign _T_1040 = _T_1036[0] ^ _T_1036[2];
  assign _T_1042 = _T_1040 ^ _T_1036[3];
  assign _T_1044 = _T_1042 ^ _T_1036[5];
  assign _T_1046 = {_T_1044,_T_1036[15:1]};
  assign _T_1049 = _T_1048 == 16'h0;
  assign _T_1052 = _T_1048[0] ^ _T_1048[2];
  assign _T_1054 = _T_1052 ^ _T_1048[3];
  assign _T_1056 = _T_1054 ^ _T_1048[5];
  assign _T_1058 = {_T_1056,_T_1048[15:1]};
  assign _T_1061 = _T_1060 == 16'h0;
  assign _T_1064 = _T_1060[0] ^ _T_1060[2];
  assign _T_1066 = _T_1064 ^ _T_1060[3];
  assign _T_1068 = _T_1066 ^ _T_1060[5];
  assign _T_1070 = {_T_1068,_T_1060[15:1]};
  assign _T_1073 = _T_1072 == 16'h0;
  assign _T_1076 = _T_1072[0] ^ _T_1072[2];
  assign _T_1078 = _T_1076 ^ _T_1072[3];
  assign _T_1080 = _T_1078 ^ _T_1072[5];
  assign _T_1082 = {_T_1080,_T_1072[15:1]};
  assign _T_1085 = _T_1084 == 16'h0;
  assign _T_1088 = _T_1084[0] ^ _T_1084[2];
  assign _T_1090 = _T_1088 ^ _T_1084[3];
  assign _T_1092 = _T_1090 ^ _T_1084[5];
  assign _T_1094 = {_T_1092,_T_1084[15:1]};
  assign _T_1097 = _T_1096 == 16'h0;
  assign _T_1100 = _T_1096[0] ^ _T_1096[2];
  assign _T_1102 = _T_1100 ^ _T_1096[3];
  assign _T_1104 = _T_1102 ^ _T_1096[5];
  assign _T_1106 = {_T_1104,_T_1096[15:1]};
  assign _T_1109 = _T_1108 == 16'h0;
  assign _T_1112 = _T_1108[0] ^ _T_1108[2];
  assign _T_1114 = _T_1112 ^ _T_1108[3];
  assign _T_1116 = _T_1114 ^ _T_1108[5];
  assign _T_1118 = {_T_1116,_T_1108[15:1]};
  assign _T_1121 = _T_1120 == 16'h0;
  assign _T_1124 = _T_1120[0] ^ _T_1120[2];
  assign _T_1126 = _T_1124 ^ _T_1120[3];
  assign _T_1128 = _T_1126 ^ _T_1120[5];
  assign _T_1130 = {_T_1128,_T_1120[15:1]};
  assign _T_1133 = _T_1132 == 16'h0;
  assign _T_1136 = _T_1132[0] ^ _T_1132[2];
  assign _T_1138 = _T_1136 ^ _T_1132[3];
  assign _T_1140 = _T_1138 ^ _T_1132[5];
  assign _T_1142 = {_T_1140,_T_1132[15:1]};
  assign _T_1145 = _T_1144 == 16'h0;
  assign _T_1148 = _T_1144[0] ^ _T_1144[2];
  assign _T_1150 = _T_1148 ^ _T_1144[3];
  assign _T_1152 = _T_1150 ^ _T_1144[5];
  assign _T_1154 = {_T_1152,_T_1144[15:1]};
  assign _T_1157 = _T_1156 == 16'h0;
  assign _T_1160 = _T_1156[0] ^ _T_1156[2];
  assign _T_1162 = _T_1160 ^ _T_1156[3];
  assign _T_1164 = _T_1162 ^ _T_1156[5];
  assign _T_1166 = {_T_1164,_T_1156[15:1]};
  assign _T_1169 = _T_1168 == 16'h0;
  assign _T_1172 = _T_1168[0] ^ _T_1168[2];
  assign _T_1174 = _T_1172 ^ _T_1168[3];
  assign _T_1176 = _T_1174 ^ _T_1168[5];
  assign _T_1178 = {_T_1176,_T_1168[15:1]};
  assign _T_1181 = _T_1180 == 16'h0;
  assign _T_1184 = _T_1180[0] ^ _T_1180[2];
  assign _T_1186 = _T_1184 ^ _T_1180[3];
  assign _T_1188 = _T_1186 ^ _T_1180[5];
  assign _T_1190 = {_T_1188,_T_1180[15:1]};
  assign _T_1193 = _T_1192 == 16'h0;
  assign _T_1196 = _T_1192[0] ^ _T_1192[2];
  assign _T_1198 = _T_1196 ^ _T_1192[3];
  assign _T_1200 = _T_1198 ^ _T_1192[5];
  assign _T_1202 = {_T_1200,_T_1192[15:1]};
  assign _T_1205 = _T_1204 == 16'h0;
  assign _T_1208 = _T_1204[0] ^ _T_1204[2];
  assign _T_1210 = _T_1208 ^ _T_1204[3];
  assign _T_1212 = _T_1210 ^ _T_1204[5];
  assign _T_1214 = {_T_1212,_T_1204[15:1]};
  assign _T_1217 = _T_1216 == 16'h0;
  assign _T_1220 = _T_1216[0] ^ _T_1216[2];
  assign _T_1222 = _T_1220 ^ _T_1216[3];
  assign _T_1224 = _T_1222 ^ _T_1216[5];
  assign _T_1226 = {_T_1224,_T_1216[15:1]};
  assign _T_1229 = _T_1228 == 16'h0;
  assign _T_1232 = _T_1228[0] ^ _T_1228[2];
  assign _T_1234 = _T_1232 ^ _T_1228[3];
  assign _T_1236 = _T_1234 ^ _T_1228[5];
  assign _T_1238 = {_T_1236,_T_1228[15:1]};
  assign _T_1241 = _T_1240 == 16'h0;
  assign _T_1244 = _T_1240[0] ^ _T_1240[2];
  assign _T_1246 = _T_1244 ^ _T_1240[3];
  assign _T_1248 = _T_1246 ^ _T_1240[5];
  assign _T_1250 = {_T_1248,_T_1240[15:1]};
  assign _T_1253 = _T_1252 == 16'h0;
  assign _T_1256 = _T_1252[0] ^ _T_1252[2];
  assign _T_1258 = _T_1256 ^ _T_1252[3];
  assign _T_1260 = _T_1258 ^ _T_1252[5];
  assign _T_1262 = {_T_1260,_T_1252[15:1]};
  assign _T_1265 = _T_1264 == 16'h0;
  assign _T_1268 = _T_1264[0] ^ _T_1264[2];
  assign _T_1270 = _T_1268 ^ _T_1264[3];
  assign _T_1272 = _T_1270 ^ _T_1264[5];
  assign _T_1274 = {_T_1272,_T_1264[15:1]};
  assign _T_1277 = _T_1276 == 16'h0;
  assign _T_1280 = _T_1276[0] ^ _T_1276[2];
  assign _T_1282 = _T_1280 ^ _T_1276[3];
  assign _T_1284 = _T_1282 ^ _T_1276[5];
  assign _T_1286 = {_T_1284,_T_1276[15:1]};
  assign _T_1289 = _T_1288 == 16'h0;
  assign _T_1292 = _T_1288[0] ^ _T_1288[2];
  assign _T_1294 = _T_1292 ^ _T_1288[3];
  assign _T_1296 = _T_1294 ^ _T_1288[5];
  assign _T_1298 = {_T_1296,_T_1288[15:1]};
  assign _T_1301 = _T_1300 == 16'h0;
  assign _T_1304 = _T_1300[0] ^ _T_1300[2];
  assign _T_1306 = _T_1304 ^ _T_1300[3];
  assign _T_1308 = _T_1306 ^ _T_1300[5];
  assign _T_1310 = {_T_1308,_T_1300[15:1]};
  assign _T_1313 = _T_1312 == 16'h0;
  assign _T_1316 = _T_1312[0] ^ _T_1312[2];
  assign _T_1318 = _T_1316 ^ _T_1312[3];
  assign _T_1320 = _T_1318 ^ _T_1312[5];
  assign _T_1322 = {_T_1320,_T_1312[15:1]};
  assign _T_1325 = _T_1324 == 16'h0;
  assign _T_1328 = _T_1324[0] ^ _T_1324[2];
  assign _T_1330 = _T_1328 ^ _T_1324[3];
  assign _T_1332 = _T_1330 ^ _T_1324[5];
  assign _T_1334 = {_T_1332,_T_1324[15:1]};
  assign _T_1337 = _T_1336 == 16'h0;
  assign _T_1340 = _T_1336[0] ^ _T_1336[2];
  assign _T_1342 = _T_1340 ^ _T_1336[3];
  assign _T_1344 = _T_1342 ^ _T_1336[5];
  assign _T_1346 = {_T_1344,_T_1336[15:1]};
  assign _T_1349 = _T_1348 == 16'h0;
  assign _T_1352 = _T_1348[0] ^ _T_1348[2];
  assign _T_1354 = _T_1352 ^ _T_1348[3];
  assign _T_1356 = _T_1354 ^ _T_1348[5];
  assign _T_1358 = {_T_1356,_T_1348[15:1]};
  assign _T_1361 = _T_1360 == 16'h0;
  assign _T_1364 = _T_1360[0] ^ _T_1360[2];
  assign _T_1366 = _T_1364 ^ _T_1360[3];
  assign _T_1368 = _T_1366 ^ _T_1360[5];
  assign _T_1370 = {_T_1368,_T_1360[15:1]};
  assign _T_1373 = _T_1372 == 16'h0;
  assign _T_1376 = _T_1372[0] ^ _T_1372[2];
  assign _T_1378 = _T_1376 ^ _T_1372[3];
  assign _T_1380 = _T_1378 ^ _T_1372[5];
  assign _T_1382 = {_T_1380,_T_1372[15:1]};
  assign _T_1385 = _T_1384 == 16'h0;
  assign _T_1388 = _T_1384[0] ^ _T_1384[2];
  assign _T_1390 = _T_1388 ^ _T_1384[3];
  assign _T_1392 = _T_1390 ^ _T_1384[5];
  assign _T_1394 = {_T_1392,_T_1384[15:1]};
  assign _T_1397 = _T_1396 == 16'h0;
  assign _T_1400 = _T_1396[0] ^ _T_1396[2];
  assign _T_1402 = _T_1400 ^ _T_1396[3];
  assign _T_1404 = _T_1402 ^ _T_1396[5];
  assign _T_1406 = {_T_1404,_T_1396[15:1]};
  assign _T_1409 = _T_1408 == 16'h0;
  assign _T_1412 = _T_1408[0] ^ _T_1408[2];
  assign _T_1414 = _T_1412 ^ _T_1408[3];
  assign _T_1416 = _T_1414 ^ _T_1408[5];
  assign _T_1418 = {_T_1416,_T_1408[15:1]};
  assign _T_1421 = _T_1420 == 16'h0;
  assign _T_1424 = _T_1420[0] ^ _T_1420[2];
  assign _T_1426 = _T_1424 ^ _T_1420[3];
  assign _T_1428 = _T_1426 ^ _T_1420[5];
  assign _T_1430 = {_T_1428,_T_1420[15:1]};
  assign _T_1433 = _T_1432 == 16'h0;
  assign _T_1436 = _T_1432[0] ^ _T_1432[2];
  assign _T_1438 = _T_1436 ^ _T_1432[3];
  assign _T_1440 = _T_1438 ^ _T_1432[5];
  assign _T_1442 = {_T_1440,_T_1432[15:1]};
  assign _T_1445 = _T_1444 == 16'h0;
  assign _T_1448 = _T_1444[0] ^ _T_1444[2];
  assign _T_1450 = _T_1448 ^ _T_1444[3];
  assign _T_1452 = _T_1450 ^ _T_1444[5];
  assign _T_1454 = {_T_1452,_T_1444[15:1]};
  assign _T_1457 = _T_1456 == 16'h0;
  assign _T_1460 = _T_1456[0] ^ _T_1456[2];
  assign _T_1462 = _T_1460 ^ _T_1456[3];
  assign _T_1464 = _T_1462 ^ _T_1456[5];
  assign _T_1466 = {_T_1464,_T_1456[15:1]};
  assign _T_1469 = _T_1468 == 16'h0;
  assign _T_1472 = _T_1468[0] ^ _T_1468[2];
  assign _T_1474 = _T_1472 ^ _T_1468[3];
  assign _T_1476 = _T_1474 ^ _T_1468[5];
  assign _T_1478 = {_T_1476,_T_1468[15:1]};
  assign _T_1481 = _T_1480 == 16'h0;
  assign _T_1484 = _T_1480[0] ^ _T_1480[2];
  assign _T_1486 = _T_1484 ^ _T_1480[3];
  assign _T_1488 = _T_1486 ^ _T_1480[5];
  assign _T_1490 = {_T_1488,_T_1480[15:1]};
  assign _T_1493 = _T_1492 == 16'h0;
  assign _T_1496 = _T_1492[0] ^ _T_1492[2];
  assign _T_1498 = _T_1496 ^ _T_1492[3];
  assign _T_1500 = _T_1498 ^ _T_1492[5];
  assign _T_1502 = {_T_1500,_T_1492[15:1]};
  assign _T_1505 = _T_1504 == 16'h0;
  assign _T_1508 = _T_1504[0] ^ _T_1504[2];
  assign _T_1510 = _T_1508 ^ _T_1504[3];
  assign _T_1512 = _T_1510 ^ _T_1504[5];
  assign _T_1514 = {_T_1512,_T_1504[15:1]};
  assign _T_1517 = _T_1516 == 16'h0;
  assign _T_1520 = _T_1516[0] ^ _T_1516[2];
  assign _T_1522 = _T_1520 ^ _T_1516[3];
  assign _T_1524 = _T_1522 ^ _T_1516[5];
  assign _T_1526 = {_T_1524,_T_1516[15:1]};
  assign _T_1529 = _T_1528 == 16'h0;
  assign _T_1532 = _T_1528[0] ^ _T_1528[2];
  assign _T_1534 = _T_1532 ^ _T_1528[3];
  assign _T_1536 = _T_1534 ^ _T_1528[5];
  assign _T_1538 = {_T_1536,_T_1528[15:1]};
  assign _T_1541 = _T_1540 == 16'h0;
  assign _T_1544 = _T_1540[0] ^ _T_1540[2];
  assign _T_1546 = _T_1544 ^ _T_1540[3];
  assign _T_1548 = _T_1546 ^ _T_1540[5];
  assign _T_1550 = {_T_1548,_T_1540[15:1]};
  assign _T_1553 = _T_1552 == 16'h0;
  assign _T_1556 = _T_1552[0] ^ _T_1552[2];
  assign _T_1558 = _T_1556 ^ _T_1552[3];
  assign _T_1560 = _T_1558 ^ _T_1552[5];
  assign _T_1562 = {_T_1560,_T_1552[15:1]};
  assign _T_1565 = _T_1564 == 16'h0;
  assign _T_1568 = _T_1564[0] ^ _T_1564[2];
  assign _T_1570 = _T_1568 ^ _T_1564[3];
  assign _T_1572 = _T_1570 ^ _T_1564[5];
  assign _T_1574 = {_T_1572,_T_1564[15:1]};
  assign _T_1577 = _T_1576 == 16'h0;
  assign _T_1580 = _T_1576[0] ^ _T_1576[2];
  assign _T_1582 = _T_1580 ^ _T_1576[3];
  assign _T_1584 = _T_1582 ^ _T_1576[5];
  assign _T_1586 = {_T_1584,_T_1576[15:1]};
  assign _T_1589 = _T_1588 == 16'h0;
  assign _T_1592 = _T_1588[0] ^ _T_1588[2];
  assign _T_1594 = _T_1592 ^ _T_1588[3];
  assign _T_1596 = _T_1594 ^ _T_1588[5];
  assign _T_1598 = {_T_1596,_T_1588[15:1]};
  assign _T_1601 = _T_1600 == 16'h0;
  assign _T_1604 = _T_1600[0] ^ _T_1600[2];
  assign _T_1606 = _T_1604 ^ _T_1600[3];
  assign _T_1608 = _T_1606 ^ _T_1600[5];
  assign _T_1610 = {_T_1608,_T_1600[15:1]};
  assign _T_1613 = _T_1612 == 16'h0;
  assign _T_1616 = _T_1612[0] ^ _T_1612[2];
  assign _T_1618 = _T_1616 ^ _T_1612[3];
  assign _T_1620 = _T_1618 ^ _T_1612[5];
  assign _T_1622 = {_T_1620,_T_1612[15:1]};
  assign _T_1625 = _T_1624 == 16'h0;
  assign _T_1628 = _T_1624[0] ^ _T_1624[2];
  assign _T_1630 = _T_1628 ^ _T_1624[3];
  assign _T_1632 = _T_1630 ^ _T_1624[5];
  assign _T_1634 = {_T_1632,_T_1624[15:1]};
  assign _T_1637 = _T_1636 == 16'h0;
  assign _T_1640 = _T_1636[0] ^ _T_1636[2];
  assign _T_1642 = _T_1640 ^ _T_1636[3];
  assign _T_1644 = _T_1642 ^ _T_1636[5];
  assign _T_1646 = {_T_1644,_T_1636[15:1]};
  assign _T_1649 = _T_1648 == 16'h0;
  assign _T_1652 = _T_1648[0] ^ _T_1648[2];
  assign _T_1654 = _T_1652 ^ _T_1648[3];
  assign _T_1656 = _T_1654 ^ _T_1648[5];
  assign _T_1658 = {_T_1656,_T_1648[15:1]};
  assign _T_1661 = _T_1660 == 16'h0;
  assign _T_1664 = _T_1660[0] ^ _T_1660[2];
  assign _T_1666 = _T_1664 ^ _T_1660[3];
  assign _T_1668 = _T_1666 ^ _T_1660[5];
  assign _T_1670 = {_T_1668,_T_1660[15:1]};
  assign _T_1673 = _T_1672 == 16'h0;
  assign _T_1676 = _T_1672[0] ^ _T_1672[2];
  assign _T_1678 = _T_1676 ^ _T_1672[3];
  assign _T_1680 = _T_1678 ^ _T_1672[5];
  assign _T_1682 = {_T_1680,_T_1672[15:1]};
  assign _T_1685 = _T_1684 == 16'h0;
  assign _T_1688 = _T_1684[0] ^ _T_1684[2];
  assign _T_1690 = _T_1688 ^ _T_1684[3];
  assign _T_1692 = _T_1690 ^ _T_1684[5];
  assign _T_1694 = {_T_1692,_T_1684[15:1]};
  assign _T_1697 = _T_1696 == 16'h0;
  assign _T_1700 = _T_1696[0] ^ _T_1696[2];
  assign _T_1702 = _T_1700 ^ _T_1696[3];
  assign _T_1704 = _T_1702 ^ _T_1696[5];
  assign _T_1706 = {_T_1704,_T_1696[15:1]};
  assign _T_1715 = {_T_256[0],_T_244[0],_T_232[0],_T_220[0],_T_208[0],_T_196[0],_T_184[0]};
  assign _T_1723 = {_T_352[0],_T_340[0],_T_328[0],_T_316[0],_T_304[0],_T_292[0],_T_280[0],_T_268[0],_T_1715};
  assign _T_1730 = {_T_448[0],_T_436[0],_T_424[0],_T_412[0],_T_400[0],_T_388[0],_T_376[0],_T_364[0]};
  assign _T_1739 = {_T_544[0],_T_532[0],_T_520[0],_T_508[0],_T_496[0],_T_484[0],_T_472[0],_T_460[0],_T_1730,_T_1723};
  assign _T_1746 = {_T_640[0],_T_628[0],_T_616[0],_T_604[0],_T_592[0],_T_580[0],_T_568[0],_T_556[0]};
  assign _T_1754 = {_T_736[0],_T_724[0],_T_712[0],_T_700[0],_T_688[0],_T_676[0],_T_664[0],_T_652[0],_T_1746};
  assign _T_1761 = {_T_832[0],_T_820[0],_T_808[0],_T_796[0],_T_784[0],_T_772[0],_T_760[0],_T_748[0]};
  assign _T_1770 = {_T_928[0],_T_916[0],_T_904[0],_T_892[0],_T_880[0],_T_868[0],_T_856[0],_T_844[0],_T_1761,_T_1754};
  assign _T_1778 = {_T_1024[0],_T_1012[0],_T_1000[0],_T_988[0],_T_976[0],_T_964[0],_T_952[0],_T_940[0]};
  assign _T_1786 = {_T_1120[0],_T_1108[0],_T_1096[0],_T_1084[0],_T_1072[0],_T_1060[0],_T_1048[0],_T_1036[0],_T_1778};
  assign _T_1793 = {_T_1216[0],_T_1204[0],_T_1192[0],_T_1180[0],_T_1168[0],_T_1156[0],_T_1144[0],_T_1132[0]};
  assign _T_1802 = {_T_1312[0],_T_1300[0],_T_1288[0],_T_1276[0],_T_1264[0],_T_1252[0],_T_1240[0],_T_1228[0],_T_1793,_T_1786};
  assign _T_1809 = {_T_1408[0],_T_1396[0],_T_1384[0],_T_1372[0],_T_1360[0],_T_1348[0],_T_1336[0],_T_1324[0]};
  assign _T_1817 = {_T_1504[0],_T_1492[0],_T_1480[0],_T_1468[0],_T_1456[0],_T_1444[0],_T_1432[0],_T_1420[0],_T_1809};
  assign _T_1824 = {_T_1600[0],_T_1588[0],_T_1576[0],_T_1564[0],_T_1552[0],_T_1540[0],_T_1528[0],_T_1516[0]};
  assign _T_1833 = {_T_1696[0],_T_1684[0],_T_1672[0],_T_1660[0],_T_1648[0],_T_1636[0],_T_1624[0],_T_1612[0],_T_1824,_T_1817};
  assign _T_1835 = {_T_1833,_T_1802,_T_1770,_T_1739};
  assign _T_1836 = _T_42 == 32'h5;
  assign _T_1837 = system_wfi_from_tile_0;
  assign _T_1839 = _T_1838 == 16'h0;
  assign _T_1842 = _T_1838[0] ^ _T_1838[2];
  assign _T_1844 = _T_1842 ^ _T_1838[3];
  assign _T_1846 = _T_1844 ^ _T_1838[5];
  assign _T_1848 = {_T_1846,_T_1838[15:1]};
  assign _T_1851 = _T_1850 == 16'h0;
  assign _T_1854 = _T_1850[0] ^ _T_1850[2];
  assign _T_1856 = _T_1854 ^ _T_1850[3];
  assign _T_1858 = _T_1856 ^ _T_1850[5];
  assign _T_1860 = {_T_1858,_T_1850[15:1]};
  assign _T_1863 = _T_1862 == 16'h0;
  assign _T_1866 = _T_1862[0] ^ _T_1862[2];
  assign _T_1868 = _T_1866 ^ _T_1862[3];
  assign _T_1870 = _T_1868 ^ _T_1862[5];
  assign _T_1872 = {_T_1870,_T_1862[15:1]};
  assign _T_1875 = _T_1874 == 16'h0;
  assign _T_1878 = _T_1874[0] ^ _T_1874[2];
  assign _T_1880 = _T_1878 ^ _T_1874[3];
  assign _T_1882 = _T_1880 ^ _T_1874[5];
  assign _T_1884 = {_T_1882,_T_1874[15:1]};
  assign _T_1887 = _T_1886 == 16'h0;
  assign _T_1890 = _T_1886[0] ^ _T_1886[2];
  assign _T_1892 = _T_1890 ^ _T_1886[3];
  assign _T_1894 = _T_1892 ^ _T_1886[5];
  assign _T_1896 = {_T_1894,_T_1886[15:1]};
  assign _T_1899 = _T_1898 == 16'h0;
  assign _T_1902 = _T_1898[0] ^ _T_1898[2];
  assign _T_1904 = _T_1902 ^ _T_1898[3];
  assign _T_1906 = _T_1904 ^ _T_1898[5];
  assign _T_1908 = {_T_1906,_T_1898[15:1]};
  assign _T_1911 = _T_1910 == 16'h0;
  assign _T_1914 = _T_1910[0] ^ _T_1910[2];
  assign _T_1916 = _T_1914 ^ _T_1910[3];
  assign _T_1918 = _T_1916 ^ _T_1910[5];
  assign _T_1920 = {_T_1918,_T_1910[15:1]};
  assign _T_1923 = _T_1922 == 16'h0;
  assign _T_1926 = _T_1922[0] ^ _T_1922[2];
  assign _T_1928 = _T_1926 ^ _T_1922[3];
  assign _T_1930 = _T_1928 ^ _T_1922[5];
  assign _T_1932 = {_T_1930,_T_1922[15:1]};
  assign _T_1935 = _T_1934 == 16'h0;
  assign _T_1938 = _T_1934[0] ^ _T_1934[2];
  assign _T_1940 = _T_1938 ^ _T_1934[3];
  assign _T_1942 = _T_1940 ^ _T_1934[5];
  assign _T_1944 = {_T_1942,_T_1934[15:1]};
  assign _T_1947 = _T_1946 == 16'h0;
  assign _T_1950 = _T_1946[0] ^ _T_1946[2];
  assign _T_1952 = _T_1950 ^ _T_1946[3];
  assign _T_1954 = _T_1952 ^ _T_1946[5];
  assign _T_1956 = {_T_1954,_T_1946[15:1]};
  assign _T_1959 = _T_1958 == 16'h0;
  assign _T_1962 = _T_1958[0] ^ _T_1958[2];
  assign _T_1964 = _T_1962 ^ _T_1958[3];
  assign _T_1966 = _T_1964 ^ _T_1958[5];
  assign _T_1968 = {_T_1966,_T_1958[15:1]};
  assign _T_1971 = _T_1970 == 16'h0;
  assign _T_1974 = _T_1970[0] ^ _T_1970[2];
  assign _T_1976 = _T_1974 ^ _T_1970[3];
  assign _T_1978 = _T_1976 ^ _T_1970[5];
  assign _T_1980 = {_T_1978,_T_1970[15:1]};
  assign _T_1983 = _T_1982 == 16'h0;
  assign _T_1986 = _T_1982[0] ^ _T_1982[2];
  assign _T_1988 = _T_1986 ^ _T_1982[3];
  assign _T_1990 = _T_1988 ^ _T_1982[5];
  assign _T_1992 = {_T_1990,_T_1982[15:1]};
  assign _T_1995 = _T_1994 == 16'h0;
  assign _T_1998 = _T_1994[0] ^ _T_1994[2];
  assign _T_2000 = _T_1998 ^ _T_1994[3];
  assign _T_2002 = _T_2000 ^ _T_1994[5];
  assign _T_2004 = {_T_2002,_T_1994[15:1]};
  assign _T_2007 = _T_2006 == 16'h0;
  assign _T_2010 = _T_2006[0] ^ _T_2006[2];
  assign _T_2012 = _T_2010 ^ _T_2006[3];
  assign _T_2014 = _T_2012 ^ _T_2006[5];
  assign _T_2016 = {_T_2014,_T_2006[15:1]};
  assign _T_2019 = _T_2018 == 16'h0;
  assign _T_2022 = _T_2018[0] ^ _T_2018[2];
  assign _T_2024 = _T_2022 ^ _T_2018[3];
  assign _T_2026 = _T_2024 ^ _T_2018[5];
  assign _T_2028 = {_T_2026,_T_2018[15:1]};
  assign _T_2031 = _T_2030 == 16'h0;
  assign _T_2034 = _T_2030[0] ^ _T_2030[2];
  assign _T_2036 = _T_2034 ^ _T_2030[3];
  assign _T_2038 = _T_2036 ^ _T_2030[5];
  assign _T_2040 = {_T_2038,_T_2030[15:1]};
  assign _T_2043 = _T_2042 == 16'h0;
  assign _T_2046 = _T_2042[0] ^ _T_2042[2];
  assign _T_2048 = _T_2046 ^ _T_2042[3];
  assign _T_2050 = _T_2048 ^ _T_2042[5];
  assign _T_2052 = {_T_2050,_T_2042[15:1]};
  assign _T_2055 = _T_2054 == 16'h0;
  assign _T_2058 = _T_2054[0] ^ _T_2054[2];
  assign _T_2060 = _T_2058 ^ _T_2054[3];
  assign _T_2062 = _T_2060 ^ _T_2054[5];
  assign _T_2064 = {_T_2062,_T_2054[15:1]};
  assign _T_2067 = _T_2066 == 16'h0;
  assign _T_2070 = _T_2066[0] ^ _T_2066[2];
  assign _T_2072 = _T_2070 ^ _T_2066[3];
  assign _T_2074 = _T_2072 ^ _T_2066[5];
  assign _T_2076 = {_T_2074,_T_2066[15:1]};
  assign _T_2079 = _T_2078 == 16'h0;
  assign _T_2082 = _T_2078[0] ^ _T_2078[2];
  assign _T_2084 = _T_2082 ^ _T_2078[3];
  assign _T_2086 = _T_2084 ^ _T_2078[5];
  assign _T_2088 = {_T_2086,_T_2078[15:1]};
  assign _T_2091 = _T_2090 == 16'h0;
  assign _T_2094 = _T_2090[0] ^ _T_2090[2];
  assign _T_2096 = _T_2094 ^ _T_2090[3];
  assign _T_2098 = _T_2096 ^ _T_2090[5];
  assign _T_2100 = {_T_2098,_T_2090[15:1]};
  assign _T_2103 = _T_2102 == 16'h0;
  assign _T_2106 = _T_2102[0] ^ _T_2102[2];
  assign _T_2108 = _T_2106 ^ _T_2102[3];
  assign _T_2110 = _T_2108 ^ _T_2102[5];
  assign _T_2112 = {_T_2110,_T_2102[15:1]};
  assign _T_2115 = _T_2114 == 16'h0;
  assign _T_2118 = _T_2114[0] ^ _T_2114[2];
  assign _T_2120 = _T_2118 ^ _T_2114[3];
  assign _T_2122 = _T_2120 ^ _T_2114[5];
  assign _T_2124 = {_T_2122,_T_2114[15:1]};
  assign _T_2127 = _T_2126 == 16'h0;
  assign _T_2130 = _T_2126[0] ^ _T_2126[2];
  assign _T_2132 = _T_2130 ^ _T_2126[3];
  assign _T_2134 = _T_2132 ^ _T_2126[5];
  assign _T_2136 = {_T_2134,_T_2126[15:1]};
  assign _T_2139 = _T_2138 == 16'h0;
  assign _T_2142 = _T_2138[0] ^ _T_2138[2];
  assign _T_2144 = _T_2142 ^ _T_2138[3];
  assign _T_2146 = _T_2144 ^ _T_2138[5];
  assign _T_2148 = {_T_2146,_T_2138[15:1]};
  assign _T_2151 = _T_2150 == 16'h0;
  assign _T_2154 = _T_2150[0] ^ _T_2150[2];
  assign _T_2156 = _T_2154 ^ _T_2150[3];
  assign _T_2158 = _T_2156 ^ _T_2150[5];
  assign _T_2160 = {_T_2158,_T_2150[15:1]};
  assign _T_2163 = _T_2162 == 16'h0;
  assign _T_2166 = _T_2162[0] ^ _T_2162[2];
  assign _T_2168 = _T_2166 ^ _T_2162[3];
  assign _T_2170 = _T_2168 ^ _T_2162[5];
  assign _T_2172 = {_T_2170,_T_2162[15:1]};
  assign _T_2175 = _T_2174 == 16'h0;
  assign _T_2178 = _T_2174[0] ^ _T_2174[2];
  assign _T_2180 = _T_2178 ^ _T_2174[3];
  assign _T_2182 = _T_2180 ^ _T_2174[5];
  assign _T_2184 = {_T_2182,_T_2174[15:1]};
  assign _T_2187 = _T_2186 == 16'h0;
  assign _T_2190 = _T_2186[0] ^ _T_2186[2];
  assign _T_2192 = _T_2190 ^ _T_2186[3];
  assign _T_2194 = _T_2192 ^ _T_2186[5];
  assign _T_2196 = {_T_2194,_T_2186[15:1]};
  assign _T_2199 = _T_2198 == 16'h0;
  assign _T_2202 = _T_2198[0] ^ _T_2198[2];
  assign _T_2204 = _T_2202 ^ _T_2198[3];
  assign _T_2206 = _T_2204 ^ _T_2198[5];
  assign _T_2208 = {_T_2206,_T_2198[15:1]};
  assign _T_2211 = _T_2210 == 16'h0;
  assign _T_2214 = _T_2210[0] ^ _T_2210[2];
  assign _T_2216 = _T_2214 ^ _T_2210[3];
  assign _T_2218 = _T_2216 ^ _T_2210[5];
  assign _T_2220 = {_T_2218,_T_2210[15:1]};
  assign _T_2223 = _T_2222 == 16'h0;
  assign _T_2226 = _T_2222[0] ^ _T_2222[2];
  assign _T_2228 = _T_2226 ^ _T_2222[3];
  assign _T_2230 = _T_2228 ^ _T_2222[5];
  assign _T_2232 = {_T_2230,_T_2222[15:1]};
  assign _T_2235 = _T_2234 == 16'h0;
  assign _T_2238 = _T_2234[0] ^ _T_2234[2];
  assign _T_2240 = _T_2238 ^ _T_2234[3];
  assign _T_2242 = _T_2240 ^ _T_2234[5];
  assign _T_2244 = {_T_2242,_T_2234[15:1]};
  assign _T_2247 = _T_2246 == 16'h0;
  assign _T_2250 = _T_2246[0] ^ _T_2246[2];
  assign _T_2252 = _T_2250 ^ _T_2246[3];
  assign _T_2254 = _T_2252 ^ _T_2246[5];
  assign _T_2256 = {_T_2254,_T_2246[15:1]};
  assign _T_2259 = _T_2258 == 16'h0;
  assign _T_2262 = _T_2258[0] ^ _T_2258[2];
  assign _T_2264 = _T_2262 ^ _T_2258[3];
  assign _T_2266 = _T_2264 ^ _T_2258[5];
  assign _T_2268 = {_T_2266,_T_2258[15:1]};
  assign _T_2271 = _T_2270 == 16'h0;
  assign _T_2274 = _T_2270[0] ^ _T_2270[2];
  assign _T_2276 = _T_2274 ^ _T_2270[3];
  assign _T_2278 = _T_2276 ^ _T_2270[5];
  assign _T_2280 = {_T_2278,_T_2270[15:1]};
  assign _T_2283 = _T_2282 == 16'h0;
  assign _T_2286 = _T_2282[0] ^ _T_2282[2];
  assign _T_2288 = _T_2286 ^ _T_2282[3];
  assign _T_2290 = _T_2288 ^ _T_2282[5];
  assign _T_2292 = {_T_2290,_T_2282[15:1]};
  assign _T_2295 = _T_2294 == 16'h0;
  assign _T_2298 = _T_2294[0] ^ _T_2294[2];
  assign _T_2300 = _T_2298 ^ _T_2294[3];
  assign _T_2302 = _T_2300 ^ _T_2294[5];
  assign _T_2304 = {_T_2302,_T_2294[15:1]};
  assign _T_2307 = _T_2306 == 16'h0;
  assign _T_2310 = _T_2306[0] ^ _T_2306[2];
  assign _T_2312 = _T_2310 ^ _T_2306[3];
  assign _T_2314 = _T_2312 ^ _T_2306[5];
  assign _T_2316 = {_T_2314,_T_2306[15:1]};
  assign _T_2319 = _T_2318 == 16'h0;
  assign _T_2322 = _T_2318[0] ^ _T_2318[2];
  assign _T_2324 = _T_2322 ^ _T_2318[3];
  assign _T_2326 = _T_2324 ^ _T_2318[5];
  assign _T_2328 = {_T_2326,_T_2318[15:1]};
  assign _T_2331 = _T_2330 == 16'h0;
  assign _T_2334 = _T_2330[0] ^ _T_2330[2];
  assign _T_2336 = _T_2334 ^ _T_2330[3];
  assign _T_2338 = _T_2336 ^ _T_2330[5];
  assign _T_2340 = {_T_2338,_T_2330[15:1]};
  assign _T_2343 = _T_2342 == 16'h0;
  assign _T_2346 = _T_2342[0] ^ _T_2342[2];
  assign _T_2348 = _T_2346 ^ _T_2342[3];
  assign _T_2350 = _T_2348 ^ _T_2342[5];
  assign _T_2352 = {_T_2350,_T_2342[15:1]};
  assign _T_2355 = _T_2354 == 16'h0;
  assign _T_2358 = _T_2354[0] ^ _T_2354[2];
  assign _T_2360 = _T_2358 ^ _T_2354[3];
  assign _T_2362 = _T_2360 ^ _T_2354[5];
  assign _T_2364 = {_T_2362,_T_2354[15:1]};
  assign _T_2367 = _T_2366 == 16'h0;
  assign _T_2370 = _T_2366[0] ^ _T_2366[2];
  assign _T_2372 = _T_2370 ^ _T_2366[3];
  assign _T_2374 = _T_2372 ^ _T_2366[5];
  assign _T_2376 = {_T_2374,_T_2366[15:1]};
  assign _T_2379 = _T_2378 == 16'h0;
  assign _T_2382 = _T_2378[0] ^ _T_2378[2];
  assign _T_2384 = _T_2382 ^ _T_2378[3];
  assign _T_2386 = _T_2384 ^ _T_2378[5];
  assign _T_2388 = {_T_2386,_T_2378[15:1]};
  assign _T_2391 = _T_2390 == 16'h0;
  assign _T_2394 = _T_2390[0] ^ _T_2390[2];
  assign _T_2396 = _T_2394 ^ _T_2390[3];
  assign _T_2398 = _T_2396 ^ _T_2390[5];
  assign _T_2400 = {_T_2398,_T_2390[15:1]};
  assign _T_2403 = _T_2402 == 16'h0;
  assign _T_2406 = _T_2402[0] ^ _T_2402[2];
  assign _T_2408 = _T_2406 ^ _T_2402[3];
  assign _T_2410 = _T_2408 ^ _T_2402[5];
  assign _T_2412 = {_T_2410,_T_2402[15:1]};
  assign _T_2415 = _T_2414 == 16'h0;
  assign _T_2418 = _T_2414[0] ^ _T_2414[2];
  assign _T_2420 = _T_2418 ^ _T_2414[3];
  assign _T_2422 = _T_2420 ^ _T_2414[5];
  assign _T_2424 = {_T_2422,_T_2414[15:1]};
  assign _T_2427 = _T_2426 == 16'h0;
  assign _T_2430 = _T_2426[0] ^ _T_2426[2];
  assign _T_2432 = _T_2430 ^ _T_2426[3];
  assign _T_2434 = _T_2432 ^ _T_2426[5];
  assign _T_2436 = {_T_2434,_T_2426[15:1]};
  assign _T_2439 = _T_2438 == 16'h0;
  assign _T_2442 = _T_2438[0] ^ _T_2438[2];
  assign _T_2444 = _T_2442 ^ _T_2438[3];
  assign _T_2446 = _T_2444 ^ _T_2438[5];
  assign _T_2448 = {_T_2446,_T_2438[15:1]};
  assign _T_2451 = _T_2450 == 16'h0;
  assign _T_2454 = _T_2450[0] ^ _T_2450[2];
  assign _T_2456 = _T_2454 ^ _T_2450[3];
  assign _T_2458 = _T_2456 ^ _T_2450[5];
  assign _T_2460 = {_T_2458,_T_2450[15:1]};
  assign _T_2463 = _T_2462 == 16'h0;
  assign _T_2466 = _T_2462[0] ^ _T_2462[2];
  assign _T_2468 = _T_2466 ^ _T_2462[3];
  assign _T_2470 = _T_2468 ^ _T_2462[5];
  assign _T_2472 = {_T_2470,_T_2462[15:1]};
  assign _T_2475 = _T_2474 == 16'h0;
  assign _T_2478 = _T_2474[0] ^ _T_2474[2];
  assign _T_2480 = _T_2478 ^ _T_2474[3];
  assign _T_2482 = _T_2480 ^ _T_2474[5];
  assign _T_2484 = {_T_2482,_T_2474[15:1]};
  assign _T_2487 = _T_2486 == 16'h0;
  assign _T_2490 = _T_2486[0] ^ _T_2486[2];
  assign _T_2492 = _T_2490 ^ _T_2486[3];
  assign _T_2494 = _T_2492 ^ _T_2486[5];
  assign _T_2496 = {_T_2494,_T_2486[15:1]};
  assign _T_2499 = _T_2498 == 16'h0;
  assign _T_2502 = _T_2498[0] ^ _T_2498[2];
  assign _T_2504 = _T_2502 ^ _T_2498[3];
  assign _T_2506 = _T_2504 ^ _T_2498[5];
  assign _T_2508 = {_T_2506,_T_2498[15:1]};
  assign _T_2511 = _T_2510 == 16'h0;
  assign _T_2514 = _T_2510[0] ^ _T_2510[2];
  assign _T_2516 = _T_2514 ^ _T_2510[3];
  assign _T_2518 = _T_2516 ^ _T_2510[5];
  assign _T_2520 = {_T_2518,_T_2510[15:1]};
  assign _T_2523 = _T_2522 == 16'h0;
  assign _T_2526 = _T_2522[0] ^ _T_2522[2];
  assign _T_2528 = _T_2526 ^ _T_2522[3];
  assign _T_2530 = _T_2528 ^ _T_2522[5];
  assign _T_2532 = {_T_2530,_T_2522[15:1]};
  assign _T_2535 = _T_2534 == 16'h0;
  assign _T_2538 = _T_2534[0] ^ _T_2534[2];
  assign _T_2540 = _T_2538 ^ _T_2534[3];
  assign _T_2542 = _T_2540 ^ _T_2534[5];
  assign _T_2544 = {_T_2542,_T_2534[15:1]};
  assign _T_2547 = _T_2546 == 16'h0;
  assign _T_2550 = _T_2546[0] ^ _T_2546[2];
  assign _T_2552 = _T_2550 ^ _T_2546[3];
  assign _T_2554 = _T_2552 ^ _T_2546[5];
  assign _T_2556 = {_T_2554,_T_2546[15:1]};
  assign _T_2559 = _T_2558 == 16'h0;
  assign _T_2562 = _T_2558[0] ^ _T_2558[2];
  assign _T_2564 = _T_2562 ^ _T_2558[3];
  assign _T_2566 = _T_2564 ^ _T_2558[5];
  assign _T_2568 = {_T_2566,_T_2558[15:1]};
  assign _T_2571 = _T_2570 == 16'h0;
  assign _T_2574 = _T_2570[0] ^ _T_2570[2];
  assign _T_2576 = _T_2574 ^ _T_2570[3];
  assign _T_2578 = _T_2576 ^ _T_2570[5];
  assign _T_2580 = {_T_2578,_T_2570[15:1]};
  assign _T_2583 = _T_2582 == 16'h0;
  assign _T_2586 = _T_2582[0] ^ _T_2582[2];
  assign _T_2588 = _T_2586 ^ _T_2582[3];
  assign _T_2590 = _T_2588 ^ _T_2582[5];
  assign _T_2592 = {_T_2590,_T_2582[15:1]};
  assign _T_2595 = _T_2594 == 16'h0;
  assign _T_2598 = _T_2594[0] ^ _T_2594[2];
  assign _T_2600 = _T_2598 ^ _T_2594[3];
  assign _T_2602 = _T_2600 ^ _T_2594[5];
  assign _T_2604 = {_T_2602,_T_2594[15:1]};
  assign _T_2607 = _T_2606 == 16'h0;
  assign _T_2610 = _T_2606[0] ^ _T_2606[2];
  assign _T_2612 = _T_2610 ^ _T_2606[3];
  assign _T_2614 = _T_2612 ^ _T_2606[5];
  assign _T_2616 = {_T_2614,_T_2606[15:1]};
  assign _T_2619 = _T_2618 == 16'h0;
  assign _T_2622 = _T_2618[0] ^ _T_2618[2];
  assign _T_2624 = _T_2622 ^ _T_2618[3];
  assign _T_2626 = _T_2624 ^ _T_2618[5];
  assign _T_2628 = {_T_2626,_T_2618[15:1]};
  assign _T_2631 = _T_2630 == 16'h0;
  assign _T_2634 = _T_2630[0] ^ _T_2630[2];
  assign _T_2636 = _T_2634 ^ _T_2630[3];
  assign _T_2638 = _T_2636 ^ _T_2630[5];
  assign _T_2640 = {_T_2638,_T_2630[15:1]};
  assign _T_2643 = _T_2642 == 16'h0;
  assign _T_2646 = _T_2642[0] ^ _T_2642[2];
  assign _T_2648 = _T_2646 ^ _T_2642[3];
  assign _T_2650 = _T_2648 ^ _T_2642[5];
  assign _T_2652 = {_T_2650,_T_2642[15:1]};
  assign _T_2655 = _T_2654 == 16'h0;
  assign _T_2658 = _T_2654[0] ^ _T_2654[2];
  assign _T_2660 = _T_2658 ^ _T_2654[3];
  assign _T_2662 = _T_2660 ^ _T_2654[5];
  assign _T_2664 = {_T_2662,_T_2654[15:1]};
  assign _T_2667 = _T_2666 == 16'h0;
  assign _T_2670 = _T_2666[0] ^ _T_2666[2];
  assign _T_2672 = _T_2670 ^ _T_2666[3];
  assign _T_2674 = _T_2672 ^ _T_2666[5];
  assign _T_2676 = {_T_2674,_T_2666[15:1]};
  assign _T_2679 = _T_2678 == 16'h0;
  assign _T_2682 = _T_2678[0] ^ _T_2678[2];
  assign _T_2684 = _T_2682 ^ _T_2678[3];
  assign _T_2686 = _T_2684 ^ _T_2678[5];
  assign _T_2688 = {_T_2686,_T_2678[15:1]};
  assign _T_2691 = _T_2690 == 16'h0;
  assign _T_2694 = _T_2690[0] ^ _T_2690[2];
  assign _T_2696 = _T_2694 ^ _T_2690[3];
  assign _T_2698 = _T_2696 ^ _T_2690[5];
  assign _T_2700 = {_T_2698,_T_2690[15:1]};
  assign _T_2703 = _T_2702 == 16'h0;
  assign _T_2706 = _T_2702[0] ^ _T_2702[2];
  assign _T_2708 = _T_2706 ^ _T_2702[3];
  assign _T_2710 = _T_2708 ^ _T_2702[5];
  assign _T_2712 = {_T_2710,_T_2702[15:1]};
  assign _T_2715 = _T_2714 == 16'h0;
  assign _T_2718 = _T_2714[0] ^ _T_2714[2];
  assign _T_2720 = _T_2718 ^ _T_2714[3];
  assign _T_2722 = _T_2720 ^ _T_2714[5];
  assign _T_2724 = {_T_2722,_T_2714[15:1]};
  assign _T_2727 = _T_2726 == 16'h0;
  assign _T_2730 = _T_2726[0] ^ _T_2726[2];
  assign _T_2732 = _T_2730 ^ _T_2726[3];
  assign _T_2734 = _T_2732 ^ _T_2726[5];
  assign _T_2736 = {_T_2734,_T_2726[15:1]};
  assign _T_2739 = _T_2738 == 16'h0;
  assign _T_2742 = _T_2738[0] ^ _T_2738[2];
  assign _T_2744 = _T_2742 ^ _T_2738[3];
  assign _T_2746 = _T_2744 ^ _T_2738[5];
  assign _T_2748 = {_T_2746,_T_2738[15:1]};
  assign _T_2751 = _T_2750 == 16'h0;
  assign _T_2754 = _T_2750[0] ^ _T_2750[2];
  assign _T_2756 = _T_2754 ^ _T_2750[3];
  assign _T_2758 = _T_2756 ^ _T_2750[5];
  assign _T_2760 = {_T_2758,_T_2750[15:1]};
  assign _T_2763 = _T_2762 == 16'h0;
  assign _T_2766 = _T_2762[0] ^ _T_2762[2];
  assign _T_2768 = _T_2766 ^ _T_2762[3];
  assign _T_2770 = _T_2768 ^ _T_2762[5];
  assign _T_2772 = {_T_2770,_T_2762[15:1]};
  assign _T_2775 = _T_2774 == 16'h0;
  assign _T_2778 = _T_2774[0] ^ _T_2774[2];
  assign _T_2780 = _T_2778 ^ _T_2774[3];
  assign _T_2782 = _T_2780 ^ _T_2774[5];
  assign _T_2784 = {_T_2782,_T_2774[15:1]};
  assign _T_2787 = _T_2786 == 16'h0;
  assign _T_2790 = _T_2786[0] ^ _T_2786[2];
  assign _T_2792 = _T_2790 ^ _T_2786[3];
  assign _T_2794 = _T_2792 ^ _T_2786[5];
  assign _T_2796 = {_T_2794,_T_2786[15:1]};
  assign _T_2799 = _T_2798 == 16'h0;
  assign _T_2802 = _T_2798[0] ^ _T_2798[2];
  assign _T_2804 = _T_2802 ^ _T_2798[3];
  assign _T_2806 = _T_2804 ^ _T_2798[5];
  assign _T_2808 = {_T_2806,_T_2798[15:1]};
  assign _T_2811 = _T_2810 == 16'h0;
  assign _T_2814 = _T_2810[0] ^ _T_2810[2];
  assign _T_2816 = _T_2814 ^ _T_2810[3];
  assign _T_2818 = _T_2816 ^ _T_2810[5];
  assign _T_2820 = {_T_2818,_T_2810[15:1]};
  assign _T_2823 = _T_2822 == 16'h0;
  assign _T_2826 = _T_2822[0] ^ _T_2822[2];
  assign _T_2828 = _T_2826 ^ _T_2822[3];
  assign _T_2830 = _T_2828 ^ _T_2822[5];
  assign _T_2832 = {_T_2830,_T_2822[15:1]};
  assign _T_2835 = _T_2834 == 16'h0;
  assign _T_2838 = _T_2834[0] ^ _T_2834[2];
  assign _T_2840 = _T_2838 ^ _T_2834[3];
  assign _T_2842 = _T_2840 ^ _T_2834[5];
  assign _T_2844 = {_T_2842,_T_2834[15:1]};
  assign _T_2847 = _T_2846 == 16'h0;
  assign _T_2850 = _T_2846[0] ^ _T_2846[2];
  assign _T_2852 = _T_2850 ^ _T_2846[3];
  assign _T_2854 = _T_2852 ^ _T_2846[5];
  assign _T_2856 = {_T_2854,_T_2846[15:1]};
  assign _T_2859 = _T_2858 == 16'h0;
  assign _T_2862 = _T_2858[0] ^ _T_2858[2];
  assign _T_2864 = _T_2862 ^ _T_2858[3];
  assign _T_2866 = _T_2864 ^ _T_2858[5];
  assign _T_2868 = {_T_2866,_T_2858[15:1]};
  assign _T_2871 = _T_2870 == 16'h0;
  assign _T_2874 = _T_2870[0] ^ _T_2870[2];
  assign _T_2876 = _T_2874 ^ _T_2870[3];
  assign _T_2878 = _T_2876 ^ _T_2870[5];
  assign _T_2880 = {_T_2878,_T_2870[15:1]};
  assign _T_2883 = _T_2882 == 16'h0;
  assign _T_2886 = _T_2882[0] ^ _T_2882[2];
  assign _T_2888 = _T_2886 ^ _T_2882[3];
  assign _T_2890 = _T_2888 ^ _T_2882[5];
  assign _T_2892 = {_T_2890,_T_2882[15:1]};
  assign _T_2895 = _T_2894 == 16'h0;
  assign _T_2898 = _T_2894[0] ^ _T_2894[2];
  assign _T_2900 = _T_2898 ^ _T_2894[3];
  assign _T_2902 = _T_2900 ^ _T_2894[5];
  assign _T_2904 = {_T_2902,_T_2894[15:1]};
  assign _T_2907 = _T_2906 == 16'h0;
  assign _T_2910 = _T_2906[0] ^ _T_2906[2];
  assign _T_2912 = _T_2910 ^ _T_2906[3];
  assign _T_2914 = _T_2912 ^ _T_2906[5];
  assign _T_2916 = {_T_2914,_T_2906[15:1]};
  assign _T_2919 = _T_2918 == 16'h0;
  assign _T_2922 = _T_2918[0] ^ _T_2918[2];
  assign _T_2924 = _T_2922 ^ _T_2918[3];
  assign _T_2926 = _T_2924 ^ _T_2918[5];
  assign _T_2928 = {_T_2926,_T_2918[15:1]};
  assign _T_2931 = _T_2930 == 16'h0;
  assign _T_2934 = _T_2930[0] ^ _T_2930[2];
  assign _T_2936 = _T_2934 ^ _T_2930[3];
  assign _T_2938 = _T_2936 ^ _T_2930[5];
  assign _T_2940 = {_T_2938,_T_2930[15:1]};
  assign _T_2943 = _T_2942 == 16'h0;
  assign _T_2946 = _T_2942[0] ^ _T_2942[2];
  assign _T_2948 = _T_2946 ^ _T_2942[3];
  assign _T_2950 = _T_2948 ^ _T_2942[5];
  assign _T_2952 = {_T_2950,_T_2942[15:1]};
  assign _T_2955 = _T_2954 == 16'h0;
  assign _T_2958 = _T_2954[0] ^ _T_2954[2];
  assign _T_2960 = _T_2958 ^ _T_2954[3];
  assign _T_2962 = _T_2960 ^ _T_2954[5];
  assign _T_2964 = {_T_2962,_T_2954[15:1]};
  assign _T_2967 = _T_2966 == 16'h0;
  assign _T_2970 = _T_2966[0] ^ _T_2966[2];
  assign _T_2972 = _T_2970 ^ _T_2966[3];
  assign _T_2974 = _T_2972 ^ _T_2966[5];
  assign _T_2976 = {_T_2974,_T_2966[15:1]};
  assign _T_2979 = _T_2978 == 16'h0;
  assign _T_2982 = _T_2978[0] ^ _T_2978[2];
  assign _T_2984 = _T_2982 ^ _T_2978[3];
  assign _T_2986 = _T_2984 ^ _T_2978[5];
  assign _T_2988 = {_T_2986,_T_2978[15:1]};
  assign _T_2991 = _T_2990 == 16'h0;
  assign _T_2994 = _T_2990[0] ^ _T_2990[2];
  assign _T_2996 = _T_2994 ^ _T_2990[3];
  assign _T_2998 = _T_2996 ^ _T_2990[5];
  assign _T_3000 = {_T_2998,_T_2990[15:1]};
  assign _T_3003 = _T_3002 == 16'h0;
  assign _T_3006 = _T_3002[0] ^ _T_3002[2];
  assign _T_3008 = _T_3006 ^ _T_3002[3];
  assign _T_3010 = _T_3008 ^ _T_3002[5];
  assign _T_3012 = {_T_3010,_T_3002[15:1]};
  assign _T_3015 = _T_3014 == 16'h0;
  assign _T_3018 = _T_3014[0] ^ _T_3014[2];
  assign _T_3020 = _T_3018 ^ _T_3014[3];
  assign _T_3022 = _T_3020 ^ _T_3014[5];
  assign _T_3024 = {_T_3022,_T_3014[15:1]};
  assign _T_3027 = _T_3026 == 16'h0;
  assign _T_3030 = _T_3026[0] ^ _T_3026[2];
  assign _T_3032 = _T_3030 ^ _T_3026[3];
  assign _T_3034 = _T_3032 ^ _T_3026[5];
  assign _T_3036 = {_T_3034,_T_3026[15:1]};
  assign _T_3039 = _T_3038 == 16'h0;
  assign _T_3042 = _T_3038[0] ^ _T_3038[2];
  assign _T_3044 = _T_3042 ^ _T_3038[3];
  assign _T_3046 = _T_3044 ^ _T_3038[5];
  assign _T_3048 = {_T_3046,_T_3038[15:1]};
  assign _T_3051 = _T_3050 == 16'h0;
  assign _T_3054 = _T_3050[0] ^ _T_3050[2];
  assign _T_3056 = _T_3054 ^ _T_3050[3];
  assign _T_3058 = _T_3056 ^ _T_3050[5];
  assign _T_3060 = {_T_3058,_T_3050[15:1]};
  assign _T_3063 = _T_3062 == 16'h0;
  assign _T_3066 = _T_3062[0] ^ _T_3062[2];
  assign _T_3068 = _T_3066 ^ _T_3062[3];
  assign _T_3070 = _T_3068 ^ _T_3062[5];
  assign _T_3072 = {_T_3070,_T_3062[15:1]};
  assign _T_3075 = _T_3074 == 16'h0;
  assign _T_3078 = _T_3074[0] ^ _T_3074[2];
  assign _T_3080 = _T_3078 ^ _T_3074[3];
  assign _T_3082 = _T_3080 ^ _T_3074[5];
  assign _T_3084 = {_T_3082,_T_3074[15:1]};
  assign _T_3087 = _T_3086 == 16'h0;
  assign _T_3090 = _T_3086[0] ^ _T_3086[2];
  assign _T_3092 = _T_3090 ^ _T_3086[3];
  assign _T_3094 = _T_3092 ^ _T_3086[5];
  assign _T_3096 = {_T_3094,_T_3086[15:1]};
  assign _T_3099 = _T_3098 == 16'h0;
  assign _T_3102 = _T_3098[0] ^ _T_3098[2];
  assign _T_3104 = _T_3102 ^ _T_3098[3];
  assign _T_3106 = _T_3104 ^ _T_3098[5];
  assign _T_3108 = {_T_3106,_T_3098[15:1]};
  assign _T_3111 = _T_3110 == 16'h0;
  assign _T_3114 = _T_3110[0] ^ _T_3110[2];
  assign _T_3116 = _T_3114 ^ _T_3110[3];
  assign _T_3118 = _T_3116 ^ _T_3110[5];
  assign _T_3120 = {_T_3118,_T_3110[15:1]};
  assign _T_3123 = _T_3122 == 16'h0;
  assign _T_3126 = _T_3122[0] ^ _T_3122[2];
  assign _T_3128 = _T_3126 ^ _T_3122[3];
  assign _T_3130 = _T_3128 ^ _T_3122[5];
  assign _T_3132 = {_T_3130,_T_3122[15:1]};
  assign _T_3135 = _T_3134 == 16'h0;
  assign _T_3138 = _T_3134[0] ^ _T_3134[2];
  assign _T_3140 = _T_3138 ^ _T_3134[3];
  assign _T_3142 = _T_3140 ^ _T_3134[5];
  assign _T_3144 = {_T_3142,_T_3134[15:1]};
  assign _T_3147 = _T_3146 == 16'h0;
  assign _T_3150 = _T_3146[0] ^ _T_3146[2];
  assign _T_3152 = _T_3150 ^ _T_3146[3];
  assign _T_3154 = _T_3152 ^ _T_3146[5];
  assign _T_3156 = {_T_3154,_T_3146[15:1]};
  assign _T_3159 = _T_3158 == 16'h0;
  assign _T_3162 = _T_3158[0] ^ _T_3158[2];
  assign _T_3164 = _T_3162 ^ _T_3158[3];
  assign _T_3166 = _T_3164 ^ _T_3158[5];
  assign _T_3168 = {_T_3166,_T_3158[15:1]};
  assign _T_3171 = _T_3170 == 16'h0;
  assign _T_3174 = _T_3170[0] ^ _T_3170[2];
  assign _T_3176 = _T_3174 ^ _T_3170[3];
  assign _T_3178 = _T_3176 ^ _T_3170[5];
  assign _T_3180 = {_T_3178,_T_3170[15:1]};
  assign _T_3183 = _T_3182 == 16'h0;
  assign _T_3186 = _T_3182[0] ^ _T_3182[2];
  assign _T_3188 = _T_3186 ^ _T_3182[3];
  assign _T_3190 = _T_3188 ^ _T_3182[5];
  assign _T_3192 = {_T_3190,_T_3182[15:1]};
  assign _T_3195 = _T_3194 == 16'h0;
  assign _T_3198 = _T_3194[0] ^ _T_3194[2];
  assign _T_3200 = _T_3198 ^ _T_3194[3];
  assign _T_3202 = _T_3200 ^ _T_3194[5];
  assign _T_3204 = {_T_3202,_T_3194[15:1]};
  assign _T_3207 = _T_3206 == 16'h0;
  assign _T_3210 = _T_3206[0] ^ _T_3206[2];
  assign _T_3212 = _T_3210 ^ _T_3206[3];
  assign _T_3214 = _T_3212 ^ _T_3206[5];
  assign _T_3216 = {_T_3214,_T_3206[15:1]};
  assign _T_3219 = _T_3218 == 16'h0;
  assign _T_3222 = _T_3218[0] ^ _T_3218[2];
  assign _T_3224 = _T_3222 ^ _T_3218[3];
  assign _T_3226 = _T_3224 ^ _T_3218[5];
  assign _T_3228 = {_T_3226,_T_3218[15:1]};
  assign _T_3231 = _T_3230 == 16'h0;
  assign _T_3234 = _T_3230[0] ^ _T_3230[2];
  assign _T_3236 = _T_3234 ^ _T_3230[3];
  assign _T_3238 = _T_3236 ^ _T_3230[5];
  assign _T_3240 = {_T_3238,_T_3230[15:1]};
  assign _T_3243 = _T_3242 == 16'h0;
  assign _T_3246 = _T_3242[0] ^ _T_3242[2];
  assign _T_3248 = _T_3246 ^ _T_3242[3];
  assign _T_3250 = _T_3248 ^ _T_3242[5];
  assign _T_3252 = {_T_3250,_T_3242[15:1]};
  assign _T_3255 = _T_3254 == 16'h0;
  assign _T_3258 = _T_3254[0] ^ _T_3254[2];
  assign _T_3260 = _T_3258 ^ _T_3254[3];
  assign _T_3262 = _T_3260 ^ _T_3254[5];
  assign _T_3264 = {_T_3262,_T_3254[15:1]};
  assign _T_3267 = _T_3266 == 16'h0;
  assign _T_3270 = _T_3266[0] ^ _T_3266[2];
  assign _T_3272 = _T_3270 ^ _T_3266[3];
  assign _T_3274 = _T_3272 ^ _T_3266[5];
  assign _T_3276 = {_T_3274,_T_3266[15:1]};
  assign _T_3279 = _T_3278 == 16'h0;
  assign _T_3282 = _T_3278[0] ^ _T_3278[2];
  assign _T_3284 = _T_3282 ^ _T_3278[3];
  assign _T_3286 = _T_3284 ^ _T_3278[5];
  assign _T_3288 = {_T_3286,_T_3278[15:1]};
  assign _T_3291 = _T_3290 == 16'h0;
  assign _T_3294 = _T_3290[0] ^ _T_3290[2];
  assign _T_3296 = _T_3294 ^ _T_3290[3];
  assign _T_3298 = _T_3296 ^ _T_3290[5];
  assign _T_3300 = {_T_3298,_T_3290[15:1]};
  assign _T_3303 = _T_3302 == 16'h0;
  assign _T_3306 = _T_3302[0] ^ _T_3302[2];
  assign _T_3308 = _T_3306 ^ _T_3302[3];
  assign _T_3310 = _T_3308 ^ _T_3302[5];
  assign _T_3312 = {_T_3310,_T_3302[15:1]};
  assign _T_3315 = _T_3314 == 16'h0;
  assign _T_3318 = _T_3314[0] ^ _T_3314[2];
  assign _T_3320 = _T_3318 ^ _T_3314[3];
  assign _T_3322 = _T_3320 ^ _T_3314[5];
  assign _T_3324 = {_T_3322,_T_3314[15:1]};
  assign _T_3327 = _T_3326 == 16'h0;
  assign _T_3330 = _T_3326[0] ^ _T_3326[2];
  assign _T_3332 = _T_3330 ^ _T_3326[3];
  assign _T_3334 = _T_3332 ^ _T_3326[5];
  assign _T_3336 = {_T_3334,_T_3326[15:1]};
  assign _T_3339 = _T_3338 == 16'h0;
  assign _T_3342 = _T_3338[0] ^ _T_3338[2];
  assign _T_3344 = _T_3342 ^ _T_3338[3];
  assign _T_3346 = _T_3344 ^ _T_3338[5];
  assign _T_3348 = {_T_3346,_T_3338[15:1]};
  assign _T_3351 = _T_3350 == 16'h0;
  assign _T_3354 = _T_3350[0] ^ _T_3350[2];
  assign _T_3356 = _T_3354 ^ _T_3350[3];
  assign _T_3358 = _T_3356 ^ _T_3350[5];
  assign _T_3360 = {_T_3358,_T_3350[15:1]};
  assign _T_3369 = {_T_1910[0],_T_1898[0],_T_1886[0],_T_1874[0],_T_1862[0],_T_1850[0],_T_1838[0]};
  assign _T_3377 = {_T_2006[0],_T_1994[0],_T_1982[0],_T_1970[0],_T_1958[0],_T_1946[0],_T_1934[0],_T_1922[0],_T_3369};
  assign _T_3384 = {_T_2102[0],_T_2090[0],_T_2078[0],_T_2066[0],_T_2054[0],_T_2042[0],_T_2030[0],_T_2018[0]};
  assign _T_3393 = {_T_2198[0],_T_2186[0],_T_2174[0],_T_2162[0],_T_2150[0],_T_2138[0],_T_2126[0],_T_2114[0],_T_3384,_T_3377};
  assign _T_3400 = {_T_2294[0],_T_2282[0],_T_2270[0],_T_2258[0],_T_2246[0],_T_2234[0],_T_2222[0],_T_2210[0]};
  assign _T_3408 = {_T_2390[0],_T_2378[0],_T_2366[0],_T_2354[0],_T_2342[0],_T_2330[0],_T_2318[0],_T_2306[0],_T_3400};
  assign _T_3415 = {_T_2486[0],_T_2474[0],_T_2462[0],_T_2450[0],_T_2438[0],_T_2426[0],_T_2414[0],_T_2402[0]};
  assign _T_3424 = {_T_2582[0],_T_2570[0],_T_2558[0],_T_2546[0],_T_2534[0],_T_2522[0],_T_2510[0],_T_2498[0],_T_3415,_T_3408};
  assign _T_3432 = {_T_2678[0],_T_2666[0],_T_2654[0],_T_2642[0],_T_2630[0],_T_2618[0],_T_2606[0],_T_2594[0]};
  assign _T_3440 = {_T_2774[0],_T_2762[0],_T_2750[0],_T_2738[0],_T_2726[0],_T_2714[0],_T_2702[0],_T_2690[0],_T_3432};
  assign _T_3447 = {_T_2870[0],_T_2858[0],_T_2846[0],_T_2834[0],_T_2822[0],_T_2810[0],_T_2798[0],_T_2786[0]};
  assign _T_3456 = {_T_2966[0],_T_2954[0],_T_2942[0],_T_2930[0],_T_2918[0],_T_2906[0],_T_2894[0],_T_2882[0],_T_3447,_T_3440};
  assign _T_3463 = {_T_3062[0],_T_3050[0],_T_3038[0],_T_3026[0],_T_3014[0],_T_3002[0],_T_2990[0],_T_2978[0]};
  assign _T_3471 = {_T_3158[0],_T_3146[0],_T_3134[0],_T_3122[0],_T_3110[0],_T_3098[0],_T_3086[0],_T_3074[0],_T_3463};
  assign _T_3478 = {_T_3254[0],_T_3242[0],_T_3230[0],_T_3218[0],_T_3206[0],_T_3194[0],_T_3182[0],_T_3170[0]};
  assign _T_3487 = {_T_3350[0],_T_3338[0],_T_3326[0],_T_3314[0],_T_3302[0],_T_3290[0],_T_3278[0],_T_3266[0],_T_3478,_T_3471};
  assign _T_3489 = {_T_3487,_T_3456,_T_3424,_T_3393};
  assign _GEN_514 = _T_1837 ? NullInterruptDriver_interrupts : _T_3489;
  assign _GEN_515 = _T_1836 ? _GEN_514 : 127'h0;
  assign _GEN_516 = _T_183 ? _T_1835 : _GEN_515;
  assign _GEN_517 = _T_177 ? _T_182 : {{1'd0}, _GEN_516};
  assign _GEN_518 = _T_49 ? 128'h2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa : _GEN_517;
  assign _GEN_519 = _T_47 ? 128'h7fffffffffffffffffffffffffffffff : _GEN_518;
  assign _GEN_520 = _T_46 ? {{1'd0}, NullInterruptDriver_interrupts} : _GEN_519;
  assign _T_18 = DataTap_2__0;
  assign _T_19 = DataTap_2__1;
  assign _T_25 = DataTap_2__7;
  assign io_success = 1'h1;
  assign system_clock = dpiClockGate_clock_out;
  assign system_reset = reset | system_debug_ndreset;
  assign system_psd_test_clock_enable = 1'h0;
  assign system_meip_0 = 1'h0;
  assign system_resetctrl_hartIsInReset_0 = debug_compatibility_debug_resetctrl_hartIsInReset_0;
  assign system_debug_clock = debug_compatibility_debug_clock;
  assign system_debug_reset = debug_compatibility_debug_reset;
  assign system_debug_systemjtag_jtag_TCK = 1'h1;
  assign system_debug_systemjtag_jtag_TMS = 1'h1;
  assign system_debug_systemjtag_jtag_TDI = 1'h1;
  assign system_debug_systemjtag_reset = reset;
  assign system_debug_systemjtag_mfr_id = 11'h0;
  assign system_debug_systemjtag_part_number = 16'h0;
  assign system_debug_systemjtag_version = 4'h0;
  assign system_debug_dmactiveAck = debug_compatibility_debug_dmactiveAck;
  assign system_reset_vector_0 = 32'h20000000;
  assign system_rtc_toggle = _T_3;
  assign system_local_interrupts_0 = _GEN_520[126:0];
  assign system_sys_port_ahb_0_hready = testRAM_1_io_ahb_0_hready;
  assign system_sys_port_ahb_0_hresp = testRAM_1_io_ahb_0_hresp;
  assign system_sys_port_ahb_0_hrdata = testRAM_1_io_ahb_0_hrdata;
  assign system_periph_port_ahb_0_hready = testRAM_io_ahb_0_hready;
  assign system_periph_port_ahb_0_hresp = testRAM_io_ahb_0_hresp;
  assign system_periph_port_ahb_0_hrdata = testRAM_io_ahb_0_hrdata;
  assign system_front_port_ahb_0_hmastlock = 1'h0;
  assign system_front_port_ahb_0_hsel = 1'h0;
  assign system_front_port_ahb_0_hready = 1'h0;
  assign system_front_port_ahb_0_htrans = 2'h0;
  assign system_front_port_ahb_0_hsize = 3'h0;
  assign system_front_port_ahb_0_hburst = 3'h0;
  assign system_front_port_ahb_0_hwrite = 1'h0;
  assign system_front_port_ahb_0_hprot = 4'h3;
  assign system_front_port_ahb_0_haddr = 32'h0;
  assign system_front_port_ahb_0_hwdata = 32'h0;
  assign func_clock_clock = clock;
  assign dpiClockGate_clock_in = func_clock_io_clock_out;
  assign c_core_reset_driver_clock = clock;
  assign debug_compatibility_clock = system_clock;
  assign debug_compatibility_reset = system_reset;
  assign debug_compatibility_debug_outer_reset = system_debug_systemjtag_reset;
  assign debug_compatibility_debug_dmactive = system_debug_dmactive;
  assign testRAM_clock = dpiClockGate_clock_out;
  assign testRAM_reset = _T_13 | reset;
  assign testRAM_io_ahb_0_htrans = system_periph_port_ahb_0_htrans;
  assign testRAM_io_ahb_0_hsize = system_periph_port_ahb_0_hsize;
  assign testRAM_io_ahb_0_hwrite = system_periph_port_ahb_0_hwrite;
  assign testRAM_io_ahb_0_haddr = system_periph_port_ahb_0_haddr;
  assign testRAM_io_ahb_0_hwdata = system_periph_port_ahb_0_hwdata;
  assign testRAM_1_clock = dpiClockGate_clock_out;
  assign testRAM_1_reset = _T_13 | reset;
  assign testRAM_1_io_ahb_0_htrans = system_sys_port_ahb_0_htrans;
  assign testRAM_1_io_ahb_0_hsize = system_sys_port_ahb_0_hsize;
  assign testRAM_1_io_ahb_0_hwrite = system_sys_port_ahb_0_hwrite;
  assign testRAM_1_io_ahb_0_haddr = system_sys_port_ahb_0_haddr;
  assign testRAM_1_io_ahb_0_hwdata = system_sys_port_ahb_0_hwdata;
  assign WfiChecker_reset = reset;
  assign WfiChecker_clock = clock;
  assign WfiChecker_wfi = system_wfi_from_tile_0;
  assign WfiChecker_excpt = DataTap_2__5;
  assign WfiChecker_bus_err_int = 1'h0;
  assign WfiChecker_debug_int = DataTap_2__6;
  assign WfiChecker_clint_int = _T_25[0];
  assign WfiChecker_allow_wfi = DataTap_2__8;
  assign WfiChecker_debug = DataTap_2__9;
  assign WfiChecker_singleStep = DataTap_2__10;
  assign WfiChecker_reg_mie = {{16'd0}, _T_18};
  assign WfiChecker_reg_mip = _T_19[31:0];
  assign WfiChecker_inst_vld_0 = DataTap_9__0_valid;
  assign WfiChecker_pc_0 = DataTap_9__0_pc;
  assign WfiChecker_inst_0 = DataTap_9__0_inst;
  assign core_monitor_m_0_clock = DataTap_9__0_clock;
  assign core_monitor_m_0_reset = DataTap_9__0_reset;
  assign core_monitor_m_0_excpt = DataTap_9__0_excpt;
  assign core_monitor_m_0_priv_mode = DataTap_9__0_priv_mode;
  assign core_monitor_m_0_hartid = DataTap_9__0_hartid;
  assign core_monitor_m_0_timer = DataTap_9__0_timer;
  assign core_monitor_m_0_valid = DataTap_9__0_valid;
  assign core_monitor_m_0_pc = DataTap_9__0_pc;
  assign core_monitor_m_0_wrdst = DataTap_9__0_wrdst;
  assign core_monitor_m_0_wrdata = DataTap_9__0_wrdata;
  assign core_monitor_m_0_wrenx = DataTap_9__0_wrenx;
  assign core_monitor_m_0_wrenf = DataTap_9__0_wrenf;
  assign core_monitor_m_0_rd0src = DataTap_9__0_rd0src;
  assign core_monitor_m_0_rd0val = DataTap_9__0_rd0val;
  assign core_monitor_m_0_rd1src = DataTap_9__0_rd1src;
  assign core_monitor_m_0_rd1val = DataTap_9__0_rd1val;
  assign core_monitor_m_0_inst = DataTap_9__0_inst;
  assign dpitbh_clock = 1'h0;
  assign dpitbh_reset = 1'h0;
  assign GlobalIntDriver_clock = 1'h0;
  assign GlobalIntDriver_reset = 1'h0;
  assign NullInterruptDriver_clock = 1'h0;
  assign NullInterruptDriver_reset = 1'h0;
  assign _GEN_521 = ~_T_34;
  assign _GEN_522 = ~_T_35;
  assign _GEN_523 = _GEN_521 & _GEN_522;
  assign _GEN_524 = ~_T_36;
  assign _GEN_525 = _GEN_523 & _GEN_524;
  assign _GEN_526 = ~_T_37;
  assign _GEN_527 = _GEN_525 & _GEN_526;
  assign _GEN_528 = ~_T_38;
  assign _GEN_529 = _GEN_527 & _GEN_528;
  assign _GEN_539 = ~_T_46;
  assign _GEN_540 = ~_T_47;
  assign _GEN_541 = _GEN_539 & _GEN_540;
  assign _GEN_542 = ~_T_49;
  assign _GEN_543 = _GEN_541 & _GEN_542;
  assign _GEN_544 = ~_T_177;
  assign _GEN_545 = _GEN_543 & _GEN_544;
  assign _GEN_546 = ~_T_183;
  assign _GEN_547 = _GEN_545 & _GEN_546;
  assign _GEN_548 = ~_T_1836;
  assign _GEN_549 = _GEN_547 & _GEN_548;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_3 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_2 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_184 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_196 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_208 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_220 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_232 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_244 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_256 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_268 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_280 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_292 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_304 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_316 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_328 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_340 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_352 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_364 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_376 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_388 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_400 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_412 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_424 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_436 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_448 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_460 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_472 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_484 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_496 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_508 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_520 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_532 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_544 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_556 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_568 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_580 = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_592 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_604 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_616 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_628 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_640 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_652 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_664 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_676 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_688 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_700 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_712 = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_724 = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_736 = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_748 = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_760 = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_772 = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_784 = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_796 = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_808 = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_820 = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_832 = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_844 = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_856 = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_868 = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_880 = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_892 = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_904 = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_916 = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_928 = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_940 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_952 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_964 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_976 = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_988 = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_1000 = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_1012 = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_1024 = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_1036 = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_1048 = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_1060 = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_1072 = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_1084 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_1096 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_1108 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_1120 = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_1132 = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_1144 = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_1156 = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_1168 = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_1180 = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_1192 = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_1204 = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_1216 = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_1228 = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_1240 = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_1252 = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_1264 = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_1276 = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_1288 = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_1300 = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_1312 = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_1324 = _RAND_99[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_1336 = _RAND_100[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_1348 = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_1360 = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_1372 = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_1384 = _RAND_104[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_1396 = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_1408 = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_1420 = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_1432 = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_1444 = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_1456 = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_1468 = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_1480 = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_1492 = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_1504 = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_1516 = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_1528 = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_1540 = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_1552 = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_1564 = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_1576 = _RAND_120[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_1588 = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_1600 = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_1612 = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_1624 = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_1636 = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_1648 = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_1660 = _RAND_127[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_1672 = _RAND_128[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_1684 = _RAND_129[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_1696 = _RAND_130[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_1838 = _RAND_131[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_1850 = _RAND_132[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_1862 = _RAND_133[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_1874 = _RAND_134[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_1886 = _RAND_135[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_1898 = _RAND_136[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_1910 = _RAND_137[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_1922 = _RAND_138[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_1934 = _RAND_139[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_1946 = _RAND_140[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_1958 = _RAND_141[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_1970 = _RAND_142[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_1982 = _RAND_143[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_1994 = _RAND_144[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_2006 = _RAND_145[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_2018 = _RAND_146[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_2030 = _RAND_147[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_2042 = _RAND_148[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_2054 = _RAND_149[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_2066 = _RAND_150[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_2078 = _RAND_151[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_2090 = _RAND_152[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_2102 = _RAND_153[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_2114 = _RAND_154[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_2126 = _RAND_155[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_2138 = _RAND_156[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_2150 = _RAND_157[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_2162 = _RAND_158[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_2174 = _RAND_159[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_2186 = _RAND_160[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_2198 = _RAND_161[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_2210 = _RAND_162[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_2222 = _RAND_163[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_2234 = _RAND_164[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_2246 = _RAND_165[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_2258 = _RAND_166[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_2270 = _RAND_167[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_2282 = _RAND_168[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_2294 = _RAND_169[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_2306 = _RAND_170[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_2318 = _RAND_171[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_2330 = _RAND_172[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_2342 = _RAND_173[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_2354 = _RAND_174[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_2366 = _RAND_175[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_2378 = _RAND_176[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_2390 = _RAND_177[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_2402 = _RAND_178[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_2414 = _RAND_179[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_2426 = _RAND_180[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_2438 = _RAND_181[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_2450 = _RAND_182[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_2462 = _RAND_183[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_2474 = _RAND_184[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_2486 = _RAND_185[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_2498 = _RAND_186[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_2510 = _RAND_187[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_2522 = _RAND_188[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_2534 = _RAND_189[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_2546 = _RAND_190[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_2558 = _RAND_191[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_2570 = _RAND_192[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_2582 = _RAND_193[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_2594 = _RAND_194[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_2606 = _RAND_195[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_2618 = _RAND_196[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_2630 = _RAND_197[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_2642 = _RAND_198[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_2654 = _RAND_199[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_2666 = _RAND_200[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_2678 = _RAND_201[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_2690 = _RAND_202[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_2702 = _RAND_203[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_2714 = _RAND_204[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_2726 = _RAND_205[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_2738 = _RAND_206[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_2750 = _RAND_207[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_2762 = _RAND_208[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_2774 = _RAND_209[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_2786 = _RAND_210[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_2798 = _RAND_211[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_2810 = _RAND_212[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_2822 = _RAND_213[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_2834 = _RAND_214[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_2846 = _RAND_215[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_2858 = _RAND_216[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_2870 = _RAND_217[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_2882 = _RAND_218[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_2894 = _RAND_219[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_2906 = _RAND_220[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_2918 = _RAND_221[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_2930 = _RAND_222[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_2942 = _RAND_223[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_2954 = _RAND_224[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_2966 = _RAND_225[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_2978 = _RAND_226[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_2990 = _RAND_227[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_3002 = _RAND_228[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_3014 = _RAND_229[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_3026 = _RAND_230[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_3038 = _RAND_231[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_3050 = _RAND_232[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_3062 = _RAND_233[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_3074 = _RAND_234[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_3086 = _RAND_235[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_3098 = _RAND_236[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_3110 = _RAND_237[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_3122 = _RAND_238[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_3134 = _RAND_239[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_3146 = _RAND_240[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_3158 = _RAND_241[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_3170 = _RAND_242[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_3182 = _RAND_243[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_3194 = _RAND_244[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_3206 = _RAND_245[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_3218 = _RAND_246[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_3230 = _RAND_247[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_3242 = _RAND_248[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_3254 = _RAND_249[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_3266 = _RAND_250[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_3278 = _RAND_251[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_3290 = _RAND_252[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_3302 = _RAND_253[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_3314 = _RAND_254[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_3326 = _RAND_255[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_3338 = _RAND_256[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_3350 = _RAND_257[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge dpiClockGate_clock_out) begin
    if (reset) begin
      _T_2 <= 5'h0;
    end else begin
      _T_2 <= _T_5;
    end
    if (reset) begin
      _T_3 <= 1'h0;
    end else if (_T_6) begin
      _T_3 <= _T_7;
    end
  end
  always @(posedge clock) begin
    if (reset) begin
      value_1 <= 7'h0;
    end else if (_T_43) begin
      value_1 <= 7'h0;
    end else begin
      value_1 <= _T_45;
    end
    if (reset) begin
      value_2 <= 7'h0;
    end else if (_T_43) begin
      if (_T_179) begin
        value_2 <= 7'h0;
      end else begin
        value_2 <= _T_181;
      end
    end
    if (_T_43) begin
      if (_T_185) begin
        _T_184 <= 16'h1;
      end else begin
        _T_184 <= _T_194;
      end
    end
    if (_T_43) begin
      if (_T_197) begin
        _T_196 <= 16'h1;
      end else begin
        _T_196 <= _T_206;
      end
    end
    if (_T_43) begin
      if (_T_209) begin
        _T_208 <= 16'h1;
      end else begin
        _T_208 <= _T_218;
      end
    end
    if (_T_43) begin
      if (_T_221) begin
        _T_220 <= 16'h1;
      end else begin
        _T_220 <= _T_230;
      end
    end
    if (_T_43) begin
      if (_T_233) begin
        _T_232 <= 16'h1;
      end else begin
        _T_232 <= _T_242;
      end
    end
    if (_T_43) begin
      if (_T_245) begin
        _T_244 <= 16'h1;
      end else begin
        _T_244 <= _T_254;
      end
    end
    if (_T_43) begin
      if (_T_257) begin
        _T_256 <= 16'h1;
      end else begin
        _T_256 <= _T_266;
      end
    end
    if (_T_43) begin
      if (_T_269) begin
        _T_268 <= 16'h1;
      end else begin
        _T_268 <= _T_278;
      end
    end
    if (_T_43) begin
      if (_T_281) begin
        _T_280 <= 16'h1;
      end else begin
        _T_280 <= _T_290;
      end
    end
    if (_T_43) begin
      if (_T_293) begin
        _T_292 <= 16'h1;
      end else begin
        _T_292 <= _T_302;
      end
    end
    if (_T_43) begin
      if (_T_305) begin
        _T_304 <= 16'h1;
      end else begin
        _T_304 <= _T_314;
      end
    end
    if (_T_43) begin
      if (_T_317) begin
        _T_316 <= 16'h1;
      end else begin
        _T_316 <= _T_326;
      end
    end
    if (_T_43) begin
      if (_T_329) begin
        _T_328 <= 16'h1;
      end else begin
        _T_328 <= _T_338;
      end
    end
    if (_T_43) begin
      if (_T_341) begin
        _T_340 <= 16'h1;
      end else begin
        _T_340 <= _T_350;
      end
    end
    if (_T_43) begin
      if (_T_353) begin
        _T_352 <= 16'h1;
      end else begin
        _T_352 <= _T_362;
      end
    end
    if (_T_43) begin
      if (_T_365) begin
        _T_364 <= 16'h1;
      end else begin
        _T_364 <= _T_374;
      end
    end
    if (_T_43) begin
      if (_T_377) begin
        _T_376 <= 16'h1;
      end else begin
        _T_376 <= _T_386;
      end
    end
    if (_T_43) begin
      if (_T_389) begin
        _T_388 <= 16'h1;
      end else begin
        _T_388 <= _T_398;
      end
    end
    if (_T_43) begin
      if (_T_401) begin
        _T_400 <= 16'h1;
      end else begin
        _T_400 <= _T_410;
      end
    end
    if (_T_43) begin
      if (_T_413) begin
        _T_412 <= 16'h1;
      end else begin
        _T_412 <= _T_422;
      end
    end
    if (_T_43) begin
      if (_T_425) begin
        _T_424 <= 16'h1;
      end else begin
        _T_424 <= _T_434;
      end
    end
    if (_T_43) begin
      if (_T_437) begin
        _T_436 <= 16'h1;
      end else begin
        _T_436 <= _T_446;
      end
    end
    if (_T_43) begin
      if (_T_449) begin
        _T_448 <= 16'h1;
      end else begin
        _T_448 <= _T_458;
      end
    end
    if (_T_43) begin
      if (_T_461) begin
        _T_460 <= 16'h1;
      end else begin
        _T_460 <= _T_470;
      end
    end
    if (_T_43) begin
      if (_T_473) begin
        _T_472 <= 16'h1;
      end else begin
        _T_472 <= _T_482;
      end
    end
    if (_T_43) begin
      if (_T_485) begin
        _T_484 <= 16'h1;
      end else begin
        _T_484 <= _T_494;
      end
    end
    if (_T_43) begin
      if (_T_497) begin
        _T_496 <= 16'h1;
      end else begin
        _T_496 <= _T_506;
      end
    end
    if (_T_43) begin
      if (_T_509) begin
        _T_508 <= 16'h1;
      end else begin
        _T_508 <= _T_518;
      end
    end
    if (_T_43) begin
      if (_T_521) begin
        _T_520 <= 16'h1;
      end else begin
        _T_520 <= _T_530;
      end
    end
    if (_T_43) begin
      if (_T_533) begin
        _T_532 <= 16'h1;
      end else begin
        _T_532 <= _T_542;
      end
    end
    if (_T_43) begin
      if (_T_545) begin
        _T_544 <= 16'h1;
      end else begin
        _T_544 <= _T_554;
      end
    end
    if (_T_43) begin
      if (_T_557) begin
        _T_556 <= 16'h1;
      end else begin
        _T_556 <= _T_566;
      end
    end
    if (_T_43) begin
      if (_T_569) begin
        _T_568 <= 16'h1;
      end else begin
        _T_568 <= _T_578;
      end
    end
    if (_T_43) begin
      if (_T_581) begin
        _T_580 <= 16'h1;
      end else begin
        _T_580 <= _T_590;
      end
    end
    if (_T_43) begin
      if (_T_593) begin
        _T_592 <= 16'h1;
      end else begin
        _T_592 <= _T_602;
      end
    end
    if (_T_43) begin
      if (_T_605) begin
        _T_604 <= 16'h1;
      end else begin
        _T_604 <= _T_614;
      end
    end
    if (_T_43) begin
      if (_T_617) begin
        _T_616 <= 16'h1;
      end else begin
        _T_616 <= _T_626;
      end
    end
    if (_T_43) begin
      if (_T_629) begin
        _T_628 <= 16'h1;
      end else begin
        _T_628 <= _T_638;
      end
    end
    if (_T_43) begin
      if (_T_641) begin
        _T_640 <= 16'h1;
      end else begin
        _T_640 <= _T_650;
      end
    end
    if (_T_43) begin
      if (_T_653) begin
        _T_652 <= 16'h1;
      end else begin
        _T_652 <= _T_662;
      end
    end
    if (_T_43) begin
      if (_T_665) begin
        _T_664 <= 16'h1;
      end else begin
        _T_664 <= _T_674;
      end
    end
    if (_T_43) begin
      if (_T_677) begin
        _T_676 <= 16'h1;
      end else begin
        _T_676 <= _T_686;
      end
    end
    if (_T_43) begin
      if (_T_689) begin
        _T_688 <= 16'h1;
      end else begin
        _T_688 <= _T_698;
      end
    end
    if (_T_43) begin
      if (_T_701) begin
        _T_700 <= 16'h1;
      end else begin
        _T_700 <= _T_710;
      end
    end
    if (_T_43) begin
      if (_T_713) begin
        _T_712 <= 16'h1;
      end else begin
        _T_712 <= _T_722;
      end
    end
    if (_T_43) begin
      if (_T_725) begin
        _T_724 <= 16'h1;
      end else begin
        _T_724 <= _T_734;
      end
    end
    if (_T_43) begin
      if (_T_737) begin
        _T_736 <= 16'h1;
      end else begin
        _T_736 <= _T_746;
      end
    end
    if (_T_43) begin
      if (_T_749) begin
        _T_748 <= 16'h1;
      end else begin
        _T_748 <= _T_758;
      end
    end
    if (_T_43) begin
      if (_T_761) begin
        _T_760 <= 16'h1;
      end else begin
        _T_760 <= _T_770;
      end
    end
    if (_T_43) begin
      if (_T_773) begin
        _T_772 <= 16'h1;
      end else begin
        _T_772 <= _T_782;
      end
    end
    if (_T_43) begin
      if (_T_785) begin
        _T_784 <= 16'h1;
      end else begin
        _T_784 <= _T_794;
      end
    end
    if (_T_43) begin
      if (_T_797) begin
        _T_796 <= 16'h1;
      end else begin
        _T_796 <= _T_806;
      end
    end
    if (_T_43) begin
      if (_T_809) begin
        _T_808 <= 16'h1;
      end else begin
        _T_808 <= _T_818;
      end
    end
    if (_T_43) begin
      if (_T_821) begin
        _T_820 <= 16'h1;
      end else begin
        _T_820 <= _T_830;
      end
    end
    if (_T_43) begin
      if (_T_833) begin
        _T_832 <= 16'h1;
      end else begin
        _T_832 <= _T_842;
      end
    end
    if (_T_43) begin
      if (_T_845) begin
        _T_844 <= 16'h1;
      end else begin
        _T_844 <= _T_854;
      end
    end
    if (_T_43) begin
      if (_T_857) begin
        _T_856 <= 16'h1;
      end else begin
        _T_856 <= _T_866;
      end
    end
    if (_T_43) begin
      if (_T_869) begin
        _T_868 <= 16'h1;
      end else begin
        _T_868 <= _T_878;
      end
    end
    if (_T_43) begin
      if (_T_881) begin
        _T_880 <= 16'h1;
      end else begin
        _T_880 <= _T_890;
      end
    end
    if (_T_43) begin
      if (_T_893) begin
        _T_892 <= 16'h1;
      end else begin
        _T_892 <= _T_902;
      end
    end
    if (_T_43) begin
      if (_T_905) begin
        _T_904 <= 16'h1;
      end else begin
        _T_904 <= _T_914;
      end
    end
    if (_T_43) begin
      if (_T_917) begin
        _T_916 <= 16'h1;
      end else begin
        _T_916 <= _T_926;
      end
    end
    if (_T_43) begin
      if (_T_929) begin
        _T_928 <= 16'h1;
      end else begin
        _T_928 <= _T_938;
      end
    end
    if (_T_43) begin
      if (_T_941) begin
        _T_940 <= 16'h1;
      end else begin
        _T_940 <= _T_950;
      end
    end
    if (_T_43) begin
      if (_T_953) begin
        _T_952 <= 16'h1;
      end else begin
        _T_952 <= _T_962;
      end
    end
    if (_T_43) begin
      if (_T_965) begin
        _T_964 <= 16'h1;
      end else begin
        _T_964 <= _T_974;
      end
    end
    if (_T_43) begin
      if (_T_977) begin
        _T_976 <= 16'h1;
      end else begin
        _T_976 <= _T_986;
      end
    end
    if (_T_43) begin
      if (_T_989) begin
        _T_988 <= 16'h1;
      end else begin
        _T_988 <= _T_998;
      end
    end
    if (_T_43) begin
      if (_T_1001) begin
        _T_1000 <= 16'h1;
      end else begin
        _T_1000 <= _T_1010;
      end
    end
    if (_T_43) begin
      if (_T_1013) begin
        _T_1012 <= 16'h1;
      end else begin
        _T_1012 <= _T_1022;
      end
    end
    if (_T_43) begin
      if (_T_1025) begin
        _T_1024 <= 16'h1;
      end else begin
        _T_1024 <= _T_1034;
      end
    end
    if (_T_43) begin
      if (_T_1037) begin
        _T_1036 <= 16'h1;
      end else begin
        _T_1036 <= _T_1046;
      end
    end
    if (_T_43) begin
      if (_T_1049) begin
        _T_1048 <= 16'h1;
      end else begin
        _T_1048 <= _T_1058;
      end
    end
    if (_T_43) begin
      if (_T_1061) begin
        _T_1060 <= 16'h1;
      end else begin
        _T_1060 <= _T_1070;
      end
    end
    if (_T_43) begin
      if (_T_1073) begin
        _T_1072 <= 16'h1;
      end else begin
        _T_1072 <= _T_1082;
      end
    end
    if (_T_43) begin
      if (_T_1085) begin
        _T_1084 <= 16'h1;
      end else begin
        _T_1084 <= _T_1094;
      end
    end
    if (_T_43) begin
      if (_T_1097) begin
        _T_1096 <= 16'h1;
      end else begin
        _T_1096 <= _T_1106;
      end
    end
    if (_T_43) begin
      if (_T_1109) begin
        _T_1108 <= 16'h1;
      end else begin
        _T_1108 <= _T_1118;
      end
    end
    if (_T_43) begin
      if (_T_1121) begin
        _T_1120 <= 16'h1;
      end else begin
        _T_1120 <= _T_1130;
      end
    end
    if (_T_43) begin
      if (_T_1133) begin
        _T_1132 <= 16'h1;
      end else begin
        _T_1132 <= _T_1142;
      end
    end
    if (_T_43) begin
      if (_T_1145) begin
        _T_1144 <= 16'h1;
      end else begin
        _T_1144 <= _T_1154;
      end
    end
    if (_T_43) begin
      if (_T_1157) begin
        _T_1156 <= 16'h1;
      end else begin
        _T_1156 <= _T_1166;
      end
    end
    if (_T_43) begin
      if (_T_1169) begin
        _T_1168 <= 16'h1;
      end else begin
        _T_1168 <= _T_1178;
      end
    end
    if (_T_43) begin
      if (_T_1181) begin
        _T_1180 <= 16'h1;
      end else begin
        _T_1180 <= _T_1190;
      end
    end
    if (_T_43) begin
      if (_T_1193) begin
        _T_1192 <= 16'h1;
      end else begin
        _T_1192 <= _T_1202;
      end
    end
    if (_T_43) begin
      if (_T_1205) begin
        _T_1204 <= 16'h1;
      end else begin
        _T_1204 <= _T_1214;
      end
    end
    if (_T_43) begin
      if (_T_1217) begin
        _T_1216 <= 16'h1;
      end else begin
        _T_1216 <= _T_1226;
      end
    end
    if (_T_43) begin
      if (_T_1229) begin
        _T_1228 <= 16'h1;
      end else begin
        _T_1228 <= _T_1238;
      end
    end
    if (_T_43) begin
      if (_T_1241) begin
        _T_1240 <= 16'h1;
      end else begin
        _T_1240 <= _T_1250;
      end
    end
    if (_T_43) begin
      if (_T_1253) begin
        _T_1252 <= 16'h1;
      end else begin
        _T_1252 <= _T_1262;
      end
    end
    if (_T_43) begin
      if (_T_1265) begin
        _T_1264 <= 16'h1;
      end else begin
        _T_1264 <= _T_1274;
      end
    end
    if (_T_43) begin
      if (_T_1277) begin
        _T_1276 <= 16'h1;
      end else begin
        _T_1276 <= _T_1286;
      end
    end
    if (_T_43) begin
      if (_T_1289) begin
        _T_1288 <= 16'h1;
      end else begin
        _T_1288 <= _T_1298;
      end
    end
    if (_T_43) begin
      if (_T_1301) begin
        _T_1300 <= 16'h1;
      end else begin
        _T_1300 <= _T_1310;
      end
    end
    if (_T_43) begin
      if (_T_1313) begin
        _T_1312 <= 16'h1;
      end else begin
        _T_1312 <= _T_1322;
      end
    end
    if (_T_43) begin
      if (_T_1325) begin
        _T_1324 <= 16'h1;
      end else begin
        _T_1324 <= _T_1334;
      end
    end
    if (_T_43) begin
      if (_T_1337) begin
        _T_1336 <= 16'h1;
      end else begin
        _T_1336 <= _T_1346;
      end
    end
    if (_T_43) begin
      if (_T_1349) begin
        _T_1348 <= 16'h1;
      end else begin
        _T_1348 <= _T_1358;
      end
    end
    if (_T_43) begin
      if (_T_1361) begin
        _T_1360 <= 16'h1;
      end else begin
        _T_1360 <= _T_1370;
      end
    end
    if (_T_43) begin
      if (_T_1373) begin
        _T_1372 <= 16'h1;
      end else begin
        _T_1372 <= _T_1382;
      end
    end
    if (_T_43) begin
      if (_T_1385) begin
        _T_1384 <= 16'h1;
      end else begin
        _T_1384 <= _T_1394;
      end
    end
    if (_T_43) begin
      if (_T_1397) begin
        _T_1396 <= 16'h1;
      end else begin
        _T_1396 <= _T_1406;
      end
    end
    if (_T_43) begin
      if (_T_1409) begin
        _T_1408 <= 16'h1;
      end else begin
        _T_1408 <= _T_1418;
      end
    end
    if (_T_43) begin
      if (_T_1421) begin
        _T_1420 <= 16'h1;
      end else begin
        _T_1420 <= _T_1430;
      end
    end
    if (_T_43) begin
      if (_T_1433) begin
        _T_1432 <= 16'h1;
      end else begin
        _T_1432 <= _T_1442;
      end
    end
    if (_T_43) begin
      if (_T_1445) begin
        _T_1444 <= 16'h1;
      end else begin
        _T_1444 <= _T_1454;
      end
    end
    if (_T_43) begin
      if (_T_1457) begin
        _T_1456 <= 16'h1;
      end else begin
        _T_1456 <= _T_1466;
      end
    end
    if (_T_43) begin
      if (_T_1469) begin
        _T_1468 <= 16'h1;
      end else begin
        _T_1468 <= _T_1478;
      end
    end
    if (_T_43) begin
      if (_T_1481) begin
        _T_1480 <= 16'h1;
      end else begin
        _T_1480 <= _T_1490;
      end
    end
    if (_T_43) begin
      if (_T_1493) begin
        _T_1492 <= 16'h1;
      end else begin
        _T_1492 <= _T_1502;
      end
    end
    if (_T_43) begin
      if (_T_1505) begin
        _T_1504 <= 16'h1;
      end else begin
        _T_1504 <= _T_1514;
      end
    end
    if (_T_43) begin
      if (_T_1517) begin
        _T_1516 <= 16'h1;
      end else begin
        _T_1516 <= _T_1526;
      end
    end
    if (_T_43) begin
      if (_T_1529) begin
        _T_1528 <= 16'h1;
      end else begin
        _T_1528 <= _T_1538;
      end
    end
    if (_T_43) begin
      if (_T_1541) begin
        _T_1540 <= 16'h1;
      end else begin
        _T_1540 <= _T_1550;
      end
    end
    if (_T_43) begin
      if (_T_1553) begin
        _T_1552 <= 16'h1;
      end else begin
        _T_1552 <= _T_1562;
      end
    end
    if (_T_43) begin
      if (_T_1565) begin
        _T_1564 <= 16'h1;
      end else begin
        _T_1564 <= _T_1574;
      end
    end
    if (_T_43) begin
      if (_T_1577) begin
        _T_1576 <= 16'h1;
      end else begin
        _T_1576 <= _T_1586;
      end
    end
    if (_T_43) begin
      if (_T_1589) begin
        _T_1588 <= 16'h1;
      end else begin
        _T_1588 <= _T_1598;
      end
    end
    if (_T_43) begin
      if (_T_1601) begin
        _T_1600 <= 16'h1;
      end else begin
        _T_1600 <= _T_1610;
      end
    end
    if (_T_43) begin
      if (_T_1613) begin
        _T_1612 <= 16'h1;
      end else begin
        _T_1612 <= _T_1622;
      end
    end
    if (_T_43) begin
      if (_T_1625) begin
        _T_1624 <= 16'h1;
      end else begin
        _T_1624 <= _T_1634;
      end
    end
    if (_T_43) begin
      if (_T_1637) begin
        _T_1636 <= 16'h1;
      end else begin
        _T_1636 <= _T_1646;
      end
    end
    if (_T_43) begin
      if (_T_1649) begin
        _T_1648 <= 16'h1;
      end else begin
        _T_1648 <= _T_1658;
      end
    end
    if (_T_43) begin
      if (_T_1661) begin
        _T_1660 <= 16'h1;
      end else begin
        _T_1660 <= _T_1670;
      end
    end
    if (_T_43) begin
      if (_T_1673) begin
        _T_1672 <= 16'h1;
      end else begin
        _T_1672 <= _T_1682;
      end
    end
    if (_T_43) begin
      if (_T_1685) begin
        _T_1684 <= 16'h1;
      end else begin
        _T_1684 <= _T_1694;
      end
    end
    if (_T_43) begin
      if (_T_1697) begin
        _T_1696 <= 16'h1;
      end else begin
        _T_1696 <= _T_1706;
      end
    end
    if (_T_43) begin
      if (_T_1839) begin
        _T_1838 <= 16'h1;
      end else begin
        _T_1838 <= _T_1848;
      end
    end
    if (_T_43) begin
      if (_T_1851) begin
        _T_1850 <= 16'h1;
      end else begin
        _T_1850 <= _T_1860;
      end
    end
    if (_T_43) begin
      if (_T_1863) begin
        _T_1862 <= 16'h1;
      end else begin
        _T_1862 <= _T_1872;
      end
    end
    if (_T_43) begin
      if (_T_1875) begin
        _T_1874 <= 16'h1;
      end else begin
        _T_1874 <= _T_1884;
      end
    end
    if (_T_43) begin
      if (_T_1887) begin
        _T_1886 <= 16'h1;
      end else begin
        _T_1886 <= _T_1896;
      end
    end
    if (_T_43) begin
      if (_T_1899) begin
        _T_1898 <= 16'h1;
      end else begin
        _T_1898 <= _T_1908;
      end
    end
    if (_T_43) begin
      if (_T_1911) begin
        _T_1910 <= 16'h1;
      end else begin
        _T_1910 <= _T_1920;
      end
    end
    if (_T_43) begin
      if (_T_1923) begin
        _T_1922 <= 16'h1;
      end else begin
        _T_1922 <= _T_1932;
      end
    end
    if (_T_43) begin
      if (_T_1935) begin
        _T_1934 <= 16'h1;
      end else begin
        _T_1934 <= _T_1944;
      end
    end
    if (_T_43) begin
      if (_T_1947) begin
        _T_1946 <= 16'h1;
      end else begin
        _T_1946 <= _T_1956;
      end
    end
    if (_T_43) begin
      if (_T_1959) begin
        _T_1958 <= 16'h1;
      end else begin
        _T_1958 <= _T_1968;
      end
    end
    if (_T_43) begin
      if (_T_1971) begin
        _T_1970 <= 16'h1;
      end else begin
        _T_1970 <= _T_1980;
      end
    end
    if (_T_43) begin
      if (_T_1983) begin
        _T_1982 <= 16'h1;
      end else begin
        _T_1982 <= _T_1992;
      end
    end
    if (_T_43) begin
      if (_T_1995) begin
        _T_1994 <= 16'h1;
      end else begin
        _T_1994 <= _T_2004;
      end
    end
    if (_T_43) begin
      if (_T_2007) begin
        _T_2006 <= 16'h1;
      end else begin
        _T_2006 <= _T_2016;
      end
    end
    if (_T_43) begin
      if (_T_2019) begin
        _T_2018 <= 16'h1;
      end else begin
        _T_2018 <= _T_2028;
      end
    end
    if (_T_43) begin
      if (_T_2031) begin
        _T_2030 <= 16'h1;
      end else begin
        _T_2030 <= _T_2040;
      end
    end
    if (_T_43) begin
      if (_T_2043) begin
        _T_2042 <= 16'h1;
      end else begin
        _T_2042 <= _T_2052;
      end
    end
    if (_T_43) begin
      if (_T_2055) begin
        _T_2054 <= 16'h1;
      end else begin
        _T_2054 <= _T_2064;
      end
    end
    if (_T_43) begin
      if (_T_2067) begin
        _T_2066 <= 16'h1;
      end else begin
        _T_2066 <= _T_2076;
      end
    end
    if (_T_43) begin
      if (_T_2079) begin
        _T_2078 <= 16'h1;
      end else begin
        _T_2078 <= _T_2088;
      end
    end
    if (_T_43) begin
      if (_T_2091) begin
        _T_2090 <= 16'h1;
      end else begin
        _T_2090 <= _T_2100;
      end
    end
    if (_T_43) begin
      if (_T_2103) begin
        _T_2102 <= 16'h1;
      end else begin
        _T_2102 <= _T_2112;
      end
    end
    if (_T_43) begin
      if (_T_2115) begin
        _T_2114 <= 16'h1;
      end else begin
        _T_2114 <= _T_2124;
      end
    end
    if (_T_43) begin
      if (_T_2127) begin
        _T_2126 <= 16'h1;
      end else begin
        _T_2126 <= _T_2136;
      end
    end
    if (_T_43) begin
      if (_T_2139) begin
        _T_2138 <= 16'h1;
      end else begin
        _T_2138 <= _T_2148;
      end
    end
    if (_T_43) begin
      if (_T_2151) begin
        _T_2150 <= 16'h1;
      end else begin
        _T_2150 <= _T_2160;
      end
    end
    if (_T_43) begin
      if (_T_2163) begin
        _T_2162 <= 16'h1;
      end else begin
        _T_2162 <= _T_2172;
      end
    end
    if (_T_43) begin
      if (_T_2175) begin
        _T_2174 <= 16'h1;
      end else begin
        _T_2174 <= _T_2184;
      end
    end
    if (_T_43) begin
      if (_T_2187) begin
        _T_2186 <= 16'h1;
      end else begin
        _T_2186 <= _T_2196;
      end
    end
    if (_T_43) begin
      if (_T_2199) begin
        _T_2198 <= 16'h1;
      end else begin
        _T_2198 <= _T_2208;
      end
    end
    if (_T_43) begin
      if (_T_2211) begin
        _T_2210 <= 16'h1;
      end else begin
        _T_2210 <= _T_2220;
      end
    end
    if (_T_43) begin
      if (_T_2223) begin
        _T_2222 <= 16'h1;
      end else begin
        _T_2222 <= _T_2232;
      end
    end
    if (_T_43) begin
      if (_T_2235) begin
        _T_2234 <= 16'h1;
      end else begin
        _T_2234 <= _T_2244;
      end
    end
    if (_T_43) begin
      if (_T_2247) begin
        _T_2246 <= 16'h1;
      end else begin
        _T_2246 <= _T_2256;
      end
    end
    if (_T_43) begin
      if (_T_2259) begin
        _T_2258 <= 16'h1;
      end else begin
        _T_2258 <= _T_2268;
      end
    end
    if (_T_43) begin
      if (_T_2271) begin
        _T_2270 <= 16'h1;
      end else begin
        _T_2270 <= _T_2280;
      end
    end
    if (_T_43) begin
      if (_T_2283) begin
        _T_2282 <= 16'h1;
      end else begin
        _T_2282 <= _T_2292;
      end
    end
    if (_T_43) begin
      if (_T_2295) begin
        _T_2294 <= 16'h1;
      end else begin
        _T_2294 <= _T_2304;
      end
    end
    if (_T_43) begin
      if (_T_2307) begin
        _T_2306 <= 16'h1;
      end else begin
        _T_2306 <= _T_2316;
      end
    end
    if (_T_43) begin
      if (_T_2319) begin
        _T_2318 <= 16'h1;
      end else begin
        _T_2318 <= _T_2328;
      end
    end
    if (_T_43) begin
      if (_T_2331) begin
        _T_2330 <= 16'h1;
      end else begin
        _T_2330 <= _T_2340;
      end
    end
    if (_T_43) begin
      if (_T_2343) begin
        _T_2342 <= 16'h1;
      end else begin
        _T_2342 <= _T_2352;
      end
    end
    if (_T_43) begin
      if (_T_2355) begin
        _T_2354 <= 16'h1;
      end else begin
        _T_2354 <= _T_2364;
      end
    end
    if (_T_43) begin
      if (_T_2367) begin
        _T_2366 <= 16'h1;
      end else begin
        _T_2366 <= _T_2376;
      end
    end
    if (_T_43) begin
      if (_T_2379) begin
        _T_2378 <= 16'h1;
      end else begin
        _T_2378 <= _T_2388;
      end
    end
    if (_T_43) begin
      if (_T_2391) begin
        _T_2390 <= 16'h1;
      end else begin
        _T_2390 <= _T_2400;
      end
    end
    if (_T_43) begin
      if (_T_2403) begin
        _T_2402 <= 16'h1;
      end else begin
        _T_2402 <= _T_2412;
      end
    end
    if (_T_43) begin
      if (_T_2415) begin
        _T_2414 <= 16'h1;
      end else begin
        _T_2414 <= _T_2424;
      end
    end
    if (_T_43) begin
      if (_T_2427) begin
        _T_2426 <= 16'h1;
      end else begin
        _T_2426 <= _T_2436;
      end
    end
    if (_T_43) begin
      if (_T_2439) begin
        _T_2438 <= 16'h1;
      end else begin
        _T_2438 <= _T_2448;
      end
    end
    if (_T_43) begin
      if (_T_2451) begin
        _T_2450 <= 16'h1;
      end else begin
        _T_2450 <= _T_2460;
      end
    end
    if (_T_43) begin
      if (_T_2463) begin
        _T_2462 <= 16'h1;
      end else begin
        _T_2462 <= _T_2472;
      end
    end
    if (_T_43) begin
      if (_T_2475) begin
        _T_2474 <= 16'h1;
      end else begin
        _T_2474 <= _T_2484;
      end
    end
    if (_T_43) begin
      if (_T_2487) begin
        _T_2486 <= 16'h1;
      end else begin
        _T_2486 <= _T_2496;
      end
    end
    if (_T_43) begin
      if (_T_2499) begin
        _T_2498 <= 16'h1;
      end else begin
        _T_2498 <= _T_2508;
      end
    end
    if (_T_43) begin
      if (_T_2511) begin
        _T_2510 <= 16'h1;
      end else begin
        _T_2510 <= _T_2520;
      end
    end
    if (_T_43) begin
      if (_T_2523) begin
        _T_2522 <= 16'h1;
      end else begin
        _T_2522 <= _T_2532;
      end
    end
    if (_T_43) begin
      if (_T_2535) begin
        _T_2534 <= 16'h1;
      end else begin
        _T_2534 <= _T_2544;
      end
    end
    if (_T_43) begin
      if (_T_2547) begin
        _T_2546 <= 16'h1;
      end else begin
        _T_2546 <= _T_2556;
      end
    end
    if (_T_43) begin
      if (_T_2559) begin
        _T_2558 <= 16'h1;
      end else begin
        _T_2558 <= _T_2568;
      end
    end
    if (_T_43) begin
      if (_T_2571) begin
        _T_2570 <= 16'h1;
      end else begin
        _T_2570 <= _T_2580;
      end
    end
    if (_T_43) begin
      if (_T_2583) begin
        _T_2582 <= 16'h1;
      end else begin
        _T_2582 <= _T_2592;
      end
    end
    if (_T_43) begin
      if (_T_2595) begin
        _T_2594 <= 16'h1;
      end else begin
        _T_2594 <= _T_2604;
      end
    end
    if (_T_43) begin
      if (_T_2607) begin
        _T_2606 <= 16'h1;
      end else begin
        _T_2606 <= _T_2616;
      end
    end
    if (_T_43) begin
      if (_T_2619) begin
        _T_2618 <= 16'h1;
      end else begin
        _T_2618 <= _T_2628;
      end
    end
    if (_T_43) begin
      if (_T_2631) begin
        _T_2630 <= 16'h1;
      end else begin
        _T_2630 <= _T_2640;
      end
    end
    if (_T_43) begin
      if (_T_2643) begin
        _T_2642 <= 16'h1;
      end else begin
        _T_2642 <= _T_2652;
      end
    end
    if (_T_43) begin
      if (_T_2655) begin
        _T_2654 <= 16'h1;
      end else begin
        _T_2654 <= _T_2664;
      end
    end
    if (_T_43) begin
      if (_T_2667) begin
        _T_2666 <= 16'h1;
      end else begin
        _T_2666 <= _T_2676;
      end
    end
    if (_T_43) begin
      if (_T_2679) begin
        _T_2678 <= 16'h1;
      end else begin
        _T_2678 <= _T_2688;
      end
    end
    if (_T_43) begin
      if (_T_2691) begin
        _T_2690 <= 16'h1;
      end else begin
        _T_2690 <= _T_2700;
      end
    end
    if (_T_43) begin
      if (_T_2703) begin
        _T_2702 <= 16'h1;
      end else begin
        _T_2702 <= _T_2712;
      end
    end
    if (_T_43) begin
      if (_T_2715) begin
        _T_2714 <= 16'h1;
      end else begin
        _T_2714 <= _T_2724;
      end
    end
    if (_T_43) begin
      if (_T_2727) begin
        _T_2726 <= 16'h1;
      end else begin
        _T_2726 <= _T_2736;
      end
    end
    if (_T_43) begin
      if (_T_2739) begin
        _T_2738 <= 16'h1;
      end else begin
        _T_2738 <= _T_2748;
      end
    end
    if (_T_43) begin
      if (_T_2751) begin
        _T_2750 <= 16'h1;
      end else begin
        _T_2750 <= _T_2760;
      end
    end
    if (_T_43) begin
      if (_T_2763) begin
        _T_2762 <= 16'h1;
      end else begin
        _T_2762 <= _T_2772;
      end
    end
    if (_T_43) begin
      if (_T_2775) begin
        _T_2774 <= 16'h1;
      end else begin
        _T_2774 <= _T_2784;
      end
    end
    if (_T_43) begin
      if (_T_2787) begin
        _T_2786 <= 16'h1;
      end else begin
        _T_2786 <= _T_2796;
      end
    end
    if (_T_43) begin
      if (_T_2799) begin
        _T_2798 <= 16'h1;
      end else begin
        _T_2798 <= _T_2808;
      end
    end
    if (_T_43) begin
      if (_T_2811) begin
        _T_2810 <= 16'h1;
      end else begin
        _T_2810 <= _T_2820;
      end
    end
    if (_T_43) begin
      if (_T_2823) begin
        _T_2822 <= 16'h1;
      end else begin
        _T_2822 <= _T_2832;
      end
    end
    if (_T_43) begin
      if (_T_2835) begin
        _T_2834 <= 16'h1;
      end else begin
        _T_2834 <= _T_2844;
      end
    end
    if (_T_43) begin
      if (_T_2847) begin
        _T_2846 <= 16'h1;
      end else begin
        _T_2846 <= _T_2856;
      end
    end
    if (_T_43) begin
      if (_T_2859) begin
        _T_2858 <= 16'h1;
      end else begin
        _T_2858 <= _T_2868;
      end
    end
    if (_T_43) begin
      if (_T_2871) begin
        _T_2870 <= 16'h1;
      end else begin
        _T_2870 <= _T_2880;
      end
    end
    if (_T_43) begin
      if (_T_2883) begin
        _T_2882 <= 16'h1;
      end else begin
        _T_2882 <= _T_2892;
      end
    end
    if (_T_43) begin
      if (_T_2895) begin
        _T_2894 <= 16'h1;
      end else begin
        _T_2894 <= _T_2904;
      end
    end
    if (_T_43) begin
      if (_T_2907) begin
        _T_2906 <= 16'h1;
      end else begin
        _T_2906 <= _T_2916;
      end
    end
    if (_T_43) begin
      if (_T_2919) begin
        _T_2918 <= 16'h1;
      end else begin
        _T_2918 <= _T_2928;
      end
    end
    if (_T_43) begin
      if (_T_2931) begin
        _T_2930 <= 16'h1;
      end else begin
        _T_2930 <= _T_2940;
      end
    end
    if (_T_43) begin
      if (_T_2943) begin
        _T_2942 <= 16'h1;
      end else begin
        _T_2942 <= _T_2952;
      end
    end
    if (_T_43) begin
      if (_T_2955) begin
        _T_2954 <= 16'h1;
      end else begin
        _T_2954 <= _T_2964;
      end
    end
    if (_T_43) begin
      if (_T_2967) begin
        _T_2966 <= 16'h1;
      end else begin
        _T_2966 <= _T_2976;
      end
    end
    if (_T_43) begin
      if (_T_2979) begin
        _T_2978 <= 16'h1;
      end else begin
        _T_2978 <= _T_2988;
      end
    end
    if (_T_43) begin
      if (_T_2991) begin
        _T_2990 <= 16'h1;
      end else begin
        _T_2990 <= _T_3000;
      end
    end
    if (_T_43) begin
      if (_T_3003) begin
        _T_3002 <= 16'h1;
      end else begin
        _T_3002 <= _T_3012;
      end
    end
    if (_T_43) begin
      if (_T_3015) begin
        _T_3014 <= 16'h1;
      end else begin
        _T_3014 <= _T_3024;
      end
    end
    if (_T_43) begin
      if (_T_3027) begin
        _T_3026 <= 16'h1;
      end else begin
        _T_3026 <= _T_3036;
      end
    end
    if (_T_43) begin
      if (_T_3039) begin
        _T_3038 <= 16'h1;
      end else begin
        _T_3038 <= _T_3048;
      end
    end
    if (_T_43) begin
      if (_T_3051) begin
        _T_3050 <= 16'h1;
      end else begin
        _T_3050 <= _T_3060;
      end
    end
    if (_T_43) begin
      if (_T_3063) begin
        _T_3062 <= 16'h1;
      end else begin
        _T_3062 <= _T_3072;
      end
    end
    if (_T_43) begin
      if (_T_3075) begin
        _T_3074 <= 16'h1;
      end else begin
        _T_3074 <= _T_3084;
      end
    end
    if (_T_43) begin
      if (_T_3087) begin
        _T_3086 <= 16'h1;
      end else begin
        _T_3086 <= _T_3096;
      end
    end
    if (_T_43) begin
      if (_T_3099) begin
        _T_3098 <= 16'h1;
      end else begin
        _T_3098 <= _T_3108;
      end
    end
    if (_T_43) begin
      if (_T_3111) begin
        _T_3110 <= 16'h1;
      end else begin
        _T_3110 <= _T_3120;
      end
    end
    if (_T_43) begin
      if (_T_3123) begin
        _T_3122 <= 16'h1;
      end else begin
        _T_3122 <= _T_3132;
      end
    end
    if (_T_43) begin
      if (_T_3135) begin
        _T_3134 <= 16'h1;
      end else begin
        _T_3134 <= _T_3144;
      end
    end
    if (_T_43) begin
      if (_T_3147) begin
        _T_3146 <= 16'h1;
      end else begin
        _T_3146 <= _T_3156;
      end
    end
    if (_T_43) begin
      if (_T_3159) begin
        _T_3158 <= 16'h1;
      end else begin
        _T_3158 <= _T_3168;
      end
    end
    if (_T_43) begin
      if (_T_3171) begin
        _T_3170 <= 16'h1;
      end else begin
        _T_3170 <= _T_3180;
      end
    end
    if (_T_43) begin
      if (_T_3183) begin
        _T_3182 <= 16'h1;
      end else begin
        _T_3182 <= _T_3192;
      end
    end
    if (_T_43) begin
      if (_T_3195) begin
        _T_3194 <= 16'h1;
      end else begin
        _T_3194 <= _T_3204;
      end
    end
    if (_T_43) begin
      if (_T_3207) begin
        _T_3206 <= 16'h1;
      end else begin
        _T_3206 <= _T_3216;
      end
    end
    if (_T_43) begin
      if (_T_3219) begin
        _T_3218 <= 16'h1;
      end else begin
        _T_3218 <= _T_3228;
      end
    end
    if (_T_43) begin
      if (_T_3231) begin
        _T_3230 <= 16'h1;
      end else begin
        _T_3230 <= _T_3240;
      end
    end
    if (_T_43) begin
      if (_T_3243) begin
        _T_3242 <= 16'h1;
      end else begin
        _T_3242 <= _T_3252;
      end
    end
    if (_T_43) begin
      if (_T_3255) begin
        _T_3254 <= 16'h1;
      end else begin
        _T_3254 <= _T_3264;
      end
    end
    if (_T_43) begin
      if (_T_3267) begin
        _T_3266 <= 16'h1;
      end else begin
        _T_3266 <= _T_3276;
      end
    end
    if (_T_43) begin
      if (_T_3279) begin
        _T_3278 <= 16'h1;
      end else begin
        _T_3278 <= _T_3288;
      end
    end
    if (_T_43) begin
      if (_T_3291) begin
        _T_3290 <= 16'h1;
      end else begin
        _T_3290 <= _T_3300;
      end
    end
    if (_T_43) begin
      if (_T_3303) begin
        _T_3302 <= 16'h1;
      end else begin
        _T_3302 <= _T_3312;
      end
    end
    if (_T_43) begin
      if (_T_3315) begin
        _T_3314 <= 16'h1;
      end else begin
        _T_3314 <= _T_3324;
      end
    end
    if (_T_43) begin
      if (_T_3327) begin
        _T_3326 <= 16'h1;
      end else begin
        _T_3326 <= _T_3336;
      end
    end
    if (_T_43) begin
      if (_T_3339) begin
        _T_3338 <= 16'h1;
      end else begin
        _T_3338 <= _T_3348;
      end
    end
    if (_T_43) begin
      if (_T_3351) begin
        _T_3350 <= 16'h1;
      end else begin
        _T_3350 <= _T_3360;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_529 & _T_41) begin
          $fwrite(32'h80000002,"Assertion failed: DriveInterruptType.%d not supported yet\n    at Interrupts.scala:201 assert(false.B, \"DriveInterruptType.%%d not supported yet\", drive_interrupt_type)\n",_T_30);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_529 & _T_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_549 & _T_41) begin
          $fwrite(32'h80000002,"Assertion failed: DriveInterruptType.%d not supported yet\n    at InterruptDriver.scala:83 assert(false.B, \"DriveInterruptType.%%d not supported yet\", drive_interrupt_type)\n",_T_42);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_549 & _T_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
