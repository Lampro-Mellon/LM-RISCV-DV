//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_93(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input  [1:0]  _EVAL_1,
  output        _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [29:0] _EVAL_5,
  input  [2:0]  _EVAL_6,
  output [31:0] _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  output [1:0]  _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  output        _EVAL_13,
  output        _EVAL_14,
  input  [31:0] _EVAL_15,
  output [1:0]  _EVAL_16,
  input  [2:0]  _EVAL_17,
  input         _EVAL_18,
  input  [1:0]  _EVAL_19,
  output        _EVAL_20,
  input         _EVAL_21,
  output        _EVAL_22,
  output        _EVAL_23,
  output        _EVAL_24,
  output [2:0]  _EVAL_25,
  input  [31:0] _EVAL_26,
  input         _EVAL_27,
  input  [2:0]  _EVAL_28,
  output        _EVAL_29,
  output [31:0] _EVAL_30,
  input  [3:0]  _EVAL_31,
  output [2:0]  _EVAL_32,
  output        _EVAL_33,
  input         _EVAL_34,
  output [2:0]  _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  output [3:0]  _EVAL_38,
  output [29:0] _EVAL_39,
  input         _EVAL_40,
  output [2:0]  _EVAL_41,
  output [1:0]  _EVAL_42,
  output        _EVAL_43,
  input  [1:0]  _EVAL_44,
  output        _EVAL_45,
  input  [2:0]  _EVAL_46,
  output        _EVAL_47,
  output [2:0]  _EVAL_48
);
  assign _EVAL_10 = _EVAL_19;
  assign _EVAL_25 = _EVAL_6;
  assign _EVAL_47 = _EVAL_18;
  assign _EVAL_33 = _EVAL_3;
  assign _EVAL_32 = _EVAL_28;
  assign _EVAL_7 = _EVAL_15;
  assign _EVAL_22 = _EVAL_37;
  assign _EVAL_35 = _EVAL_17;
  assign _EVAL_24 = _EVAL_36;
  assign _EVAL_16 = _EVAL_44;
  assign _EVAL_39 = _EVAL_5;
  assign _EVAL_43 = _EVAL_11;
  assign _EVAL_45 = _EVAL_9;
  assign _EVAL_23 = _EVAL_12;
  assign _EVAL_13 = _EVAL_8;
  assign _EVAL_42 = _EVAL_1;
  assign _EVAL_20 = _EVAL_4;
  assign _EVAL_48 = _EVAL_46;
  assign _EVAL_29 = _EVAL_21;
  assign _EVAL_41 = _EVAL;
  assign _EVAL_30 = _EVAL_26;
  assign _EVAL_2 = _EVAL_27;
  assign _EVAL_14 = _EVAL_0;
  assign _EVAL_38 = _EVAL_31;
endmodule
