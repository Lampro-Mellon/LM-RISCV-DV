//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_43(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  output [2:0]  _EVAL_3,
  input         _EVAL_4,
  output        _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  output        _EVAL_8,
  output [3:0]  _EVAL_9,
  input  [31:0] _EVAL_10,
  output [2:0]  _EVAL_11,
  input  [31:0] _EVAL_12,
  output        _EVAL_13,
  output        _EVAL_14,
  output [3:0]  _EVAL_15,
  output        _EVAL_16,
  output [31:0] _EVAL_17,
  input         _EVAL_18,
  output        _EVAL_19,
  output        _EVAL_20,
  output        _EVAL_21,
  input         _EVAL_22,
  output        _EVAL_23,
  input  [3:0]  _EVAL_24,
  input         _EVAL_25,
  input  [3:0]  _EVAL_26,
  output        _EVAL_27,
  output [31:0] _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  output        _EVAL_31,
  input  [2:0]  _EVAL_32,
  input  [2:0]  _EVAL_33,
  input         _EVAL_34
);
  wire [1:0] _EVAL_35;
  reg  _EVAL_36;
  reg [31:0] _RAND_0;
  reg  _EVAL_37 [0:1];
  reg [31:0] _RAND_1;
  wire  _EVAL_37__EVAL_38_data;
  wire  _EVAL_37__EVAL_38_addr;
  wire  _EVAL_37__EVAL_39_data;
  wire  _EVAL_37__EVAL_39_addr;
  wire  _EVAL_37__EVAL_39_mask;
  wire  _EVAL_37__EVAL_39_en;
  reg  _EVAL_40 [0:1];
  reg [31:0] _RAND_2;
  wire  _EVAL_40__EVAL_41_data;
  wire  _EVAL_40__EVAL_41_addr;
  wire  _EVAL_40__EVAL_42_data;
  wire  _EVAL_40__EVAL_42_addr;
  wire  _EVAL_40__EVAL_42_mask;
  wire  _EVAL_40__EVAL_42_en;
  reg [2:0] _EVAL_43 [0:1];
  reg [31:0] _RAND_3;
  wire [2:0] _EVAL_43__EVAL_44_data;
  wire  _EVAL_43__EVAL_44_addr;
  wire [2:0] _EVAL_43__EVAL_45_data;
  wire  _EVAL_43__EVAL_45_addr;
  wire  _EVAL_43__EVAL_45_mask;
  wire  _EVAL_43__EVAL_45_en;
  wire  _EVAL_46;
  reg [3:0] _EVAL_47 [0:1];
  reg [31:0] _RAND_4;
  wire [3:0] _EVAL_47__EVAL_48_data;
  wire  _EVAL_47__EVAL_48_addr;
  wire [3:0] _EVAL_47__EVAL_49_data;
  wire  _EVAL_47__EVAL_49_addr;
  wire  _EVAL_47__EVAL_49_mask;
  wire  _EVAL_47__EVAL_49_en;
  wire  _EVAL_50;
  reg  _EVAL_51 [0:1];
  reg [31:0] _RAND_5;
  wire  _EVAL_51__EVAL_52_data;
  wire  _EVAL_51__EVAL_52_addr;
  wire  _EVAL_51__EVAL_53_data;
  wire  _EVAL_51__EVAL_53_addr;
  wire  _EVAL_51__EVAL_53_mask;
  wire  _EVAL_51__EVAL_53_en;
  reg [31:0] _EVAL_54 [0:1];
  reg [31:0] _RAND_6;
  wire [31:0] _EVAL_54__EVAL_55_data;
  wire  _EVAL_54__EVAL_55_addr;
  wire [31:0] _EVAL_54__EVAL_56_data;
  wire  _EVAL_54__EVAL_56_addr;
  wire  _EVAL_54__EVAL_56_mask;
  wire  _EVAL_54__EVAL_56_en;
  reg [2:0] _EVAL_57 [0:1];
  reg [31:0] _RAND_7;
  wire [2:0] _EVAL_57__EVAL_58_data;
  wire  _EVAL_57__EVAL_58_addr;
  wire [2:0] _EVAL_57__EVAL_59_data;
  wire  _EVAL_57__EVAL_59_addr;
  wire  _EVAL_57__EVAL_59_mask;
  wire  _EVAL_57__EVAL_59_en;
  wire  _EVAL_60;
  reg  _EVAL_61;
  reg [31:0] _RAND_8;
  reg  _EVAL_63;
  reg [31:0] _RAND_9;
  wire  _EVAL_64;
  reg  _EVAL_65 [0:1];
  reg [31:0] _RAND_10;
  wire  _EVAL_65__EVAL_66_data;
  wire  _EVAL_65__EVAL_66_addr;
  wire  _EVAL_65__EVAL_67_data;
  wire  _EVAL_65__EVAL_67_addr;
  wire  _EVAL_65__EVAL_67_mask;
  wire  _EVAL_65__EVAL_67_en;
  wire [1:0] _EVAL_68;
  wire  _EVAL_69;
  reg [31:0] _EVAL_71 [0:1];
  reg [31:0] _RAND_11;
  wire [31:0] _EVAL_71__EVAL_72_data;
  wire  _EVAL_71__EVAL_72_addr;
  wire [31:0] _EVAL_71__EVAL_73_data;
  wire  _EVAL_71__EVAL_73_addr;
  wire  _EVAL_71__EVAL_73_mask;
  wire  _EVAL_71__EVAL_73_en;
  reg  _EVAL_74 [0:1];
  reg [31:0] _RAND_12;
  wire  _EVAL_74__EVAL_75_data;
  wire  _EVAL_74__EVAL_75_addr;
  wire  _EVAL_74__EVAL_76_data;
  wire  _EVAL_74__EVAL_76_addr;
  wire  _EVAL_74__EVAL_76_mask;
  wire  _EVAL_74__EVAL_76_en;
  wire  _EVAL_78;
  reg  _EVAL_79 [0:1];
  reg [31:0] _RAND_13;
  wire  _EVAL_79__EVAL_80_data;
  wire  _EVAL_79__EVAL_80_addr;
  wire  _EVAL_79__EVAL_81_data;
  wire  _EVAL_79__EVAL_81_addr;
  wire  _EVAL_79__EVAL_81_mask;
  wire  _EVAL_79__EVAL_81_en;
  reg  _EVAL_82 [0:1];
  reg [31:0] _RAND_14;
  wire  _EVAL_82__EVAL_83_data;
  wire  _EVAL_82__EVAL_83_addr;
  wire  _EVAL_82__EVAL_84_data;
  wire  _EVAL_82__EVAL_84_addr;
  wire  _EVAL_82__EVAL_84_mask;
  wire  _EVAL_82__EVAL_84_en;
  wire  _EVAL_85;
  reg [3:0] _EVAL_86 [0:1];
  reg [31:0] _RAND_15;
  wire [3:0] _EVAL_86__EVAL_87_data;
  wire  _EVAL_86__EVAL_87_addr;
  wire [3:0] _EVAL_86__EVAL_88_data;
  wire  _EVAL_86__EVAL_88_addr;
  wire  _EVAL_86__EVAL_88_mask;
  wire  _EVAL_86__EVAL_88_en;
  reg  _EVAL_89 [0:1];
  reg [31:0] _RAND_16;
  wire  _EVAL_89__EVAL_90_data;
  wire  _EVAL_89__EVAL_90_addr;
  wire  _EVAL_89__EVAL_91_data;
  wire  _EVAL_89__EVAL_91_addr;
  wire  _EVAL_89__EVAL_91_mask;
  wire  _EVAL_89__EVAL_91_en;
  reg  _EVAL_92 [0:1];
  reg [31:0] _RAND_17;
  wire  _EVAL_92__EVAL_93_data;
  wire  _EVAL_92__EVAL_93_addr;
  wire  _EVAL_92__EVAL_94_data;
  wire  _EVAL_92__EVAL_94_addr;
  wire  _EVAL_92__EVAL_94_mask;
  wire  _EVAL_92__EVAL_94_en;
  wire  _EVAL_95;
  wire  _EVAL_96;
  assign _EVAL_37__EVAL_38_addr = _EVAL_61;
  assign _EVAL_37__EVAL_38_data = _EVAL_37[_EVAL_37__EVAL_38_addr];
  assign _EVAL_37__EVAL_39_data = _EVAL_30;
  assign _EVAL_37__EVAL_39_addr = _EVAL_63;
  assign _EVAL_37__EVAL_39_mask = 1'h1;
  assign _EVAL_37__EVAL_39_en = _EVAL_31 & _EVAL_0;
  assign _EVAL_40__EVAL_41_addr = _EVAL_61;
  assign _EVAL_40__EVAL_41_data = _EVAL_40[_EVAL_40__EVAL_41_addr];
  assign _EVAL_40__EVAL_42_data = _EVAL_34;
  assign _EVAL_40__EVAL_42_addr = _EVAL_63;
  assign _EVAL_40__EVAL_42_mask = 1'h1;
  assign _EVAL_40__EVAL_42_en = _EVAL_31 & _EVAL_0;
  assign _EVAL_43__EVAL_44_addr = _EVAL_61;
  assign _EVAL_43__EVAL_44_data = _EVAL_43[_EVAL_43__EVAL_44_addr];
  assign _EVAL_43__EVAL_45_data = _EVAL_33;
  assign _EVAL_43__EVAL_45_addr = _EVAL_63;
  assign _EVAL_43__EVAL_45_mask = 1'h1;
  assign _EVAL_43__EVAL_45_en = _EVAL_31 & _EVAL_0;
  assign _EVAL_47__EVAL_48_addr = _EVAL_61;
  assign _EVAL_47__EVAL_48_data = _EVAL_47[_EVAL_47__EVAL_48_addr];
  assign _EVAL_47__EVAL_49_data = _EVAL_24;
  assign _EVAL_47__EVAL_49_addr = _EVAL_63;
  assign _EVAL_47__EVAL_49_mask = 1'h1;
  assign _EVAL_47__EVAL_49_en = _EVAL_31 & _EVAL_0;
  assign _EVAL_51__EVAL_52_addr = _EVAL_61;
  assign _EVAL_51__EVAL_52_data = _EVAL_51[_EVAL_51__EVAL_52_addr];
  assign _EVAL_51__EVAL_53_data = _EVAL_6;
  assign _EVAL_51__EVAL_53_addr = _EVAL_63;
  assign _EVAL_51__EVAL_53_mask = 1'h1;
  assign _EVAL_51__EVAL_53_en = _EVAL_31 & _EVAL_0;
  assign _EVAL_54__EVAL_55_addr = _EVAL_61;
  assign _EVAL_54__EVAL_55_data = _EVAL_54[_EVAL_54__EVAL_55_addr];
  assign _EVAL_54__EVAL_56_data = _EVAL_12;
  assign _EVAL_54__EVAL_56_addr = _EVAL_63;
  assign _EVAL_54__EVAL_56_mask = 1'h1;
  assign _EVAL_54__EVAL_56_en = _EVAL_31 & _EVAL_0;
  assign _EVAL_57__EVAL_58_addr = _EVAL_61;
  assign _EVAL_57__EVAL_58_data = _EVAL_57[_EVAL_57__EVAL_58_addr];
  assign _EVAL_57__EVAL_59_data = _EVAL_32;
  assign _EVAL_57__EVAL_59_addr = _EVAL_63;
  assign _EVAL_57__EVAL_59_mask = 1'h1;
  assign _EVAL_57__EVAL_59_en = _EVAL_31 & _EVAL_0;
  assign _EVAL_65__EVAL_66_addr = _EVAL_61;
  assign _EVAL_65__EVAL_66_data = _EVAL_65[_EVAL_65__EVAL_66_addr];
  assign _EVAL_65__EVAL_67_data = _EVAL_1;
  assign _EVAL_65__EVAL_67_addr = _EVAL_63;
  assign _EVAL_65__EVAL_67_mask = 1'h1;
  assign _EVAL_65__EVAL_67_en = _EVAL_31 & _EVAL_0;
  assign _EVAL_71__EVAL_72_addr = _EVAL_61;
  assign _EVAL_71__EVAL_72_data = _EVAL_71[_EVAL_71__EVAL_72_addr];
  assign _EVAL_71__EVAL_73_data = _EVAL_10;
  assign _EVAL_71__EVAL_73_addr = _EVAL_63;
  assign _EVAL_71__EVAL_73_mask = 1'h1;
  assign _EVAL_71__EVAL_73_en = _EVAL_31 & _EVAL_0;
  assign _EVAL_74__EVAL_75_addr = _EVAL_61;
  assign _EVAL_74__EVAL_75_data = _EVAL_74[_EVAL_74__EVAL_75_addr];
  assign _EVAL_74__EVAL_76_data = _EVAL_7;
  assign _EVAL_74__EVAL_76_addr = _EVAL_63;
  assign _EVAL_74__EVAL_76_mask = 1'h1;
  assign _EVAL_74__EVAL_76_en = _EVAL_31 & _EVAL_0;
  assign _EVAL_79__EVAL_80_addr = _EVAL_61;
  assign _EVAL_79__EVAL_80_data = _EVAL_79[_EVAL_79__EVAL_80_addr];
  assign _EVAL_79__EVAL_81_data = _EVAL;
  assign _EVAL_79__EVAL_81_addr = _EVAL_63;
  assign _EVAL_79__EVAL_81_mask = 1'h1;
  assign _EVAL_79__EVAL_81_en = _EVAL_31 & _EVAL_0;
  assign _EVAL_82__EVAL_83_addr = _EVAL_61;
  assign _EVAL_82__EVAL_83_data = _EVAL_82[_EVAL_82__EVAL_83_addr];
  assign _EVAL_82__EVAL_84_data = _EVAL_4;
  assign _EVAL_82__EVAL_84_addr = _EVAL_63;
  assign _EVAL_82__EVAL_84_mask = 1'h1;
  assign _EVAL_82__EVAL_84_en = _EVAL_31 & _EVAL_0;
  assign _EVAL_86__EVAL_87_addr = _EVAL_61;
  assign _EVAL_86__EVAL_87_data = _EVAL_86[_EVAL_86__EVAL_87_addr];
  assign _EVAL_86__EVAL_88_data = _EVAL_26;
  assign _EVAL_86__EVAL_88_addr = _EVAL_63;
  assign _EVAL_86__EVAL_88_mask = 1'h1;
  assign _EVAL_86__EVAL_88_en = _EVAL_31 & _EVAL_0;
  assign _EVAL_89__EVAL_90_addr = _EVAL_61;
  assign _EVAL_89__EVAL_90_data = _EVAL_89[_EVAL_89__EVAL_90_addr];
  assign _EVAL_89__EVAL_91_data = _EVAL_22;
  assign _EVAL_89__EVAL_91_addr = _EVAL_63;
  assign _EVAL_89__EVAL_91_mask = 1'h1;
  assign _EVAL_89__EVAL_91_en = _EVAL_31 & _EVAL_0;
  assign _EVAL_92__EVAL_93_addr = _EVAL_61;
  assign _EVAL_92__EVAL_93_data = _EVAL_92[_EVAL_92__EVAL_93_addr];
  assign _EVAL_92__EVAL_94_data = _EVAL_18;
  assign _EVAL_92__EVAL_94_addr = _EVAL_63;
  assign _EVAL_92__EVAL_94_mask = 1'h1;
  assign _EVAL_92__EVAL_94_en = _EVAL_31 & _EVAL_0;
  assign _EVAL_64 = _EVAL_95 & _EVAL_96;
  assign _EVAL_14 = _EVAL_51__EVAL_52_data;
  assign _EVAL_5 = _EVAL_37__EVAL_38_data;
  assign _EVAL_27 = _EVAL_40__EVAL_41_data;
  assign _EVAL_69 = _EVAL_68[0];
  assign _EVAL_17 = _EVAL_71__EVAL_72_data;
  assign _EVAL_8 = _EVAL_89__EVAL_90_data;
  assign _EVAL_16 = _EVAL_74__EVAL_75_data;
  assign _EVAL_46 = _EVAL_29 & _EVAL_23;
  assign _EVAL_96 = ~_EVAL_36;
  assign _EVAL_15 = _EVAL_47__EVAL_48_data;
  assign _EVAL_9 = _EVAL_86__EVAL_87_data;
  assign _EVAL_31 = ~_EVAL_60;
  assign _EVAL_13 = _EVAL_82__EVAL_83_data;
  assign _EVAL_20 = _EVAL_65__EVAL_66_data;
  assign _EVAL_78 = _EVAL_35[0];
  assign _EVAL_21 = _EVAL_79__EVAL_80_data;
  assign _EVAL_3 = _EVAL_57__EVAL_58_data;
  assign _EVAL_11 = _EVAL_43__EVAL_44_data;
  assign _EVAL_60 = _EVAL_95 & _EVAL_36;
  assign _EVAL_68 = _EVAL_63 + 1'h1;
  assign _EVAL_19 = _EVAL_92__EVAL_93_data;
  assign _EVAL_85 = _EVAL_31 & _EVAL_0;
  assign _EVAL_95 = _EVAL_63 == _EVAL_61;
  assign _EVAL_35 = _EVAL_61 + 1'h1;
  assign _EVAL_23 = ~_EVAL_64;
  assign _EVAL_28 = _EVAL_54__EVAL_55_data;
  assign _EVAL_50 = _EVAL_85 != _EVAL_46;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_36 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_37[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_40[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_43[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_47[initvar] = _RAND_4[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_51[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_54[initvar] = _RAND_6[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_57[initvar] = _RAND_7[2:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_61 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_63 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_65[initvar] = _RAND_10[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_11 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_71[initvar] = _RAND_11[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_74[initvar] = _RAND_12[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_13 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_79[initvar] = _RAND_13[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_14 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_82[initvar] = _RAND_14[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_15 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_86[initvar] = _RAND_15[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_16 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_89[initvar] = _RAND_16[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_17 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_92[initvar] = _RAND_17[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_2) begin
    if (_EVAL_25) begin
      _EVAL_36 <= 1'h0;
    end else if (_EVAL_50) begin
      _EVAL_36 <= _EVAL_85;
    end
    if(_EVAL_37__EVAL_39_en & _EVAL_37__EVAL_39_mask) begin
      _EVAL_37[_EVAL_37__EVAL_39_addr] <= _EVAL_37__EVAL_39_data;
    end
    if(_EVAL_40__EVAL_42_en & _EVAL_40__EVAL_42_mask) begin
      _EVAL_40[_EVAL_40__EVAL_42_addr] <= _EVAL_40__EVAL_42_data;
    end
    if(_EVAL_43__EVAL_45_en & _EVAL_43__EVAL_45_mask) begin
      _EVAL_43[_EVAL_43__EVAL_45_addr] <= _EVAL_43__EVAL_45_data;
    end
    if(_EVAL_47__EVAL_49_en & _EVAL_47__EVAL_49_mask) begin
      _EVAL_47[_EVAL_47__EVAL_49_addr] <= _EVAL_47__EVAL_49_data;
    end
    if(_EVAL_51__EVAL_53_en & _EVAL_51__EVAL_53_mask) begin
      _EVAL_51[_EVAL_51__EVAL_53_addr] <= _EVAL_51__EVAL_53_data;
    end
    if(_EVAL_54__EVAL_56_en & _EVAL_54__EVAL_56_mask) begin
      _EVAL_54[_EVAL_54__EVAL_56_addr] <= _EVAL_54__EVAL_56_data;
    end
    if(_EVAL_57__EVAL_59_en & _EVAL_57__EVAL_59_mask) begin
      _EVAL_57[_EVAL_57__EVAL_59_addr] <= _EVAL_57__EVAL_59_data;
    end
    if (_EVAL_25) begin
      _EVAL_61 <= 1'h0;
    end else if (_EVAL_46) begin
      _EVAL_61 <= _EVAL_78;
    end
    if (_EVAL_25) begin
      _EVAL_63 <= 1'h0;
    end else if (_EVAL_85) begin
      _EVAL_63 <= _EVAL_69;
    end
    if(_EVAL_65__EVAL_67_en & _EVAL_65__EVAL_67_mask) begin
      _EVAL_65[_EVAL_65__EVAL_67_addr] <= _EVAL_65__EVAL_67_data;
    end
    if(_EVAL_71__EVAL_73_en & _EVAL_71__EVAL_73_mask) begin
      _EVAL_71[_EVAL_71__EVAL_73_addr] <= _EVAL_71__EVAL_73_data;
    end
    if(_EVAL_74__EVAL_76_en & _EVAL_74__EVAL_76_mask) begin
      _EVAL_74[_EVAL_74__EVAL_76_addr] <= _EVAL_74__EVAL_76_data;
    end
    if(_EVAL_79__EVAL_81_en & _EVAL_79__EVAL_81_mask) begin
      _EVAL_79[_EVAL_79__EVAL_81_addr] <= _EVAL_79__EVAL_81_data;
    end
    if(_EVAL_82__EVAL_84_en & _EVAL_82__EVAL_84_mask) begin
      _EVAL_82[_EVAL_82__EVAL_84_addr] <= _EVAL_82__EVAL_84_data;
    end
    if(_EVAL_86__EVAL_88_en & _EVAL_86__EVAL_88_mask) begin
      _EVAL_86[_EVAL_86__EVAL_88_addr] <= _EVAL_86__EVAL_88_data;
    end
    if(_EVAL_89__EVAL_91_en & _EVAL_89__EVAL_91_mask) begin
      _EVAL_89[_EVAL_89__EVAL_91_addr] <= _EVAL_89__EVAL_91_data;
    end
    if(_EVAL_92__EVAL_94_en & _EVAL_92__EVAL_94_mask) begin
      _EVAL_92[_EVAL_92__EVAL_94_addr] <= _EVAL_92__EVAL_94_data;
    end
  end
endmodule
