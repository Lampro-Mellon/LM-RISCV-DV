//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_42_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [1:0]  _EVAL_3,
  input  [3:0]  _EVAL_4,
  input         _EVAL_5,
  input  [3:0]  _EVAL_6,
  input  [31:0] _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input  [3:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15
);
  reg [2:0] _EVAL_16;
  reg [31:0] _RAND_0;
  wire [31:0] _EVAL_17;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire [32:0] _EVAL_25;
  wire  _EVAL_26;
  wire [32:0] _EVAL_27;
  wire [7:0] _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire [31:0] _EVAL_31;
  wire [1:0] _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire [31:0] _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire [3:0] _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire [32:0] _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire [5:0] _EVAL_66;
  reg [3:0] _EVAL_67;
  reg [31:0] _RAND_1;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire [6:0] _EVAL_75;
  wire [32:0] _EVAL_76;
  wire [32:0] _EVAL_77;
  wire [31:0] _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire [1:0] _EVAL_84;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire [3:0] _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  reg [2:0] _EVAL_92;
  reg [31:0] _RAND_2;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire [5:0] _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire [31:0] _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire [6:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire [32:0] _EVAL_107;
  reg [1:0] _EVAL_108;
  reg [31:0] _RAND_3;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  reg [5:0] _EVAL_123;
  reg [31:0] _RAND_4;
  wire [5:0] _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_131;
  wire [32:0] _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  reg  _EVAL_143;
  reg [31:0] _RAND_5;
  wire [1:0] _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire [32:0] _EVAL_148;
  wire  _EVAL_149;
  wire [7:0] _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  reg [5:0] _EVAL_157;
  reg [31:0] _RAND_6;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire [32:0] _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire [6:0] _EVAL_166;
  wire  _EVAL_167;
  wire [1:0] _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire [32:0] _EVAL_172;
  wire  _EVAL_173;
  reg [5:0] _EVAL_174;
  reg [31:0] _RAND_7;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire [31:0] _EVAL_186;
  wire [32:0] _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  reg  _EVAL_194;
  reg [31:0] _RAND_8;
  wire [32:0] _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire [32:0] _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire [32:0] _EVAL_214;
  wire [32:0] _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire [22:0] _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire [22:0] _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  reg  _EVAL_232;
  reg [31:0] _RAND_9;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire [32:0] _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire [5:0] _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire [3:0] _EVAL_251;
  reg  _EVAL_252;
  reg [31:0] _RAND_10;
  wire [7:0] _EVAL_253;
  wire [31:0] _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire [6:0] _EVAL_257;
  wire  _EVAL_258;
  wire [32:0] _EVAL_259;
  reg [31:0] _EVAL_260;
  reg [31:0] _RAND_11;
  wire  _EVAL_261;
  wire [1:0] _EVAL_262;
  wire  _EVAL_263;
  wire [32:0] _EVAL_264;
  wire [3:0] _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire [5:0] _EVAL_268;
  reg [31:0] _EVAL_269;
  reg [31:0] _RAND_12;
  reg [5:0] _EVAL_270;
  reg [31:0] _RAND_13;
  reg [3:0] _EVAL_271;
  reg [31:0] _RAND_14;
  wire [5:0] _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire [7:0] _EVAL_276;
  wire  _EVAL_277;
  wire [32:0] _EVAL_278;
  wire  _EVAL_279;
  wire [31:0] _EVAL_280;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_71 = ~_EVAL_70;
  assign _EVAL_200 = _EVAL_46 & _EVAL_86;
  assign _EVAL_33 = _EVAL_262 | 2'h1;
  assign _EVAL_205 = ~_EVAL_232;
  assign _EVAL_176 = _EVAL_5 == _EVAL_194;
  assign _EVAL_140 = _EVAL_3 == _EVAL_108;
  assign _EVAL_220 = _EVAL_6 <= 4'h6;
  assign _EVAL_169 = ~_EVAL_226;
  assign _EVAL_285 = ~_EVAL_113;
  assign _EVAL_198 = ~_EVAL_203;
  assign _EVAL_242 = _EVAL_276[7:2];
  assign _EVAL_254 = _EVAL_161[31:0];
  assign _EVAL_90 = _EVAL_10 == 3'h2;
  assign _EVAL_167 = _EVAL_4 >= 4'h2;
  assign _EVAL_263 = _EVAL_251 == 4'h0;
  assign _EVAL_64 = _EVAL_22 & _EVAL_261;
  assign _EVAL_21 = ~_EVAL_43;
  assign _EVAL_203 = _EVAL_69 | _EVAL_0;
  assign _EVAL_117 = _EVAL_154 | _EVAL_0;
  assign _EVAL_60 = ~_EVAL_44;
  assign _EVAL_91 = ~_EVAL_233;
  assign _EVAL_73 = _EVAL_275 & _EVAL_81;
  assign _EVAL_160 = ~_EVAL_206;
  assign _EVAL_49 = _EVAL_105 | _EVAL_81;
  assign _EVAL_26 = _EVAL_10 == 3'h0;
  assign _EVAL_240 = $signed(_EVAL_58) == 33'sh0;
  assign _EVAL_207 = $signed(_EVAL_278) & -33'sh1000;
  assign _EVAL_251 = ~_EVAL_12;
  assign _EVAL_97 = _EVAL_196 | _EVAL_216;
  assign _EVAL_291 = ~_EVAL_136;
  assign _EVAL_23 = _EVAL_220 & _EVAL_228;
  assign _EVAL_65 = ~_EVAL_115;
  assign _EVAL_69 = _EVAL_7 == _EVAL_269;
  assign _EVAL_83 = $signed(_EVAL_148) == 33'sh0;
  assign _EVAL_189 = ~_EVAL_110;
  assign _EVAL_126 = _EVAL_101 | _EVAL_0;
  assign _EVAL_289 = plusarg_reader_out == 32'h0;
  assign _EVAL_208 = _EVAL_275 & _EVAL_49;
  assign _EVAL_245 = ~_EVAL_231;
  assign _EVAL_228 = $signed(_EVAL_27) == 33'sh0;
  assign _EVAL_235 = _EVAL_199 & _EVAL_206;
  assign _EVAL_79 = ~_EVAL_283;
  assign _EVAL_80 = _EVAL_8 & _EVAL_111;
  assign _EVAL_262 = 2'h1 << _EVAL_151;
  assign _EVAL_213 = _EVAL_165 | _EVAL_232;
  assign _EVAL_233 = _EVAL_125 | _EVAL_0;
  assign _EVAL_104 = ~_EVAL_0;
  assign _EVAL_199 = _EVAL_7[1];
  assign _EVAL_44 = _EVAL_176 | _EVAL_0;
  assign _EVAL_146 = _EVAL_8 & _EVAL_102;
  assign _EVAL_19 = _EVAL_11 & _EVAL_9;
  assign _EVAL_246 = _EVAL_8 & _EVAL_274;
  assign _EVAL_149 = _EVAL_8 & _EVAL_26;
  assign _EVAL_154 = _EVAL_3 <= 2'h2;
  assign _EVAL_51 = _EVAL_8 & _EVAL_139;
  assign _EVAL_114 = _EVAL_275 & _EVAL_54;
  assign _EVAL_150 = _EVAL_218[7:0];
  assign _EVAL_30 = _EVAL_183 | _EVAL_0;
  assign _EVAL_139 = _EVAL_10 == 3'h4;
  assign _EVAL_132 = $signed(_EVAL_215) & -33'shc000;
  assign _EVAL_278 = {1'b0,$signed(_EVAL_31)};
  assign _EVAL_57 = _EVAL_213 >> _EVAL_5;
  assign _EVAL_264 = {1'b0,$signed(_EVAL_280)};
  assign _EVAL_28 = ~_EVAL_150;
  assign _EVAL_185 = _EVAL_179 & _EVAL_199;
  assign _EVAL_202 = _EVAL_59 | _EVAL_0;
  assign _EVAL_211 = _EVAL_197 | _EVAL_185;
  assign _EVAL_219 = _EVAL_163 & _EVAL_201;
  assign _EVAL_256 = _EVAL_56 | _EVAL_0;
  assign _EVAL_166 = _EVAL_123 - 6'h1;
  assign _EVAL_217 = _EVAL_2 == 3'h6;
  assign _EVAL_201 = ~_EVAL_217;
  assign _EVAL_234 = _EVAL_97 | _EVAL_0;
  assign _EVAL_152 = ~_EVAL_52;
  assign _EVAL_224 = _EVAL_8 & _EVAL_190;
  assign _EVAL_20 = _EVAL_2 == 3'h1;
  assign _EVAL_249 = _EVAL_212 & _EVAL_29;
  assign _EVAL_54 = _EVAL_243 | _EVAL_81;
  assign _EVAL_141 = _EVAL_131 | _EVAL_0;
  assign _EVAL_287 = _EVAL_179 & _EVAL_223;
  assign _EVAL_115 = _EVAL_127 | _EVAL_0;
  assign _EVAL_124 = _EVAL_103[5:0];
  assign _EVAL_120 = ~_EVAL_184;
  assign _EVAL_243 = _EVAL_229 | _EVAL_83;
  assign _EVAL_214 = _EVAL_237;
  assign _EVAL_231 = _EVAL_208 | _EVAL_0;
  assign _EVAL_147 = _EVAL_38 | _EVAL_0;
  assign _EVAL_144 = 2'h1 << _EVAL_5;
  assign _EVAL_61 = _EVAL_53 | _EVAL_0;
  assign _EVAL_36 = _EVAL_138 & _EVAL_72;
  assign _EVAL_180 = _EVAL_8 & _EVAL_285;
  assign _EVAL_248 = _EVAL == _EVAL_143;
  assign _EVAL_39 = _EVAL_19 & _EVAL_70;
  assign _EVAL_148 = _EVAL_195;
  assign _EVAL_24 = _EVAL_211 | _EVAL_99;
  assign _EVAL_158 = ~_EVAL_234;
  assign _EVAL_31 = _EVAL_7 ^ 32'h3000;
  assign _EVAL_86 = ~_EVAL_119;
  assign _EVAL_280 = _EVAL_7 ^ 32'h40000000;
  assign _EVAL_82 = ~_EVAL_30;
  assign _EVAL_192 = _EVAL_9 & _EVAL_288;
  assign _EVAL_52 = _EVAL_98 | _EVAL_0;
  assign _EVAL_268 = _EVAL_166[5:0];
  assign _EVAL_43 = _EVAL_239 | _EVAL_0;
  assign _EVAL_267 = ~_EVAL_221;
  assign _EVAL_284 = _EVAL_23 | _EVAL_249;
  assign _EVAL_175 = _EVAL_199 & _EVAL_160;
  assign _EVAL_215 = {1'b0,$signed(_EVAL_50)};
  assign _EVAL_101 = _EVAL_3 != 2'h2;
  assign _EVAL_197 = _EVAL_6 >= 4'h2;
  assign _EVAL_145 = _EVAL_10[2];
  assign _EVAL_42 = _EVAL_9 & _EVAL_71;
  assign _EVAL_179 = _EVAL_33[1];
  assign _EVAL_138 = _EVAL_33[0];
  assign _EVAL_276 = ~_EVAL_253;
  assign _EVAL_34 = _EVAL_9 & _EVAL_217;
  assign _EVAL_255 = _EVAL_9 & _EVAL_95;
  assign _EVAL_109 = ~_EVAL_145;
  assign _EVAL_212 = _EVAL_6 <= 4'h8;
  assign _EVAL_195 = $signed(_EVAL_259) & -33'sh5000;
  assign _EVAL_121 = _EVAL_167 | _EVAL_0;
  assign _EVAL_273 = _EVAL_22 | _EVAL_19;
  assign _EVAL_279 = _EVAL_45 | _EVAL_133;
  assign _EVAL_163 = _EVAL_19 & _EVAL_209;
  assign _EVAL_237 = $signed(_EVAL_187) & -33'sh2000;
  assign _EVAL_188 = ~_EVAL_121;
  assign _EVAL_177 = _EVAL_22 & _EVAL_113;
  assign _EVAL_209 = _EVAL_123 == 6'h0;
  assign _EVAL_227 = _EVAL_2 <= 3'h6;
  assign _EVAL_257 = _EVAL_270 - 6'h1;
  assign _EVAL_105 = _EVAL_173 | _EVAL_83;
  assign _EVAL_250 = _EVAL_2 == 3'h5;
  assign _EVAL_102 = _EVAL_10 == 3'h7;
  assign _EVAL_244 = _EVAL_4 == _EVAL_67;
  assign _EVAL_107 = _EVAL_207;
  assign _EVAL_238 = _EVAL_2 == 3'h0;
  assign _EVAL_290 = _EVAL_204 | _EVAL_0;
  assign _EVAL_223 = ~_EVAL_199;
  assign _EVAL_142 = $signed(_EVAL_76) == 33'sh0;
  assign _EVAL_72 = _EVAL_223 & _EVAL_206;
  assign _EVAL_230 = ~_EVAL_141;
  assign _EVAL_74 = ~_EVAL_147;
  assign _EVAL_286 = _EVAL_8 & _EVAL_90;
  assign _EVAL_78 = _EVAL_7 ^ 32'h20000000;
  assign _EVAL_38 = _EVAL_10 == _EVAL_16;
  assign _EVAL_183 = _EVAL_2 == _EVAL_92;
  assign _EVAL_122 = ~_EVAL_266;
  assign _EVAL_171 = _EVAL_263 | _EVAL_0;
  assign _EVAL_48 = _EVAL_138 & _EVAL_235;
  assign _EVAL_165 = _EVAL_168[0];
  assign _EVAL_35 = ~_EVAL_290;
  assign _EVAL_272 = _EVAL_28[7:2];
  assign _EVAL_56 = _EVAL_1 == _EVAL_252;
  assign _EVAL_283 = _EVAL_244 | _EVAL_0;
  assign _EVAL_66 = _EVAL_257[5:0];
  assign _EVAL_59 = _EVAL_247 | _EVAL_14;
  assign _EVAL_84 = _EVAL_219 ? _EVAL_144 : 2'h0;
  assign _EVAL_88 = {_EVAL_225,_EVAL_24,_EVAL_241,_EVAL_155};
  assign _EVAL_173 = _EVAL_29 | _EVAL_240;
  assign _EVAL_113 = _EVAL_270 == 6'h0;
  assign _EVAL_93 = ~_EVAL_182;
  assign _EVAL_128 = _EVAL_248 | _EVAL_0;
  assign _EVAL_241 = _EVAL_63 | _EVAL_36;
  assign _EVAL_110 = _EVAL_57 | _EVAL_0;
  assign _EVAL_170 = _EVAL_9 & _EVAL_250;
  assign _EVAL_186 = {{24'd0}, _EVAL_28};
  assign _EVAL_181 = _EVAL_138 & _EVAL_40;
  assign _EVAL_100 = _EVAL_7 & _EVAL_186;
  assign _EVAL_89 = ~_EVAL_117;
  assign _EVAL_96 = _EVAL_75[5:0];
  assign _EVAL_226 = _EVAL_279 | _EVAL_0;
  assign _EVAL_168 = _EVAL_64 ? 2'h1 : 2'h0;
  assign _EVAL_190 = _EVAL_10 == 3'h1;
  assign _EVAL_206 = _EVAL_7[0];
  assign _EVAL_216 = ~_EVAL_165;
  assign _EVAL_95 = _EVAL_2 == 3'h2;
  assign _EVAL_193 = ~_EVAL_171;
  assign _EVAL_247 = ~_EVAL_1;
  assign _EVAL_46 = _EVAL_232 | _EVAL_165;
  assign _EVAL_81 = $signed(_EVAL_214) == 33'sh0;
  assign _EVAL_94 = _EVAL_162 | _EVAL_249;
  assign _EVAL_288 = _EVAL_2 == 3'h4;
  assign _EVAL_259 = {1'b0,$signed(_EVAL_7)};
  assign _EVAL_127 = _EVAL_159 | _EVAL_249;
  assign _EVAL_182 = _EVAL_140 | _EVAL_0;
  assign _EVAL_75 = _EVAL_157 - 6'h1;
  assign _EVAL_134 = ~_EVAL_61;
  assign _EVAL_125 = _EVAL_12 == _EVAL_88;
  assign _EVAL_253 = _EVAL_222[7:0];
  assign _EVAL_62 = ~_EVAL_178;
  assign _EVAL_178 = _EVAL_227 | _EVAL_0;
  assign _EVAL_135 = ~_EVAL_256;
  assign _EVAL_17 = _EVAL_7 ^ 32'h2000000;
  assign _EVAL_265 = ~_EVAL_88;
  assign _EVAL_151 = _EVAL_6[0];
  assign _EVAL_55 = _EVAL_12 & _EVAL_265;
  assign _EVAL_204 = _EVAL_55 == 4'h0;
  assign _EVAL_221 = _EVAL_205 | _EVAL_0;
  assign _EVAL_118 = _EVAL_9 & _EVAL_20;
  assign _EVAL_111 = _EVAL_10 == 3'h6;
  assign _EVAL_70 = _EVAL_174 == 6'h0;
  assign _EVAL_22 = _EVAL_15 & _EVAL_8;
  assign _EVAL_63 = _EVAL_197 | _EVAL_287;
  assign _EVAL_98 = _EVAL_100 == 32'h0;
  assign _EVAL_87 = ~_EVAL_153;
  assign _EVAL_37 = _EVAL_8 & _EVAL_41;
  assign _EVAL_266 = _EVAL_197 | _EVAL_0;
  assign _EVAL_119 = _EVAL_84[0];
  assign _EVAL_261 = _EVAL_157 == 6'h0;
  assign _EVAL_133 = _EVAL_260 < plusarg_reader_out;
  assign _EVAL_68 = ~_EVAL_128;
  assign _EVAL_153 = _EVAL_94 | _EVAL_0;
  assign _EVAL_218 = 23'hff << _EVAL_6;
  assign _EVAL_155 = _EVAL_63 | _EVAL_181;
  assign _EVAL_225 = _EVAL_211 | _EVAL_48;
  assign _EVAL_172 = $signed(_EVAL_264) & -33'sh2000;
  assign _EVAL_136 = _EVAL_247 | _EVAL_0;
  assign _EVAL_162 = _EVAL_114 | _EVAL_23;
  assign _EVAL_58 = _EVAL_77;
  assign _EVAL_77 = $signed(_EVAL_25) & -33'sh1000000;
  assign _EVAL_191 = ~_EVAL_112;
  assign _EVAL_222 = 23'hff << _EVAL_4;
  assign _EVAL_229 = _EVAL_142 | _EVAL_240;
  assign _EVAL_239 = _EVAL_284 | _EVAL_73;
  assign _EVAL_47 = _EVAL_9 & _EVAL_238;
  assign _EVAL_40 = _EVAL_223 & _EVAL_160;
  assign _EVAL_277 = ~_EVAL_202;
  assign _EVAL_164 = ~_EVAL_5;
  assign _EVAL_53 = _EVAL_6 == _EVAL_271;
  assign _EVAL_112 = _EVAL_164 | _EVAL_0;
  assign _EVAL_196 = _EVAL_165 != _EVAL_119;
  assign _EVAL_274 = _EVAL_10 == 3'h5;
  assign _EVAL_184 = _EVAL_156 | _EVAL_0;
  assign _EVAL_41 = _EVAL_10 == 3'h3;
  assign _EVAL_29 = $signed(_EVAL_107) == 33'sh0;
  assign _EVAL_156 = _EVAL_3 == 2'h0;
  assign _EVAL_258 = _EVAL_2[0];
  assign _EVAL_27 = _EVAL_172;
  assign _EVAL_25 = {1'b0,$signed(_EVAL_17)};
  assign _EVAL_161 = _EVAL_260 + 32'h1;
  assign _EVAL_187 = {1'b0,$signed(_EVAL_78)};
  assign _EVAL_275 = _EVAL_6 <= 4'h2;
  assign _EVAL_45 = _EVAL_205 | _EVAL_289;
  assign _EVAL_99 = _EVAL_138 & _EVAL_175;
  assign _EVAL_131 = ~_EVAL_14;
  assign _EVAL_282 = ~_EVAL_126;
  assign _EVAL_50 = _EVAL_7 ^ 32'h80000000;
  assign _EVAL_103 = _EVAL_174 - 6'h1;
  assign _EVAL_76 = _EVAL_132;
  assign _EVAL_159 = _EVAL_275 & _EVAL_243;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_16 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_67 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_92 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_108 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_123 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_143 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_157 = _RAND_6[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_174 = _RAND_7[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_194 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_232 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_252 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_260 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_269 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_270 = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_271 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_13) begin
    if (_EVAL_177) begin
      _EVAL_16 <= _EVAL_10;
    end
    if (_EVAL_39) begin
      _EVAL_67 <= _EVAL_4;
    end
    if (_EVAL_39) begin
      _EVAL_92 <= _EVAL_2;
    end
    if (_EVAL_39) begin
      _EVAL_108 <= _EVAL_3;
    end
    if (_EVAL_0) begin
      _EVAL_123 <= 6'h0;
    end else if (_EVAL_19) begin
      if (_EVAL_209) begin
        if (_EVAL_258) begin
          _EVAL_123 <= _EVAL_242;
        end else begin
          _EVAL_123 <= 6'h0;
        end
      end else begin
        _EVAL_123 <= _EVAL_268;
      end
    end
    if (_EVAL_39) begin
      _EVAL_143 <= _EVAL;
    end
    if (_EVAL_0) begin
      _EVAL_157 <= 6'h0;
    end else if (_EVAL_22) begin
      if (_EVAL_261) begin
        if (_EVAL_109) begin
          _EVAL_157 <= _EVAL_272;
        end else begin
          _EVAL_157 <= 6'h0;
        end
      end else begin
        _EVAL_157 <= _EVAL_96;
      end
    end
    if (_EVAL_0) begin
      _EVAL_174 <= 6'h0;
    end else if (_EVAL_19) begin
      if (_EVAL_70) begin
        if (_EVAL_258) begin
          _EVAL_174 <= _EVAL_242;
        end else begin
          _EVAL_174 <= 6'h0;
        end
      end else begin
        _EVAL_174 <= _EVAL_124;
      end
    end
    if (_EVAL_39) begin
      _EVAL_194 <= _EVAL_5;
    end
    if (_EVAL_0) begin
      _EVAL_232 <= 1'h0;
    end else begin
      _EVAL_232 <= _EVAL_200;
    end
    if (_EVAL_39) begin
      _EVAL_252 <= _EVAL_1;
    end
    if (_EVAL_0) begin
      _EVAL_260 <= 32'h0;
    end else if (_EVAL_273) begin
      _EVAL_260 <= 32'h0;
    end else begin
      _EVAL_260 <= _EVAL_254;
    end
    if (_EVAL_177) begin
      _EVAL_269 <= _EVAL_7;
    end
    if (_EVAL_0) begin
      _EVAL_270 <= 6'h0;
    end else if (_EVAL_22) begin
      if (_EVAL_113) begin
        if (_EVAL_109) begin
          _EVAL_270 <= _EVAL_272;
        end else begin
          _EVAL_270 <= 6'h0;
        end
      end else begin
        _EVAL_270 <= _EVAL_66;
      end
    end
    if (_EVAL_177) begin
      _EVAL_271 <= _EVAL_6;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bb6972e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40c14615)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b834eea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c61f405e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2073ecb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8df11474)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32ff9a96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(671ce092)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8c1001a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dbc7f3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ed42ade)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(def11daf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ceacb6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6c64264)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc19f687)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b6cb77e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2f10fe4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c07adb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acb3216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c55f1c6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec234d87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(938c35e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c059267f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec593925)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ced67d36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(406a448)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5aa117df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e627e5bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57a8056)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(529591c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acd748ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15cd8c81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f04df650)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db39f0fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eba8b6a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(314e9901)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dda2a4b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55c208f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(757e96e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c0d5a70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c8e85f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb5bc18e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ad08a1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc6cbf5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ea8faf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77e5f6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df20f1bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9feab58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7891642e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4f7ae6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15fe3dc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea288f78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3cde5cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52ce0a1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(809e63b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa1838e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(271517d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69499c98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6116768)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2369a476)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(164cbbcf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e02f95f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4a81e98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e12f974a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4dfb4222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(109ce97c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d0e15a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25bc7447)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b893ca6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
