//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_118(
  input  [2:0]  _EVAL,
  input  [31:0] _EVAL_0,
  output        _EVAL_1,
  output [3:0]  _EVAL_2,
  input         _EVAL_3,
  output [31:0] _EVAL_4,
  input  [31:0] _EVAL_5,
  input  [2:0]  _EVAL_6,
  output [3:0]  _EVAL_7,
  output        _EVAL_8,
  output        _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input  [8:0]  _EVAL_12,
  input         _EVAL_13,
  output        _EVAL_14,
  output        _EVAL_15,
  input         _EVAL_16,
  input  [1:0]  _EVAL_17,
  output [31:0] _EVAL_18,
  input  [1:0]  _EVAL_19,
  output        _EVAL_20,
  input         _EVAL_21,
  output [8:0]  _EVAL_22,
  input  [31:0] _EVAL_23,
  input  [3:0]  _EVAL_24,
  output        _EVAL_25,
  input         _EVAL_26,
  output [2:0]  _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  output [2:0]  _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  output        _EVAL_33,
  input         _EVAL_34,
  output [31:0] _EVAL_35,
  output [6:0]  _EVAL_36,
  input         _EVAL_37
);
  wire [1:0] _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire [42:0] _EVAL_41;
  wire [42:0] _EVAL_42;
  wire [2:0] _EVAL_43;
  wire [9:0] _EVAL_44;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire [3:0] _EVAL_48;
  wire [9:0] _EVAL_50;
  wire [9:0] _EVAL_51;
  wire [9:0] _EVAL_52;
  wire  _EVAL_54;
  reg  _EVAL_55;
  reg [31:0] _RAND_0;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire [42:0] _EVAL_59;
  wire  _EVAL_60;
  wire [1:0] _EVAL_61;
  wire  _EVAL_62;
  wire [8:0] _EVAL_63;
  wire [9:0] _EVAL_64;
  wire  _EVAL_65;
  wire [9:0] _EVAL_66;
  wire [3:0] _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire [9:0] _EVAL_70;
  wire  _EVAL_71;
  wire [1:0] _EVAL_72;
  wire [42:0] _EVAL_73;
  wire [8:0] _EVAL_75;
  wire  _EVAL_77;
  wire [8:0] _EVAL_78;
  wire [8:0] _EVAL_79;
  wire [1:0] _EVAL_80;
  wire [8:0] _EVAL_81;
  wire [9:0] _EVAL_82;
  wire  _EVAL_83;
  wire [1:0] _EVAL_84;
  wire [9:0] _EVAL_85;
  wire [8:0] _EVAL_86;
  wire [1:0] _EVAL_87;
  wire [9:0] _EVAL_89;
  wire [2:0] _EVAL_90;
  wire [9:0] _EVAL_91;
  wire [8:0] _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire [9:0] _EVAL_95;
  wire  _EVAL_96;
  wire [3:0] _EVAL_97;
  wire [9:0] _EVAL_98;
  wire [3:0] _EVAL_99;
  wire [42:0] _EVAL_100;
  wire  _EVAL_101;
  wire [9:0] _EVAL_103;
  wire [3:0] _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  reg  _EVAL_107;
  reg [31:0] _RAND_1;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire [1:0] _EVAL_111;
  wire  _EVAL_112;
  wire [9:0] _EVAL_113;
  wire [9:0] _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire [1:0] _EVAL_117;
  wire  _EVAL_119;
  wire [1:0] _EVAL_121;
  reg  _EVAL_122;
  reg [31:0] _RAND_2;
  wire [3:0] _EVAL_123;
  wire [9:0] _EVAL_125;
  wire  _EVAL_126;
  wire [1:0] _EVAL_127;
  wire [2:0] _EVAL_128;
  wire [9:0] _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire [9:0] _EVAL_133;
  wire [9:0] _EVAL_134;
  reg [1:0] _EVAL_135;
  reg [31:0] _RAND_3;
  wire [9:0] _EVAL_136;
  wire [9:0] _EVAL_137;
  wire  _EVAL_138;
  wire [9:0] _EVAL_139;
  wire  _EVAL_140;
  wire [9:0] _EVAL_141;
  wire  _EVAL_142;
  wire [1:0] _EVAL_143;
  assign _EVAL_130 = _EVAL_38[0];
  assign _EVAL_94 = $signed(_EVAL_51) == 10'sh0;
  assign _EVAL_90 = _EVAL_123[3:1];
  assign _EVAL_97 = {{1'd0}, _EVAL_90};
  assign _EVAL_87 = _EVAL_67[3:2];
  assign _EVAL_133 = _EVAL_113;
  assign _EVAL_96 = _EVAL_77 ? _EVAL_101 : _EVAL_107;
  assign _EVAL_127 = _EVAL_111 & _EVAL_72;
  assign _EVAL_93 = _EVAL_71 | _EVAL_142;
  assign _EVAL_106 = _EVAL_69 | _EVAL_119;
  assign _EVAL_20 = _EVAL_3 & _EVAL_106;
  assign _EVAL_72 = ~_EVAL_135;
  assign _EVAL_33 = _EVAL_31 & _EVAL_108;
  assign _EVAL_115 = _EVAL_122 & _EVAL_28;
  assign _EVAL_63 = _EVAL_12 ^ 9'h80;
  assign _EVAL_110 = _EVAL_77 & _EVAL_31;
  assign _EVAL_18 = _EVAL_0;
  assign _EVAL_56 = _EVAL_11 | _EVAL_28;
  assign _EVAL_57 = _EVAL_38[1];
  assign _EVAL_59 = {_EVAL_10,_EVAL_19,_EVAL_17,_EVAL_29,_EVAL_34,_EVAL_16,_EVAL_5,_EVAL_32};
  assign _EVAL_142 = $signed(_EVAL_64) == 10'sh0;
  assign _EVAL_111 = {_EVAL_28,_EVAL_11};
  assign _EVAL_65 = _EVAL_80[0];
  assign _EVAL_117 = _EVAL_87 & _EVAL_61;
  assign _EVAL_69 = _EVAL_140 | _EVAL_109;
  assign _EVAL_123 = {_EVAL_127,_EVAL_28,_EVAL_11};
  assign _EVAL_82 = $signed(_EVAL_139) & 10'sh1fc;
  assign _EVAL_116 = _EVAL_77 ? _EVAL_56 : _EVAL_58;
  assign _EVAL_89 = {1'b0,$signed(_EVAL_86)};
  assign _EVAL_131 = _EVAL_77 ? _EVAL_130 : _EVAL_107;
  assign _EVAL_75 = _EVAL_12 ^ 9'h54;
  assign _EVAL_39 = $signed(_EVAL_133) == 10'sh0;
  assign _EVAL_109 = $signed(_EVAL_95) == 10'sh0;
  assign _EVAL_66 = {1'b0,$signed(_EVAL_12)};
  assign _EVAL_44 = $signed(_EVAL_89) & 10'sh1e8;
  assign _EVAL_77 = ~_EVAL_55;
  assign _EVAL_126 = $signed(_EVAL_52) == 10'sh0;
  assign _EVAL_22 = _EVAL_12;
  assign _EVAL_30 = _EVAL;
  assign _EVAL_4 = _EVAL_0;
  assign _EVAL_50 = $signed(_EVAL_134) & 10'sh180;
  assign _EVAL_129 = {1'b0,$signed(_EVAL_78)};
  assign _EVAL_71 = $signed(_EVAL_136) == 10'sh0;
  assign _EVAL_27 = _EVAL;
  assign _EVAL_103 = {1'b0,$signed(_EVAL_92)};
  assign _EVAL_80 = _EVAL_55 - _EVAL_105;
  assign _EVAL_99 = _EVAL_123 | _EVAL_97;
  assign _EVAL_2 = _EVAL_24;
  assign _EVAL_73 = _EVAL_96 ? _EVAL_59 : 43'h0;
  assign _EVAL_101 = _EVAL_130 & _EVAL_11;
  assign _EVAL_134 = {1'b0,$signed(_EVAL_63)};
  assign _EVAL_41 = {_EVAL_6,2'h0,3'h4,2'h0,_EVAL_23,1'h0};
  assign _EVAL_100 = _EVAL_73 | _EVAL_42;
  assign _EVAL_139 = {1'b0,$signed(_EVAL_75)};
  assign _EVAL_62 = _EVAL_68 | _EVAL_94;
  assign _EVAL_35 = _EVAL_100[32:1];
  assign _EVAL_8 = _EVAL_47 | _EVAL_138;
  assign _EVAL_68 = _EVAL_83 | _EVAL_126;
  assign _EVAL_70 = {1'b0,$signed(_EVAL_81)};
  assign _EVAL_98 = {1'b0,$signed(_EVAL_79)};
  assign _EVAL_25 = _EVAL_77 ? _EVAL_56 : _EVAL_58;
  assign _EVAL_40 = _EVAL_77 ? _EVAL_46 : _EVAL_122;
  assign _EVAL_113 = $signed(_EVAL_70) & 10'sh1e0;
  assign _EVAL_67 = _EVAL_104 | _EVAL_48;
  assign _EVAL_140 = _EVAL_62 | _EVAL_39;
  assign _EVAL_105 = _EVAL_31 & _EVAL_116;
  assign _EVAL_52 = _EVAL_114;
  assign _EVAL_64 = _EVAL_82;
  assign _EVAL_85 = $signed(_EVAL_129) & 10'sh100;
  assign _EVAL_42 = _EVAL_40 ? _EVAL_41 : 43'h0;
  assign _EVAL_14 = _EVAL_100[33];
  assign _EVAL_112 = _EVAL_107 & _EVAL_11;
  assign _EVAL_78 = _EVAL_12 ^ 9'h100;
  assign _EVAL_136 = _EVAL_125;
  assign _EVAL_119 = $signed(_EVAL_137) == 10'sh0;
  assign _EVAL_9 = _EVAL_3 & _EVAL_93;
  assign _EVAL_51 = _EVAL_44;
  assign _EVAL_121 = _EVAL_38 & _EVAL_111;
  assign _EVAL_38 = ~_EVAL_117;
  assign _EVAL_104 = {{1'd0}, _EVAL_43};
  assign _EVAL_58 = _EVAL_112 | _EVAL_115;
  assign _EVAL_7 = _EVAL_24;
  assign _EVAL_47 = _EVAL_106 & _EVAL_26;
  assign _EVAL_60 = _EVAL_110 & _EVAL_54;
  assign _EVAL_128 = {_EVAL_121, 1'h0};
  assign _EVAL_84 = _EVAL_121 | _EVAL_143;
  assign _EVAL_79 = _EVAL_12 ^ 9'h44;
  assign _EVAL_141 = _EVAL_91;
  assign _EVAL_91 = $signed(_EVAL_66) & 10'sh1c0;
  assign _EVAL_125 = $signed(_EVAL_103) & 10'sh1ec;
  assign _EVAL_137 = _EVAL_85;
  assign _EVAL_1 = _EVAL_31 & _EVAL_131;
  assign _EVAL_83 = $signed(_EVAL_141) == 10'sh0;
  assign _EVAL_43 = _EVAL_99[3:1];
  assign _EVAL_95 = _EVAL_50;
  assign _EVAL_81 = _EVAL_12 ^ 9'h60;
  assign _EVAL_54 = _EVAL_111 != 2'h0;
  assign _EVAL_46 = _EVAL_57 & _EVAL_28;
  assign _EVAL_114 = $signed(_EVAL_98) & 10'sh1fc;
  assign _EVAL_86 = _EVAL_12 ^ 9'h48;
  assign _EVAL_48 = {_EVAL_135, 2'h0};
  assign _EVAL_36 = _EVAL_12[6:0];
  assign _EVAL_108 = _EVAL_77 ? _EVAL_57 : _EVAL_122;
  assign _EVAL_92 = _EVAL_12 ^ 9'h40;
  assign _EVAL_61 = _EVAL_67[1:0];
  assign _EVAL_138 = _EVAL_93 & _EVAL_37;
  assign _EVAL_15 = _EVAL_100[0];
  assign _EVAL_143 = _EVAL_128[1:0];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_55 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_107 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_122 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_135 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  if (_EVAL_13) begin
    _EVAL_55 = 1'h0;
  end
  if (_EVAL_13) begin
    _EVAL_107 = 1'h0;
  end
  if (_EVAL_13) begin
    _EVAL_122 = 1'h0;
  end
  if (_EVAL_13) begin
    _EVAL_135 = 2'h3;
  end
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_21 or posedge _EVAL_13) begin
    if (_EVAL_13) begin
      _EVAL_55 <= 1'h0;
    end else if (_EVAL_110) begin
      _EVAL_55 <= 1'h0;
    end else begin
      _EVAL_55 <= _EVAL_65;
    end
  end
  always @(posedge _EVAL_21 or posedge _EVAL_13) begin
    if (_EVAL_13) begin
      _EVAL_107 <= 1'h0;
    end else if (_EVAL_77) begin
      _EVAL_107 <= _EVAL_101;
    end
  end
  always @(posedge _EVAL_21 or posedge _EVAL_13) begin
    if (_EVAL_13) begin
      _EVAL_122 <= 1'h0;
    end else if (_EVAL_77) begin
      _EVAL_122 <= _EVAL_46;
    end
  end
  always @(posedge _EVAL_21 or posedge _EVAL_13) begin
    if (_EVAL_13) begin
      _EVAL_135 <= 2'h3;
    end else if (_EVAL_60) begin
      _EVAL_135 <= _EVAL_84;
    end
  end
endmodule
