//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_29(
  input         _EVAL,
  output        _EVAL_0,
  input  [2:0]  _EVAL_1,
  output [3:0]  _EVAL_2,
  output        _EVAL_3,
  input  [3:0]  _EVAL_4,
  input         _EVAL_5,
  input  [30:0] _EVAL_6,
  output [1:0]  _EVAL_7,
  output [2:0]  _EVAL_8,
  output        _EVAL_9,
  output [2:0]  _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [31:0] _EVAL_13,
  output        _EVAL_14,
  input  [2:0]  _EVAL_15,
  input  [2:0]  _EVAL_16,
  input         _EVAL_17,
  output [2:0]  _EVAL_18,
  output        _EVAL_19,
  output [31:0] _EVAL_20,
  output [30:0] _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  output        _EVAL_24,
  output [31:0] _EVAL_25,
  output [2:0]  _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  output [1:0]  _EVAL_29,
  input  [31:0] _EVAL_30,
  input  [2:0]  _EVAL_31,
  input         _EVAL_32,
  output [2:0]  _EVAL_33,
  input         _EVAL_34
);
  wire [2:0] buffer__EVAL;
  wire [31:0] buffer__EVAL_0;
  wire  buffer__EVAL_1;
  wire [2:0] buffer__EVAL_2;
  wire  buffer__EVAL_3;
  wire [3:0] buffer__EVAL_4;
  wire [2:0] buffer__EVAL_5;
  wire [1:0] buffer__EVAL_6;
  wire  buffer__EVAL_7;
  wire  buffer__EVAL_8;
  wire  buffer__EVAL_9;
  wire  buffer__EVAL_10;
  wire  buffer__EVAL_11;
  wire  buffer__EVAL_12;
  wire  buffer__EVAL_13;
  wire [2:0] buffer__EVAL_14;
  wire [2:0] buffer__EVAL_15;
  wire [2:0] buffer__EVAL_16;
  wire  buffer__EVAL_17;
  wire [2:0] buffer__EVAL_18;
  wire [2:0] buffer__EVAL_19;
  wire [2:0] buffer__EVAL_20;
  wire  buffer__EVAL_21;
  wire [2:0] buffer__EVAL_22;
  wire  buffer__EVAL_23;
  wire  buffer__EVAL_24;
  wire  buffer__EVAL_25;
  wire [2:0] buffer__EVAL_26;
  wire  buffer__EVAL_27;
  wire [1:0] buffer__EVAL_28;
  wire  buffer__EVAL_29;
  wire  buffer__EVAL_30;
  wire [2:0] buffer__EVAL_31;
  wire  buffer__EVAL_32;
  wire [3:0] buffer__EVAL_33;
  wire [30:0] buffer__EVAL_34;
  wire [31:0] buffer__EVAL_35;
  wire  buffer__EVAL_36;
  wire [30:0] buffer__EVAL_37;
  wire  buffer__EVAL_38;
  wire [2:0] buffer__EVAL_39;
  wire [2:0] buffer__EVAL_40;
  wire  buffer__EVAL_41;
  wire  buffer__EVAL_42;
  wire [31:0] buffer__EVAL_43;
  wire  buffer__EVAL_44;
  wire  buffer__EVAL_45;
  wire [31:0] buffer__EVAL_46;
  wire  buffer__EVAL_47;
  wire  buffer__EVAL_48;
  wire [31:0] widget__EVAL;
  wire  widget__EVAL_0;
  wire [2:0] widget__EVAL_1;
  wire [31:0] widget__EVAL_2;
  wire  widget__EVAL_3;
  wire [2:0] widget__EVAL_4;
  wire  widget__EVAL_5;
  wire  widget__EVAL_6;
  wire [2:0] widget__EVAL_7;
  wire [2:0] widget__EVAL_8;
  wire [2:0] widget__EVAL_9;
  wire [2:0] widget__EVAL_10;
  wire [1:0] widget__EVAL_11;
  wire  widget__EVAL_12;
  wire  widget__EVAL_13;
  wire  widget__EVAL_14;
  wire  widget__EVAL_15;
  wire  widget__EVAL_16;
  wire  widget__EVAL_17;
  wire  widget__EVAL_18;
  wire [31:0] widget__EVAL_19;
  wire [2:0] widget__EVAL_20;
  wire [2:0] widget__EVAL_21;
  wire  widget__EVAL_22;
  wire  widget__EVAL_23;
  wire [1:0] widget__EVAL_24;
  wire [2:0] widget__EVAL_25;
  wire [2:0] widget__EVAL_26;
  wire  widget__EVAL_27;
  wire  widget__EVAL_28;
  wire [3:0] widget__EVAL_29;
  wire [2:0] widget__EVAL_30;
  wire  widget__EVAL_31;
  wire  widget__EVAL_32;
  wire [30:0] widget__EVAL_33;
  wire  widget__EVAL_34;
  wire [2:0] widget__EVAL_35;
  wire  widget__EVAL_36;
  wire [30:0] widget__EVAL_37;
  wire  widget__EVAL_38;
  wire [2:0] widget__EVAL_39;
  wire  widget__EVAL_40;
  wire  widget__EVAL_41;
  wire  widget__EVAL_42;
  wire [31:0] widget__EVAL_43;
  wire  widget__EVAL_44;
  wire [2:0] widget__EVAL_45;
  wire  widget__EVAL_46;
  wire [3:0] widget__EVAL_47;
  wire  widget__EVAL_48;
  wire [2:0] buffer_1__EVAL;
  wire [1:0] buffer_1__EVAL_0;
  wire [2:0] buffer_1__EVAL_1;
  wire [3:0] buffer_1__EVAL_2;
  wire  buffer_1__EVAL_3;
  wire [30:0] buffer_1__EVAL_4;
  wire  buffer_1__EVAL_5;
  wire [3:0] buffer_1__EVAL_6;
  wire  buffer_1__EVAL_7;
  wire [2:0] buffer_1__EVAL_8;
  wire [2:0] buffer_1__EVAL_9;
  wire  buffer_1__EVAL_10;
  wire  buffer_1__EVAL_11;
  wire  buffer_1__EVAL_12;
  wire  buffer_1__EVAL_13;
  wire  buffer_1__EVAL_14;
  wire [1:0] buffer_1__EVAL_15;
  wire [31:0] buffer_1__EVAL_16;
  wire  buffer_1__EVAL_17;
  wire [30:0] buffer_1__EVAL_18;
  wire  buffer_1__EVAL_19;
  wire [31:0] buffer_1__EVAL_20;
  wire  buffer_1__EVAL_21;
  wire [2:0] buffer_1__EVAL_22;
  wire [2:0] buffer_1__EVAL_23;
  wire [2:0] buffer_1__EVAL_24;
  wire  buffer_1__EVAL_25;
  wire  buffer_1__EVAL_26;
  wire  buffer_1__EVAL_27;
  wire [2:0] buffer_1__EVAL_28;
  wire [2:0] buffer_1__EVAL_29;
  wire [2:0] buffer_1__EVAL_30;
  wire [2:0] buffer_1__EVAL_31;
  wire  buffer_1__EVAL_32;
  wire [2:0] buffer_1__EVAL_33;
  wire  buffer_1__EVAL_34;
  wire [31:0] buffer_1__EVAL_35;
  wire  buffer_1__EVAL_36;
  wire  buffer_1__EVAL_37;
  wire  buffer_1__EVAL_38;
  wire [31:0] buffer_1__EVAL_39;
  wire [2:0] buffer_1__EVAL_40;
  wire  buffer_1__EVAL_41;
  wire  buffer_1__EVAL_42;
  wire  buffer_1__EVAL_43;
  wire  buffer_1__EVAL_44;
  wire  buffer_1__EVAL_45;
  wire  buffer_1__EVAL_46;
  wire  buffer_1__EVAL_47;
  wire [2:0] buffer_1__EVAL_48;
  wire  tl2ahb__EVAL;
  wire [31:0] tl2ahb__EVAL_0;
  wire [2:0] tl2ahb__EVAL_1;
  wire [30:0] tl2ahb__EVAL_2;
  wire  tl2ahb__EVAL_3;
  wire  tl2ahb__EVAL_4;
  wire [31:0] tl2ahb__EVAL_5;
  wire [1:0] tl2ahb__EVAL_6;
  wire  tl2ahb__EVAL_7;
  wire  tl2ahb__EVAL_8;
  wire [3:0] tl2ahb__EVAL_9;
  wire [1:0] tl2ahb__EVAL_10;
  wire [30:0] tl2ahb__EVAL_11;
  wire [2:0] tl2ahb__EVAL_12;
  wire  tl2ahb__EVAL_13;
  wire [2:0] tl2ahb__EVAL_14;
  wire  tl2ahb__EVAL_15;
  wire  tl2ahb__EVAL_16;
  wire  tl2ahb__EVAL_17;
  wire  tl2ahb__EVAL_18;
  wire  tl2ahb__EVAL_19;
  wire [2:0] tl2ahb__EVAL_20;
  wire [2:0] tl2ahb__EVAL_21;
  wire  tl2ahb__EVAL_22;
  wire  tl2ahb__EVAL_23;
  wire  tl2ahb__EVAL_24;
  wire [2:0] tl2ahb__EVAL_25;
  wire [31:0] tl2ahb__EVAL_26;
  wire [3:0] tl2ahb__EVAL_27;
  wire  tl2ahb__EVAL_28;
  wire  tl2ahb__EVAL_29;
  wire [2:0] tl2ahb__EVAL_30;
  wire [2:0] tl2ahb__EVAL_31;
  wire [2:0] tl2ahb__EVAL_32;
  wire [31:0] tl2ahb__EVAL_33;
  wire  tl2ahb__EVAL_34;
  _EVAL_24 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32),
    ._EVAL_33(buffer__EVAL_33),
    ._EVAL_34(buffer__EVAL_34),
    ._EVAL_35(buffer__EVAL_35),
    ._EVAL_36(buffer__EVAL_36),
    ._EVAL_37(buffer__EVAL_37),
    ._EVAL_38(buffer__EVAL_38),
    ._EVAL_39(buffer__EVAL_39),
    ._EVAL_40(buffer__EVAL_40),
    ._EVAL_41(buffer__EVAL_41),
    ._EVAL_42(buffer__EVAL_42),
    ._EVAL_43(buffer__EVAL_43),
    ._EVAL_44(buffer__EVAL_44),
    ._EVAL_45(buffer__EVAL_45),
    ._EVAL_46(buffer__EVAL_46),
    ._EVAL_47(buffer__EVAL_47),
    ._EVAL_48(buffer__EVAL_48)
  );
  _EVAL_26 widget (
    ._EVAL(widget__EVAL),
    ._EVAL_0(widget__EVAL_0),
    ._EVAL_1(widget__EVAL_1),
    ._EVAL_2(widget__EVAL_2),
    ._EVAL_3(widget__EVAL_3),
    ._EVAL_4(widget__EVAL_4),
    ._EVAL_5(widget__EVAL_5),
    ._EVAL_6(widget__EVAL_6),
    ._EVAL_7(widget__EVAL_7),
    ._EVAL_8(widget__EVAL_8),
    ._EVAL_9(widget__EVAL_9),
    ._EVAL_10(widget__EVAL_10),
    ._EVAL_11(widget__EVAL_11),
    ._EVAL_12(widget__EVAL_12),
    ._EVAL_13(widget__EVAL_13),
    ._EVAL_14(widget__EVAL_14),
    ._EVAL_15(widget__EVAL_15),
    ._EVAL_16(widget__EVAL_16),
    ._EVAL_17(widget__EVAL_17),
    ._EVAL_18(widget__EVAL_18),
    ._EVAL_19(widget__EVAL_19),
    ._EVAL_20(widget__EVAL_20),
    ._EVAL_21(widget__EVAL_21),
    ._EVAL_22(widget__EVAL_22),
    ._EVAL_23(widget__EVAL_23),
    ._EVAL_24(widget__EVAL_24),
    ._EVAL_25(widget__EVAL_25),
    ._EVAL_26(widget__EVAL_26),
    ._EVAL_27(widget__EVAL_27),
    ._EVAL_28(widget__EVAL_28),
    ._EVAL_29(widget__EVAL_29),
    ._EVAL_30(widget__EVAL_30),
    ._EVAL_31(widget__EVAL_31),
    ._EVAL_32(widget__EVAL_32),
    ._EVAL_33(widget__EVAL_33),
    ._EVAL_34(widget__EVAL_34),
    ._EVAL_35(widget__EVAL_35),
    ._EVAL_36(widget__EVAL_36),
    ._EVAL_37(widget__EVAL_37),
    ._EVAL_38(widget__EVAL_38),
    ._EVAL_39(widget__EVAL_39),
    ._EVAL_40(widget__EVAL_40),
    ._EVAL_41(widget__EVAL_41),
    ._EVAL_42(widget__EVAL_42),
    ._EVAL_43(widget__EVAL_43),
    ._EVAL_44(widget__EVAL_44),
    ._EVAL_45(widget__EVAL_45),
    ._EVAL_46(widget__EVAL_46),
    ._EVAL_47(widget__EVAL_47),
    ._EVAL_48(widget__EVAL_48)
  );
  _EVAL_28 buffer_1 (
    ._EVAL(buffer_1__EVAL),
    ._EVAL_0(buffer_1__EVAL_0),
    ._EVAL_1(buffer_1__EVAL_1),
    ._EVAL_2(buffer_1__EVAL_2),
    ._EVAL_3(buffer_1__EVAL_3),
    ._EVAL_4(buffer_1__EVAL_4),
    ._EVAL_5(buffer_1__EVAL_5),
    ._EVAL_6(buffer_1__EVAL_6),
    ._EVAL_7(buffer_1__EVAL_7),
    ._EVAL_8(buffer_1__EVAL_8),
    ._EVAL_9(buffer_1__EVAL_9),
    ._EVAL_10(buffer_1__EVAL_10),
    ._EVAL_11(buffer_1__EVAL_11),
    ._EVAL_12(buffer_1__EVAL_12),
    ._EVAL_13(buffer_1__EVAL_13),
    ._EVAL_14(buffer_1__EVAL_14),
    ._EVAL_15(buffer_1__EVAL_15),
    ._EVAL_16(buffer_1__EVAL_16),
    ._EVAL_17(buffer_1__EVAL_17),
    ._EVAL_18(buffer_1__EVAL_18),
    ._EVAL_19(buffer_1__EVAL_19),
    ._EVAL_20(buffer_1__EVAL_20),
    ._EVAL_21(buffer_1__EVAL_21),
    ._EVAL_22(buffer_1__EVAL_22),
    ._EVAL_23(buffer_1__EVAL_23),
    ._EVAL_24(buffer_1__EVAL_24),
    ._EVAL_25(buffer_1__EVAL_25),
    ._EVAL_26(buffer_1__EVAL_26),
    ._EVAL_27(buffer_1__EVAL_27),
    ._EVAL_28(buffer_1__EVAL_28),
    ._EVAL_29(buffer_1__EVAL_29),
    ._EVAL_30(buffer_1__EVAL_30),
    ._EVAL_31(buffer_1__EVAL_31),
    ._EVAL_32(buffer_1__EVAL_32),
    ._EVAL_33(buffer_1__EVAL_33),
    ._EVAL_34(buffer_1__EVAL_34),
    ._EVAL_35(buffer_1__EVAL_35),
    ._EVAL_36(buffer_1__EVAL_36),
    ._EVAL_37(buffer_1__EVAL_37),
    ._EVAL_38(buffer_1__EVAL_38),
    ._EVAL_39(buffer_1__EVAL_39),
    ._EVAL_40(buffer_1__EVAL_40),
    ._EVAL_41(buffer_1__EVAL_41),
    ._EVAL_42(buffer_1__EVAL_42),
    ._EVAL_43(buffer_1__EVAL_43),
    ._EVAL_44(buffer_1__EVAL_44),
    ._EVAL_45(buffer_1__EVAL_45),
    ._EVAL_46(buffer_1__EVAL_46),
    ._EVAL_47(buffer_1__EVAL_47),
    ._EVAL_48(buffer_1__EVAL_48)
  );
  _EVAL_22 tl2ahb (
    ._EVAL(tl2ahb__EVAL),
    ._EVAL_0(tl2ahb__EVAL_0),
    ._EVAL_1(tl2ahb__EVAL_1),
    ._EVAL_2(tl2ahb__EVAL_2),
    ._EVAL_3(tl2ahb__EVAL_3),
    ._EVAL_4(tl2ahb__EVAL_4),
    ._EVAL_5(tl2ahb__EVAL_5),
    ._EVAL_6(tl2ahb__EVAL_6),
    ._EVAL_7(tl2ahb__EVAL_7),
    ._EVAL_8(tl2ahb__EVAL_8),
    ._EVAL_9(tl2ahb__EVAL_9),
    ._EVAL_10(tl2ahb__EVAL_10),
    ._EVAL_11(tl2ahb__EVAL_11),
    ._EVAL_12(tl2ahb__EVAL_12),
    ._EVAL_13(tl2ahb__EVAL_13),
    ._EVAL_14(tl2ahb__EVAL_14),
    ._EVAL_15(tl2ahb__EVAL_15),
    ._EVAL_16(tl2ahb__EVAL_16),
    ._EVAL_17(tl2ahb__EVAL_17),
    ._EVAL_18(tl2ahb__EVAL_18),
    ._EVAL_19(tl2ahb__EVAL_19),
    ._EVAL_20(tl2ahb__EVAL_20),
    ._EVAL_21(tl2ahb__EVAL_21),
    ._EVAL_22(tl2ahb__EVAL_22),
    ._EVAL_23(tl2ahb__EVAL_23),
    ._EVAL_24(tl2ahb__EVAL_24),
    ._EVAL_25(tl2ahb__EVAL_25),
    ._EVAL_26(tl2ahb__EVAL_26),
    ._EVAL_27(tl2ahb__EVAL_27),
    ._EVAL_28(tl2ahb__EVAL_28),
    ._EVAL_29(tl2ahb__EVAL_29),
    ._EVAL_30(tl2ahb__EVAL_30),
    ._EVAL_31(tl2ahb__EVAL_31),
    ._EVAL_32(tl2ahb__EVAL_32),
    ._EVAL_33(tl2ahb__EVAL_33),
    ._EVAL_34(tl2ahb__EVAL_34)
  );
  assign _EVAL_3 = buffer_1__EVAL_10;
  assign widget__EVAL_26 = buffer_1__EVAL_9;
  assign _EVAL_9 = buffer_1__EVAL_11;
  assign buffer_1__EVAL_17 = _EVAL_34;
  assign widget__EVAL_2 = buffer_1__EVAL_16;
  assign buffer_1__EVAL_27 = widget__EVAL_44;
  assign _EVAL_8 = tl2ahb__EVAL_12;
  assign widget__EVAL_4 = buffer_1__EVAL_22;
  assign widget__EVAL_29 = buffer_1__EVAL_6;
  assign widget__EVAL_13 = buffer__EVAL_11;
  assign buffer__EVAL_35 = widget__EVAL_43;
  assign buffer__EVAL_24 = widget__EVAL_27;
  assign buffer_1__EVAL_44 = _EVAL_11;
  assign widget__EVAL_22 = _EVAL_12;
  assign tl2ahb__EVAL_9 = buffer__EVAL_33;
  assign buffer_1__EVAL_42 = widget__EVAL_42;
  assign tl2ahb__EVAL_16 = buffer__EVAL_1;
  assign _EVAL_21 = tl2ahb__EVAL_11;
  assign buffer__EVAL_15 = tl2ahb__EVAL_32;
  assign buffer_1__EVAL_2 = _EVAL_4;
  assign buffer_1__EVAL_8 = _EVAL_1;
  assign tl2ahb__EVAL_20 = buffer__EVAL_18;
  assign buffer__EVAL_17 = _EVAL_11;
  assign buffer_1__EVAL_26 = widget__EVAL_41;
  assign widget__EVAL_28 = buffer__EVAL_45;
  assign buffer__EVAL_34 = widget__EVAL_33;
  assign _EVAL_14 = buffer_1__EVAL_14;
  assign tl2ahb__EVAL_13 = buffer__EVAL_10;
  assign buffer__EVAL_9 = tl2ahb__EVAL_7;
  assign buffer__EVAL_13 = widget__EVAL_38;
  assign buffer__EVAL_21 = widget__EVAL_0;
  assign buffer_1__EVAL_23 = widget__EVAL_45;
  assign buffer_1__EVAL_32 = widget__EVAL_23;
  assign _EVAL_0 = buffer_1__EVAL_7;
  assign buffer__EVAL_6 = tl2ahb__EVAL_10;
  assign widget__EVAL_19 = buffer__EVAL_0;
  assign buffer_1__EVAL = _EVAL_31;
  assign widget__EVAL_40 = buffer_1__EVAL_46;
  assign widget__EVAL_6 = buffer__EVAL_30;
  assign widget__EVAL_37 = buffer_1__EVAL_4;
  assign _EVAL_26 = tl2ahb__EVAL_25;
  assign tl2ahb__EVAL_33 = _EVAL_30;
  assign buffer_1__EVAL_20 = _EVAL_13;
  assign tl2ahb__EVAL_2 = buffer__EVAL_37;
  assign _EVAL_29 = buffer_1__EVAL_0;
  assign tl2ahb__EVAL_34 = buffer__EVAL_32;
  assign buffer__EVAL_47 = widget__EVAL_34;
  assign buffer__EVAL_29 = tl2ahb__EVAL_4;
  assign buffer__EVAL_40 = widget__EVAL_20;
  assign buffer_1__EVAL_47 = _EVAL_22;
  assign widget__EVAL_8 = buffer_1__EVAL_28;
  assign widget__EVAL_46 = buffer_1__EVAL_36;
  assign _EVAL_7 = tl2ahb__EVAL_6;
  assign widget__EVAL_11 = buffer__EVAL_28;
  assign buffer_1__EVAL_5 = _EVAL_27;
  assign buffer__EVAL_14 = tl2ahb__EVAL_30;
  assign buffer__EVAL_7 = widget__EVAL_5;
  assign buffer_1__EVAL_38 = widget__EVAL_17;
  assign tl2ahb__EVAL_19 = buffer__EVAL_27;
  assign widget__EVAL_3 = buffer_1__EVAL_13;
  assign widget__EVAL_32 = _EVAL_11;
  assign widget__EVAL_16 = buffer_1__EVAL_3;
  assign buffer_1__EVAL_24 = widget__EVAL_7;
  assign buffer__EVAL = tl2ahb__EVAL_21;
  assign buffer_1__EVAL_31 = _EVAL_15;
  assign buffer_1__EVAL_45 = _EVAL_5;
  assign _EVAL_20 = tl2ahb__EVAL_5;
  assign buffer__EVAL_4 = widget__EVAL_47;
  assign tl2ahb__EVAL_3 = _EVAL_28;
  assign tl2ahb__EVAL_28 = buffer__EVAL_3;
  assign _EVAL_10 = buffer_1__EVAL_30;
  assign widget__EVAL_15 = buffer__EVAL_38;
  assign buffer__EVAL_44 = tl2ahb__EVAL_23;
  assign tl2ahb__EVAL_22 = buffer__EVAL_23;
  assign _EVAL_18 = buffer_1__EVAL_1;
  assign buffer_1__EVAL_29 = _EVAL_16;
  assign widget__EVAL_1 = buffer__EVAL_39;
  assign tl2ahb__EVAL_31 = buffer__EVAL_31;
  assign tl2ahb__EVAL_26 = buffer__EVAL_43;
  assign buffer__EVAL_25 = widget__EVAL_36;
  assign buffer__EVAL_5 = widget__EVAL_25;
  assign widget__EVAL_39 = buffer__EVAL_16;
  assign buffer__EVAL_42 = tl2ahb__EVAL_8;
  assign buffer_1__EVAL_37 = _EVAL_12;
  assign buffer__EVAL_8 = widget__EVAL_48;
  assign _EVAL_2 = tl2ahb__EVAL_27;
  assign _EVAL_24 = buffer_1__EVAL_41;
  assign buffer_1__EVAL_21 = _EVAL_17;
  assign _EVAL_33 = buffer_1__EVAL_33;
  assign buffer__EVAL_48 = tl2ahb__EVAL_15;
  assign widget__EVAL_31 = buffer_1__EVAL_19;
  assign _EVAL_25 = buffer_1__EVAL_35;
  assign _EVAL_19 = tl2ahb__EVAL_18;
  assign widget__EVAL_14 = buffer__EVAL_12;
  assign buffer_1__EVAL_18 = _EVAL_6;
  assign buffer_1__EVAL_12 = _EVAL_32;
  assign buffer__EVAL_20 = widget__EVAL_30;
  assign buffer__EVAL_46 = tl2ahb__EVAL_0;
  assign buffer_1__EVAL_15 = widget__EVAL_24;
  assign tl2ahb__EVAL = _EVAL_23;
  assign buffer_1__EVAL_39 = widget__EVAL;
  assign widget__EVAL_12 = buffer_1__EVAL_34;
  assign widget__EVAL_10 = buffer__EVAL_22;
  assign tl2ahb__EVAL_1 = buffer__EVAL_19;
  assign tl2ahb__EVAL_29 = _EVAL_11;
  assign buffer__EVAL_26 = widget__EVAL_21;
  assign buffer_1__EVAL_40 = widget__EVAL_35;
  assign buffer__EVAL_36 = _EVAL_12;
  assign widget__EVAL_18 = buffer_1__EVAL_43;
  assign widget__EVAL_9 = buffer_1__EVAL_48;
  assign tl2ahb__EVAL_17 = _EVAL_12;
  assign tl2ahb__EVAL_14 = buffer__EVAL_2;
  assign buffer_1__EVAL_25 = _EVAL;
  assign tl2ahb__EVAL_24 = buffer__EVAL_41;
endmodule
