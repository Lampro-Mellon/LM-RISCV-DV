//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_24(
  input  [2:0]  _EVAL,
  output [31:0] _EVAL_0,
  output        _EVAL_1,
  output [2:0]  _EVAL_2,
  output        _EVAL_3,
  input  [3:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  input  [1:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  output        _EVAL_10,
  output        _EVAL_11,
  output        _EVAL_12,
  input         _EVAL_13,
  input  [2:0]  _EVAL_14,
  input  [2:0]  _EVAL_15,
  output [2:0]  _EVAL_16,
  input         _EVAL_17,
  output [2:0]  _EVAL_18,
  output [2:0]  _EVAL_19,
  input  [2:0]  _EVAL_20,
  input         _EVAL_21,
  output [2:0]  _EVAL_22,
  output        _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  input  [2:0]  _EVAL_26,
  output        _EVAL_27,
  output [1:0]  _EVAL_28,
  input         _EVAL_29,
  output        _EVAL_30,
  output [2:0]  _EVAL_31,
  output        _EVAL_32,
  output [3:0]  _EVAL_33,
  input  [30:0] _EVAL_34,
  input  [31:0] _EVAL_35,
  input         _EVAL_36,
  output [30:0] _EVAL_37,
  output        _EVAL_38,
  output [2:0]  _EVAL_39,
  input  [2:0]  _EVAL_40,
  output        _EVAL_41,
  input         _EVAL_42,
  output [31:0] _EVAL_43,
  input         _EVAL_44,
  output        _EVAL_45,
  input  [31:0] _EVAL_46,
  input         _EVAL_47,
  input         _EVAL_48
);
  assign _EVAL_3 = _EVAL_13;
  assign _EVAL_31 = _EVAL_20;
  assign _EVAL_10 = _EVAL_25;
  assign _EVAL_12 = _EVAL_44;
  assign _EVAL_16 = _EVAL_14;
  assign _EVAL_27 = _EVAL_7;
  assign _EVAL_22 = _EVAL;
  assign _EVAL_23 = _EVAL_21;
  assign _EVAL_30 = _EVAL_9;
  assign _EVAL_0 = _EVAL_46;
  assign _EVAL_2 = _EVAL_26;
  assign _EVAL_18 = _EVAL_40;
  assign _EVAL_43 = _EVAL_35;
  assign _EVAL_33 = _EVAL_4;
  assign _EVAL_32 = _EVAL_47;
  assign _EVAL_45 = _EVAL_29;
  assign _EVAL_28 = _EVAL_6;
  assign _EVAL_19 = _EVAL_5;
  assign _EVAL_1 = _EVAL_24;
  assign _EVAL_11 = _EVAL_42;
  assign _EVAL_41 = _EVAL_8;
  assign _EVAL_38 = _EVAL_48;
  assign _EVAL_37 = _EVAL_34;
  assign _EVAL_39 = _EVAL_15;
endmodule
