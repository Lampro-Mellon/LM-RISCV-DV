//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_181(
  output [31:0] _EVAL,
  output [1:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  output        _EVAL_4,
  output        _EVAL_5,
  output        _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [31:0] _EVAL_9,
  output [6:0]  _EVAL_10,
  input         _EVAL_11,
  input  [1:0]  _EVAL_12,
  input  [6:0]  _EVAL_13
);
  reg  _EVAL_15;
  reg [31:0] _RAND_0;
  wire  _EVAL_16;
  wire  _EVAL_18;
  reg  _EVAL_19;
  reg [31:0] _RAND_1;
  reg  _EVAL_21;
  reg [31:0] _RAND_2;
  wire  _EVAL_23;
  reg  _EVAL_24;
  reg [31:0] _RAND_3;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  reg  _EVAL_33;
  reg [31:0] _RAND_4;
  wire [9:0] _EVAL_35;
  wire  _EVAL_39;
  reg  _EVAL_44;
  reg [31:0] _RAND_5;
  reg  _EVAL_46;
  reg [31:0] _RAND_6;
  reg  _EVAL_47;
  reg [31:0] _RAND_7;
  wire  _EVAL_48;
  reg  _EVAL_50;
  reg [31:0] _RAND_8;
  reg  _EVAL_52;
  reg [31:0] _RAND_9;
  wire  _EVAL_55;
  reg  _EVAL_56;
  reg [31:0] _RAND_10;
  reg  _EVAL_59;
  reg [31:0] _RAND_11;
  reg  _EVAL_61;
  reg [31:0] _RAND_12;
  reg  _EVAL_62;
  reg [31:0] _RAND_13;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire [4:0] _EVAL_67;
  wire [9:0] _EVAL_68;
  reg  _EVAL_75;
  reg [31:0] _RAND_14;
  wire  _EVAL_76;
  wire  _EVAL_79;
  wire [40:0] _EVAL_81;
  wire  _EVAL_84;
  reg  _EVAL_87;
  reg [31:0] _RAND_15;
  wire  _EVAL_91;
  reg  _EVAL_93;
  reg [31:0] _RAND_16;
  reg  _EVAL_95;
  reg [31:0] _RAND_17;
  wire  _EVAL_98;
  reg  _EVAL_100;
  reg [31:0] _RAND_18;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_112;
  wire  _EVAL_114;
  reg  _EVAL_115;
  reg [31:0] _RAND_19;
  wire [9:0] _EVAL_116;
  reg  _EVAL_117;
  reg [31:0] _RAND_20;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  reg  _EVAL_122;
  reg [31:0] _RAND_21;
  wire  _EVAL_124;
  reg  _EVAL_125;
  reg [31:0] _RAND_22;
  wire  _EVAL_126;
  reg  _EVAL_128;
  reg [31:0] _RAND_23;
  reg  _EVAL_131;
  reg [31:0] _RAND_24;
  wire  _EVAL_134;
  wire  _EVAL_135;
  reg  _EVAL_137;
  reg [31:0] _RAND_25;
  wire  _EVAL_138;
  wire [40:0] _EVAL_139;
  reg  _EVAL_140;
  reg [31:0] _RAND_26;
  reg  _EVAL_141;
  reg [31:0] _RAND_27;
  reg  _EVAL_142;
  reg [31:0] _RAND_28;
  wire  _EVAL_144;
  wire  _EVAL_146;
  wire  _EVAL_148;
  reg  _EVAL_149;
  reg [31:0] _RAND_29;
  reg  _EVAL_151;
  reg [31:0] _RAND_30;
  reg  _EVAL_153;
  reg [31:0] _RAND_31;
  wire  _EVAL_156;
  wire  _EVAL_157;
  reg  _EVAL_158;
  reg [31:0] _RAND_32;
  reg  _EVAL_159;
  reg [31:0] _RAND_33;
  wire  _EVAL_161;
  reg  _EVAL_163;
  reg [31:0] _RAND_34;
  wire  _EVAL_175;
  reg  _EVAL_179;
  reg [31:0] _RAND_35;
  reg  _EVAL_180;
  reg [31:0] _RAND_36;
  reg  _EVAL_181;
  reg [31:0] _RAND_37;
  reg  _EVAL_183;
  reg [31:0] _RAND_38;
  wire  _EVAL_184;
  reg  _EVAL_189;
  reg [31:0] _RAND_39;
  wire  _EVAL_190;
  reg  _EVAL_191;
  reg [31:0] _RAND_40;
  wire  _EVAL_195;
  assign _EVAL_84 = _EVAL_139[40];
  assign _EVAL_35 = {_EVAL_75,_EVAL_180,_EVAL_158,_EVAL_131,_EVAL_15,_EVAL_159,_EVAL_149,_EVAL_137,_EVAL_50,_EVAL_115};
  assign _EVAL_39 = _EVAL_139[21];
  assign _EVAL_161 = _EVAL_139[20];
  assign _EVAL_76 = _EVAL_139[17];
  assign _EVAL_135 = _EVAL_139[24];
  assign _EVAL_81 = {_EVAL_56,_EVAL_93,_EVAL_95,_EVAL_189,_EVAL_183,_EVAL_141,_EVAL_67,_EVAL_35,_EVAL_68,_EVAL_116};
  assign _EVAL_64 = _EVAL_139[5];
  assign _EVAL_48 = _EVAL_139[6];
  assign _EVAL_138 = _EVAL_139[8];
  assign _EVAL_91 = _EVAL_139[36];
  assign _EVAL_32 = _EVAL_139[2];
  assign _EVAL_148 = _EVAL_139[10];
  assign _EVAL_79 = _EVAL_139[9];
  assign _EVAL_68 = {_EVAL_33,_EVAL_163,_EVAL_59,_EVAL_100,_EVAL_44,_EVAL_24,_EVAL_46,_EVAL_47,_EVAL_87,_EVAL_191};
  assign _EVAL_114 = _EVAL_139[27];
  assign _EVAL_184 = _EVAL_139[34];
  assign _EVAL_121 = _EVAL_139[28];
  assign _EVAL_175 = _EVAL_139[11];
  assign _EVAL_126 = _EVAL_139[14];
  assign _EVAL_23 = _EVAL_139[39];
  assign _EVAL = _EVAL_81[33:2];
  assign _EVAL_10 = _EVAL_81[40:34];
  assign _EVAL_67 = {_EVAL_19,_EVAL_117,_EVAL_62,_EVAL_21,_EVAL_151};
  assign _EVAL_26 = _EVAL_139[15];
  assign _EVAL_157 = _EVAL_139[29];
  assign _EVAL_190 = _EVAL_139[25];
  assign _EVAL_16 = _EVAL_139[3];
  assign _EVAL_4 = _EVAL_11;
  assign _EVAL_55 = _EVAL_139[32];
  assign _EVAL_27 = _EVAL_139[19];
  assign _EVAL_31 = _EVAL_139[4];
  assign _EVAL_18 = _EVAL_139[16];
  assign _EVAL_195 = _EVAL_139[30];
  assign _EVAL_144 = _EVAL_139[37];
  assign _EVAL_120 = _EVAL_139[31];
  assign _EVAL_98 = _EVAL_139[23];
  assign _EVAL_6 = _EVAL_11 ? 1'h0 : _EVAL_2;
  assign _EVAL_124 = _EVAL_139[13];
  assign _EVAL_30 = _EVAL_139[22];
  assign _EVAL_156 = _EVAL_139[35];
  assign _EVAL_116 = {_EVAL_122,_EVAL_179,_EVAL_61,_EVAL_142,_EVAL_181,_EVAL_140,_EVAL_153,_EVAL_125,_EVAL_52,_EVAL_128};
  assign _EVAL_139 = {_EVAL_13,_EVAL_9,_EVAL_12};
  assign _EVAL_110 = _EVAL_139[0];
  assign _EVAL_109 = _EVAL_139[1];
  assign _EVAL_28 = _EVAL_139[18];
  assign _EVAL_134 = _EVAL_139[38];
  assign _EVAL_5 = _EVAL_128;
  assign _EVAL_112 = _EVAL_139[33];
  assign _EVAL_119 = _EVAL_139[26];
  assign _EVAL_0 = _EVAL_81[1:0];
  assign _EVAL_65 = _EVAL_139[12];
  assign _EVAL_146 = _EVAL_139[7];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_19 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_21 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_24 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_33 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_44 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_46 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_47 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_50 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_52 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_56 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_59 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_61 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_62 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_75 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_87 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_93 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_95 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_100 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_115 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_117 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_122 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_125 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_128 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_131 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_137 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_140 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_141 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_142 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_149 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_151 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_153 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_158 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_159 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_163 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_179 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_180 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_181 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _EVAL_183 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _EVAL_189 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _EVAL_191 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_3) begin
    if (_EVAL_11) begin
      _EVAL_15 <= _EVAL_190;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_15 <= _EVAL_131;
      end
    end
    if (_EVAL_11) begin
      _EVAL_19 <= _EVAL_184;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_19 <= _EVAL_141;
      end
    end
    if (_EVAL_11) begin
      _EVAL_21 <= _EVAL_120;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_21 <= _EVAL_62;
      end
    end
    if (_EVAL_11) begin
      _EVAL_24 <= _EVAL_126;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_24 <= _EVAL_44;
      end
    end
    if (_EVAL_11) begin
      _EVAL_33 <= _EVAL_27;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_33 <= _EVAL_115;
      end
    end
    if (_EVAL_11) begin
      _EVAL_44 <= _EVAL_26;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_44 <= _EVAL_100;
      end
    end
    if (_EVAL_11) begin
      _EVAL_46 <= _EVAL_124;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_46 <= _EVAL_24;
      end
    end
    if (_EVAL_11) begin
      _EVAL_47 <= _EVAL_65;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_47 <= _EVAL_46;
      end
    end
    if (_EVAL_11) begin
      _EVAL_50 <= _EVAL_39;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_50 <= _EVAL_137;
      end
    end
    if (_EVAL_11) begin
      _EVAL_52 <= _EVAL_109;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_52 <= _EVAL_125;
      end
    end
    if (_EVAL_11) begin
      _EVAL_56 <= _EVAL_84;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_56 <= _EVAL_8;
      end
    end
    if (_EVAL_11) begin
      _EVAL_59 <= _EVAL_76;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_59 <= _EVAL_163;
      end
    end
    if (_EVAL_11) begin
      _EVAL_61 <= _EVAL_146;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_61 <= _EVAL_179;
      end
    end
    if (_EVAL_11) begin
      _EVAL_62 <= _EVAL_55;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_62 <= _EVAL_117;
      end
    end
    if (_EVAL_11) begin
      _EVAL_75 <= _EVAL_157;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_75 <= _EVAL_151;
      end
    end
    if (_EVAL_11) begin
      _EVAL_87 <= _EVAL_175;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_87 <= _EVAL_47;
      end
    end
    if (_EVAL_11) begin
      _EVAL_93 <= _EVAL_23;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_93 <= _EVAL_56;
      end
    end
    if (_EVAL_11) begin
      _EVAL_95 <= _EVAL_134;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_95 <= _EVAL_93;
      end
    end
    if (_EVAL_11) begin
      _EVAL_100 <= _EVAL_18;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_100 <= _EVAL_59;
      end
    end
    if (_EVAL_11) begin
      _EVAL_115 <= _EVAL_161;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_115 <= _EVAL_50;
      end
    end
    if (_EVAL_11) begin
      _EVAL_117 <= _EVAL_112;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_117 <= _EVAL_19;
      end
    end
    if (_EVAL_11) begin
      _EVAL_122 <= _EVAL_79;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_122 <= _EVAL_191;
      end
    end
    if (_EVAL_11) begin
      _EVAL_125 <= _EVAL_32;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_125 <= _EVAL_153;
      end
    end
    if (_EVAL_11) begin
      _EVAL_128 <= _EVAL_110;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_128 <= _EVAL_52;
      end
    end
    if (_EVAL_11) begin
      _EVAL_131 <= _EVAL_119;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_131 <= _EVAL_158;
      end
    end
    if (_EVAL_11) begin
      _EVAL_137 <= _EVAL_30;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_137 <= _EVAL_149;
      end
    end
    if (_EVAL_11) begin
      _EVAL_140 <= _EVAL_31;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_140 <= _EVAL_181;
      end
    end
    if (_EVAL_11) begin
      _EVAL_141 <= _EVAL_156;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_141 <= _EVAL_183;
      end
    end
    if (_EVAL_11) begin
      _EVAL_142 <= _EVAL_48;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_142 <= _EVAL_61;
      end
    end
    if (_EVAL_11) begin
      _EVAL_149 <= _EVAL_98;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_149 <= _EVAL_159;
      end
    end
    if (_EVAL_11) begin
      _EVAL_151 <= _EVAL_195;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_151 <= _EVAL_21;
      end
    end
    if (_EVAL_11) begin
      _EVAL_153 <= _EVAL_16;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_153 <= _EVAL_140;
      end
    end
    if (_EVAL_11) begin
      _EVAL_158 <= _EVAL_114;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_158 <= _EVAL_180;
      end
    end
    if (_EVAL_11) begin
      _EVAL_159 <= _EVAL_135;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_159 <= _EVAL_15;
      end
    end
    if (_EVAL_11) begin
      _EVAL_163 <= _EVAL_28;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_163 <= _EVAL_33;
      end
    end
    if (_EVAL_11) begin
      _EVAL_179 <= _EVAL_138;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_179 <= _EVAL_122;
      end
    end
    if (_EVAL_11) begin
      _EVAL_180 <= _EVAL_121;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_180 <= _EVAL_75;
      end
    end
    if (_EVAL_11) begin
      _EVAL_181 <= _EVAL_64;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_181 <= _EVAL_142;
      end
    end
    if (_EVAL_11) begin
      _EVAL_183 <= _EVAL_91;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_183 <= _EVAL_189;
      end
    end
    if (_EVAL_11) begin
      _EVAL_189 <= _EVAL_144;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_189 <= _EVAL_95;
      end
    end
    if (_EVAL_11) begin
      _EVAL_191 <= _EVAL_148;
    end else if (!(_EVAL_2)) begin
      if (_EVAL_7) begin
        _EVAL_191 <= _EVAL_87;
      end
    end
  end
endmodule
