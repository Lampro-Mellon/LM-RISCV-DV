//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_4(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  output [2:0]  _EVAL_2,
  output [29:0] _EVAL_3,
  output        _EVAL_4,
  output        _EVAL_5,
  input  [3:0]  _EVAL_6,
  input  [3:0]  _EVAL_7,
  input  [1:0]  _EVAL_8,
  output        _EVAL_9,
  output [2:0]  _EVAL_10,
  output [3:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input  [2:0]  _EVAL_15,
  output [31:0] _EVAL_16,
  output [1:0]  _EVAL_17,
  output        _EVAL_18,
  output [1:0]  _EVAL_19,
  input         _EVAL_20,
  output        _EVAL_21,
  input  [2:0]  _EVAL_22,
  input         _EVAL_23,
  output        _EVAL_24,
  input  [2:0]  _EVAL_25,
  output        _EVAL_26,
  output [2:0]  _EVAL_27,
  input         _EVAL_28,
  output [1:0]  _EVAL_29,
  input  [2:0]  _EVAL_30,
  output        _EVAL_31,
  output        _EVAL_32,
  input         _EVAL_33,
  input  [2:0]  _EVAL_34,
  output [2:0]  _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  output [1:0]  _EVAL_38,
  output [31:0] _EVAL_39,
  input         _EVAL_40,
  output [3:0]  _EVAL_41,
  output        _EVAL_42,
  output [2:0]  _EVAL_43,
  output        _EVAL_44,
  input         _EVAL_45,
  input         _EVAL_46,
  input         _EVAL_47,
  input         _EVAL_48,
  output        _EVAL_49,
  input  [31:0] _EVAL_50,
  output [2:0]  _EVAL_51,
  input  [3:0]  _EVAL_52,
  output [2:0]  _EVAL_53,
  output        _EVAL_54,
  input         _EVAL_55,
  output        _EVAL_56,
  output [31:0] _EVAL_57,
  input  [31:0] _EVAL_58,
  input  [1:0]  _EVAL_59,
  output [31:0] _EVAL_60,
  input  [3:0]  _EVAL_61,
  output        _EVAL_62,
  output        _EVAL_63,
  output        _EVAL_64,
  output [3:0]  _EVAL_65,
  output        _EVAL_66,
  output        _EVAL_67,
  output [30:0] _EVAL_68,
  input         _EVAL_69,
  output [2:0]  _EVAL_70,
  input         _EVAL_71,
  input  [31:0] _EVAL_72,
  input         _EVAL_73,
  input         _EVAL_74,
  input         _EVAL_75,
  output        _EVAL_76,
  output [31:0] _EVAL_77,
  output [2:0]  _EVAL_78,
  input  [2:0]  _EVAL_79,
  output        _EVAL_80,
  output        _EVAL_81,
  output [1:0]  _EVAL_82,
  input  [31:0] _EVAL_83,
  output        _EVAL_84,
  input  [31:0] _EVAL_85,
  input  [2:0]  _EVAL_86,
  input  [2:0]  _EVAL_87,
  output        _EVAL_88,
  input  [2:0]  _EVAL_89,
  input         _EVAL_90,
  input         _EVAL_91,
  output [3:0]  _EVAL_92,
  input  [2:0]  _EVAL_93,
  input         _EVAL_94,
  input  [1:0]  _EVAL_95,
  input         _EVAL_96,
  input         _EVAL_97,
  output        _EVAL_98,
  output [31:0] _EVAL_99,
  output [31:0] _EVAL_100,
  input  [2:0]  _EVAL_101,
  output [31:0] _EVAL_102,
  output        _EVAL_103,
  input         _EVAL_104,
  output [3:0]  _EVAL_105,
  output [2:0]  _EVAL_106,
  output        _EVAL_107,
  input         _EVAL_108,
  input         _EVAL_109,
  input  [31:0] _EVAL_110,
  input         _EVAL_111,
  input  [2:0]  _EVAL_112,
  input         _EVAL_113,
  output [2:0]  _EVAL_114,
  input  [3:0]  _EVAL_115,
  output        _EVAL_116,
  input  [31:0] _EVAL_117,
  output [2:0]  _EVAL_118,
  input         _EVAL_119,
  input  [3:0]  _EVAL_120,
  input  [2:0]  _EVAL_121,
  input         _EVAL_122,
  output [31:0] _EVAL_123,
  input         _EVAL_124,
  input         _EVAL_125,
  output        _EVAL_126,
  output        _EVAL_127,
  input  [2:0]  _EVAL_128,
  output [2:0]  _EVAL_129,
  output [3:0]  _EVAL_130,
  output [3:0]  _EVAL_131,
  input  [31:0] _EVAL_132,
  input         _EVAL_133,
  input  [31:0] _EVAL_134,
  input  [2:0]  _EVAL_135,
  input  [31:0] _EVAL_136,
  output [2:0]  _EVAL_137,
  input         _EVAL_138,
  input         _EVAL_139,
  output [2:0]  _EVAL_140,
  input  [3:0]  _EVAL_141,
  output [3:0]  _EVAL_142,
  input  [1:0]  _EVAL_143,
  output        _EVAL_144,
  output        _EVAL_145,
  output        _EVAL_146,
  output        _EVAL_147,
  input         _EVAL_148,
  input         _EVAL_149,
  input         _EVAL_150,
  output        _EVAL_151,
  input         _EVAL_152,
  output [2:0]  _EVAL_153,
  input         _EVAL_154,
  input         _EVAL_155,
  output        _EVAL_156,
  output        _EVAL_157,
  output        _EVAL_158,
  output        _EVAL_159,
  input         _EVAL_160,
  output        _EVAL_161,
  input         _EVAL_162,
  input         _EVAL_163
);
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire [32:0] _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire [22:0] _EVAL_170;
  wire  _EVAL_171;
  wire [88:0] _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire [32:0] _EVAL_180;
  wire [5:0] _EVAL_181;
  wire  _EVAL_183;
  wire [46:0] _EVAL_184;
  wire [32:0] _EVAL_185;
  wire [3:0] _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire [6:0] _EVAL_190;
  reg [2:0] _EVAL_192;
  reg [31:0] _RAND_0;
  wire  _EVAL_193;
  wire  _EVAL_195;
  wire [32:0] _EVAL_196;
  wire  _EVAL_197;
  wire [5:0] _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire [32:0] _EVAL_201;
  wire  _EVAL_202;
  wire [2:0] _EVAL_203;
  wire [3:0] _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire [20:0] _EVAL_208;
  wire [88:0] _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  reg [5:0] _EVAL_213;
  reg [31:0] _RAND_1;
  wire  _EVAL_214;
  wire [2:0] _EVAL_216;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire [5:0] _EVAL_221;
  wire [2:0] _EVAL_222;
  wire [46:0] _EVAL_223;
  wire [32:0] _EVAL_224;
  wire [5:0] _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire [3:0] _EVAL_228;
  wire [5:0] _EVAL_230;
  wire  _EVAL_231;
  wire [2:0] _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire [7:0] _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_239;
  wire [32:0] _EVAL_240;
  wire [4:0] _EVAL_241;
  wire [3:0] _EVAL_242;
  wire [32:0] _EVAL_243;
  wire  _EVAL_244;
  wire [2:0] _EVAL_245;
  wire [5:0] _EVAL_246;
  wire [31:0] _EVAL_247;
  wire [2:0] _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire [5:0] _EVAL_251;
  wire  _EVAL_252;
  wire [88:0] _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire [3:0] _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire [32:0] _EVAL_260;
  wire  _EVAL_261;
  wire [31:0] _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire [2:0] _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_273;
  wire [2:0] _EVAL_274;
  reg  _EVAL_275;
  reg [31:0] _RAND_2;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire [5:0] _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire [6:0] _EVAL_281;
  wire [3:0] _EVAL_282;
  wire  _EVAL_283;
  wire [3:0] _EVAL_284;
  wire  _EVAL_285;
  wire [2:0] _EVAL_286;
  wire [32:0] _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire [7:0] _EVAL_296;
  wire [4:0] _EVAL_297;
  wire [4:0] _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_303;
  wire [2:0] _EVAL_306;
  wire  _EVAL_307;
  wire [3:0] _EVAL_309;
  wire  _EVAL_310;
  wire [32:0] _EVAL_311;
  wire [5:0] _EVAL_312;
  wire  _EVAL_313;
  wire [3:0] _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_318;
  wire [46:0] _EVAL_319;
  wire [5:0] _EVAL_320;
  wire [88:0] _EVAL_321;
  wire  _EVAL_322;
  wire [32:0] _EVAL_323;
  wire  _EVAL_324;
  wire  _EVAL_325;
  wire [3:0] _EVAL_327;
  wire [5:0] _EVAL_328;
  wire  _EVAL_329;
  wire [6:0] _EVAL_330;
  wire  _EVAL_331;
  wire  _EVAL_332;
  reg  _EVAL_334;
  reg [31:0] _RAND_3;
  wire  _EVAL_338;
  wire [5:0] _EVAL_340;
  wire [46:0] _EVAL_341;
  reg  _EVAL_342;
  reg [31:0] _RAND_4;
  wire [32:0] _EVAL_343;
  wire  _EVAL_344;
  wire [3:0] _EVAL_345;
  wire [2:0] _EVAL_346;
  wire [46:0] _EVAL_347;
  wire  _EVAL_348;
  wire [1:0] _EVAL_349;
  reg [5:0] _EVAL_351;
  reg [31:0] _RAND_5;
  wire [88:0] _EVAL_353;
  wire  _EVAL_354;
  wire  _EVAL_355;
  wire [32:0] _EVAL_356;
  wire [5:0] _EVAL_357;
  wire  _EVAL_358;
  wire  _EVAL_359;
  reg [3:0] _EVAL_361;
  reg [31:0] _RAND_6;
  wire [2:0] _EVAL_362;
  wire  _EVAL_363;
  wire [40:0] _EVAL_364;
  wire [46:0] _EVAL_366;
  wire [5:0] _EVAL_367;
  wire [46:0] _EVAL_368;
  wire [3:0] _EVAL_369;
  wire [3:0] _EVAL_370;
  wire  _EVAL_371;
  reg  _EVAL_373;
  reg [31:0] _RAND_7;
  wire  _EVAL_374;
  wire [2:0] _EVAL_375;
  reg [3:0] _EVAL_376;
  reg [31:0] _RAND_8;
  wire  _EVAL_377;
  wire  _EVAL_378;
  wire  _EVAL_379;
  wire  _EVAL_380;
  wire [2:0] _EVAL_381;
  wire  _EVAL_382;
  wire  _EVAL_383;
  wire  _EVAL_384;
  wire [2:0] _EVAL_385;
  wire [5:0] _EVAL_386;
  wire [2:0] _EVAL_387;
  wire [88:0] _EVAL_388;
  wire  _EVAL_389;
  wire [5:0] _EVAL_391;
  wire  _EVAL_392;
  wire [2:0] _EVAL_393;
  wire  _EVAL_394;
  wire [32:0] _EVAL_396;
  wire [3:0] _EVAL_397;
  wire  _EVAL_398;
  wire [5:0] _EVAL_399;
  wire [3:0] _EVAL_401;
  wire [22:0] _EVAL_402;
  wire  _EVAL_403;
  wire [3:0] _EVAL_404;
  wire  _EVAL_405;
  wire [3:0] _EVAL_406;
  wire  _EVAL_408;
  wire [5:0] _EVAL_409;
  wire [88:0] _EVAL_410;
  wire  _EVAL_413;
  wire [5:0] _EVAL_414;
  wire [32:0] _EVAL_415;
  wire [32:0] _EVAL_416;
  wire  _EVAL_418;
  wire [32:0] _EVAL_420;
  wire [46:0] _EVAL_421;
  wire [2:0] _EVAL_422;
  wire [3:0] _EVAL_424;
  wire  _EVAL_425;
  wire  _EVAL_427;
  wire  _EVAL_429;
  wire [3:0] _EVAL_430;
  wire  _EVAL_432;
  wire [5:0] _EVAL_433;
  wire  _EVAL_434;
  wire [2:0] _EVAL_435;
  wire [46:0] _EVAL_437;
  wire  _EVAL_438;
  wire [5:0] _EVAL_439;
  wire [2:0] _EVAL_440;
  wire [5:0] _EVAL_441;
  wire [46:0] _EVAL_442;
  wire [1:0] _EVAL_443;
  wire [5:0] _EVAL_447;
  wire  _EVAL_448;
  wire  _EVAL_450;
  wire [7:0] _EVAL_451;
  wire [2:0] _EVAL_452;
  reg  _EVAL_453;
  reg [31:0] _RAND_9;
  reg  _EVAL_454;
  reg [31:0] _RAND_10;
  wire [31:0] _EVAL_456;
  wire [5:0] _EVAL_457;
  wire [2:0] _EVAL_458;
  wire [5:0] _EVAL_459;
  wire  _EVAL_460;
  wire  _EVAL_461;
  wire [88:0] _EVAL_462;
  wire [5:0] _EVAL_463;
  wire  _EVAL_464;
  wire  _EVAL_465;
  wire [46:0] _EVAL_466;
  wire [2:0] _EVAL_467;
  wire [7:0] _EVAL_469;
  wire  _EVAL_470;
  wire [5:0] _EVAL_471;
  wire  _EVAL_472;
  wire  _EVAL_473;
  wire [5:0] _EVAL_474;
  reg  _EVAL_476;
  reg [31:0] _RAND_11;
  wire [4:0] _EVAL_477;
  wire [31:0] _EVAL_478;
  wire  _EVAL_479;
  reg  _EVAL_480;
  reg [31:0] _RAND_12;
  wire  _EVAL_481;
  wire [32:0] _EVAL_482;
  wire [46:0] _EVAL_483;
  wire  _EVAL_485;
  wire  _EVAL_486;
  wire  _EVAL_487;
  wire [32:0] _EVAL_488;
  wire [5:0] _EVAL_489;
  wire [2:0] _EVAL_490;
  wire [7:0] _EVAL_491;
  reg  _EVAL_492;
  reg [31:0] _RAND_13;
  wire  _EVAL_493;
  reg [5:0] _EVAL_494;
  reg [31:0] _RAND_14;
  wire [5:0] _EVAL_495;
  wire  _EVAL_496;
  wire  _EVAL_497;
  wire [88:0] _EVAL_498;
  wire [3:0] _EVAL_499;
  wire [32:0] _EVAL_500;
  reg [2:0] _EVAL_501;
  reg [31:0] _RAND_15;
  wire  _EVAL_502;
  wire [3:0] _EVAL_503;
  wire [32:0] _EVAL_504;
  wire  _EVAL_506;
  wire [6:0] _EVAL_507;
  wire  _EVAL_509;
  wire  _EVAL_510;
  wire  _EVAL_511;
  wire  _EVAL_512;
  wire [2:0] _EVAL_513;
  wire  _EVAL_514;
  wire  _EVAL_515;
  wire [88:0] _EVAL_516;
  wire  _EVAL_517;
  reg  _EVAL_518;
  reg [31:0] _RAND_16;
  wire [3:0] _EVAL_519;
  wire  _EVAL_520;
  wire [32:0] _EVAL_522;
  wire [5:0] _EVAL_523;
  wire [2:0] _EVAL_524;
  wire  _EVAL_525;
  wire  _EVAL_526;
  wire [2:0] _EVAL_527;
  wire [3:0] _EVAL_528;
  wire [2:0] _EVAL_529;
  wire [3:0] _EVAL_530;
  wire [5:0] _EVAL_531;
  wire  _EVAL_532;
  wire  _EVAL_534;
  wire [32:0] _EVAL_536;
  wire [7:0] _EVAL_537;
  wire [5:0] _EVAL_538;
  wire [2:0] _EVAL_539;
  wire  _EVAL_540;
  wire  _EVAL_541;
  wire [2:0] _EVAL_542;
  wire  _EVAL_543;
  wire  _EVAL_544;
  wire  _EVAL_545;
  wire  _EVAL_546;
  wire  _EVAL_548;
  wire [4:0] _EVAL_550;
  wire [46:0] _EVAL_551;
  wire  _EVAL_552;
  wire  _EVAL_553;
  wire [88:0] _EVAL_554;
  reg  _EVAL_555;
  reg [31:0] _RAND_17;
  wire [3:0] _EVAL_557;
  wire  _EVAL_558;
  wire  _EVAL_559;
  wire [3:0] _EVAL_560;
  wire [4:0] _EVAL_562;
  reg  _EVAL_563;
  reg [31:0] _RAND_18;
  wire  _EVAL_564;
  wire  _EVAL_565;
  wire  _EVAL_566;
  wire [3:0] _EVAL_567;
  wire  _EVAL_568;
  wire [32:0] _EVAL_569;
  wire  _EVAL_570;
  wire  _EVAL_571;
  wire [88:0] _EVAL_572;
  wire  _EVAL_573;
  wire [3:0] _EVAL_574;
  wire [1:0] _EVAL_575;
  wire  _EVAL_577;
  wire [5:0] _EVAL_578;
  wire  _EVAL_579;
  wire [7:0] _EVAL_580;
  wire [5:0] _EVAL_583;
  wire [32:0] _EVAL_584;
  wire [7:0] _EVAL_585;
  wire [3:0] _EVAL_586;
  wire [5:0] _EVAL_587;
  wire [4:0] _EVAL_590;
  wire [2:0] _EVAL_592;
  wire  _EVAL_593;
  wire [6:0] _EVAL_594;
  wire [4:0] _EVAL_595;
  wire [5:0] _EVAL_596;
  wire  _EVAL_597;
  wire [5:0] _EVAL_598;
  wire [5:0] _EVAL_599;
  reg  _EVAL_600;
  reg [31:0] _RAND_19;
  wire [31:0] _EVAL_601;
  wire  _EVAL_602;
  wire [40:0] _EVAL_603;
  wire  _EVAL_605;
  wire [46:0] _EVAL_606;
  wire  _EVAL_607;
  wire [7:0] _EVAL_608;
  wire [5:0] _EVAL_609;
  reg  _EVAL_610;
  reg [31:0] _RAND_20;
  reg [3:0] _EVAL_611;
  reg [31:0] _RAND_21;
  wire  _EVAL_612;
  wire [5:0] _EVAL_613;
  wire [5:0] _EVAL_614;
  wire  _EVAL_615;
  wire [5:0] _EVAL_616;
  wire  _EVAL_617;
  wire [3:0] _EVAL_618;
  wire [7:0] _EVAL_619;
  wire [88:0] _EVAL_620;
  wire [6:0] _EVAL_621;
  wire [3:0] _EVAL_622;
  wire [88:0] _EVAL_623;
  wire  _EVAL_624;
  wire [2:0] _EVAL_625;
  wire [88:0] _EVAL_626;
  wire [7:0] _EVAL_627;
  wire [5:0] _EVAL_628;
  wire  _EVAL_629;
  wire [5:0] _EVAL_630;
  wire  _EVAL_631;
  wire  _EVAL_632;
  wire  _EVAL_633;
  wire  _EVAL_634;
  wire [5:0] _EVAL_635;
  wire  _EVAL_636;
  wire [1:0] _EVAL_637;
  wire  _EVAL_638;
  wire [3:0] _EVAL_639;
  wire  _EVAL_640;
  wire [2:0] _EVAL_641;
  reg [5:0] _EVAL_642;
  reg [31:0] _RAND_22;
  wire  _EVAL_643;
  wire [2:0] _EVAL_644;
  wire  _EVAL_645;
  reg  _EVAL_646;
  reg [31:0] _RAND_23;
  wire [2:0] _EVAL_648;
  wire  _EVAL_649;
  wire  _EVAL_651;
  reg [2:0] _EVAL_652;
  reg [31:0] _RAND_24;
  wire  _EVAL_653;
  wire  _EVAL_654;
  wire [88:0] _EVAL_655;
  wire  _EVAL_656;
  wire  _EVAL_657;
  wire  _EVAL_658;
  wire [7:0] _EVAL_659;
  wire [3:0] _EVAL_660;
  wire [3:0] _EVAL_661;
  wire  _EVAL_662;
  wire [5:0] _EVAL_664;
  reg  _EVAL_665;
  reg [31:0] _RAND_25;
  wire  _EVAL_666;
  wire  _EVAL_667;
  wire [3:0] _EVAL_668;
  wire [4:0] _EVAL_669;
  wire [46:0] _EVAL_670;
  wire [5:0] _EVAL_671;
  wire  _EVAL_672;
  wire [3:0] _EVAL_673;
  reg [5:0] _EVAL_674;
  reg [31:0] _RAND_26;
  wire  _EVAL_675;
  wire  _EVAL_676;
  wire [3:0] _EVAL_677;
  wire [5:0] _EVAL_678;
  reg  _EVAL_679;
  reg [31:0] _RAND_27;
  wire [3:0] _EVAL_680;
  wire  _EVAL_681;
  wire [5:0] _EVAL_682;
  wire  _EVAL_683;
  wire [3:0] _EVAL_684;
  wire  _EVAL_685;
  wire [2:0] _EVAL_687;
  wire [5:0] _EVAL_689;
  wire [1:0] _EVAL_690;
  wire [46:0] _EVAL_691;
  wire [3:0] _EVAL_693;
  wire [5:0] _EVAL_694;
  wire [5:0] _EVAL_695;
  wire [2:0] _EVAL_696;
  wire [31:0] _EVAL_698;
  wire [7:0] _EVAL_700;
  wire  _EVAL_701;
  wire [5:0] _EVAL_702;
  wire [7:0] _EVAL_703;
  wire [7:0] _EVAL_704;
  wire  _EVAL_705;
  wire [3:0] _EVAL_706;
  wire [2:0] _EVAL_707;
  wire [5:0] _EVAL_708;
  wire  _EVAL_709;
  wire  _EVAL_710;
  wire [5:0] _EVAL_711;
  wire [88:0] _EVAL_712;
  wire [7:0] _EVAL_714;
  wire [5:0] _EVAL_715;
  wire [22:0] _EVAL_716;
  wire [5:0] _EVAL_717;
  wire  _EVAL_718;
  wire  _EVAL_720;
  wire [2:0] _EVAL_721;
  wire [88:0] _EVAL_722;
  wire  _EVAL_723;
  wire [7:0] _EVAL_724;
  wire [3:0] _EVAL_726;
  wire  _EVAL_727;
  wire [46:0] _EVAL_728;
  wire [7:0] _EVAL_729;
  wire [3:0] _EVAL_730;
  wire [5:0] _EVAL_731;
  wire [6:0] _EVAL_732;
  wire  _EVAL_733;
  wire [6:0] _EVAL_735;
  reg  _EVAL_737;
  reg [31:0] _RAND_28;
  wire [1:0] _EVAL_738;
  wire [3:0] _EVAL_739;
  wire [5:0] _EVAL_740;
  wire [2:0] _EVAL_742;
  wire  _EVAL_743;
  wire [3:0] _EVAL_744;
  wire [5:0] _EVAL_746;
  wire [5:0] _EVAL_747;
  wire  _EVAL_749;
  wire [32:0] _EVAL_750;
  wire [7:0] _EVAL_751;
  wire [46:0] _EVAL_752;
  wire  _EVAL_753;
  wire  _EVAL_754;
  wire  _EVAL_755;
  wire  _EVAL_756;
  wire [2:0] _EVAL_757;
  wire [32:0] _EVAL_758;
  wire [2:0] _EVAL_759;
  wire  _EVAL_760;
  wire  _EVAL_761;
  wire  _EVAL_762;
  wire  _EVAL_763;
  wire [5:0] _EVAL_765;
  wire [46:0] _EVAL_767;
  wire  _EVAL_768;
  wire [5:0] _EVAL_769;
  wire  _EVAL_770;
  reg  _EVAL_771;
  reg [31:0] _RAND_29;
  wire  _EVAL_772;
  wire [5:0] _EVAL_773;
  wire  _EVAL_776;
  wire  _EVAL_777;
  wire [7:0] _EVAL_778;
  wire  _EVAL_779;
  wire [5:0] _EVAL_781;
  wire [3:0] _EVAL_783;
  wire [5:0] _EVAL_784;
  wire [2:0] _EVAL_785;
  wire [3:0] _EVAL_786;
  wire  _EVAL_787;
  wire  _EVAL_788;
  wire [32:0] _EVAL_789;
  wire [22:0] _EVAL_790;
  wire [4:0] _EVAL_791;
  wire  _EVAL_792;
  wire [5:0] _EVAL_793;
  wire  _EVAL_794;
  wire [32:0] _EVAL_796;
  wire  _EVAL_797;
  wire [88:0] _EVAL_798;
  wire  _EVAL_799;
  wire  _EVAL_802;
  wire  _EVAL_803;
  wire [32:0] _EVAL_804;
  wire  _EVAL_806;
  wire  _EVAL_808;
  wire  _EVAL_809;
  wire [2:0] _EVAL_810;
  wire [6:0] _EVAL_811;
  wire [2:0] _EVAL_813;
  wire [3:0] _EVAL_814;
  wire [7:0] _EVAL_817;
  wire [6:0] _EVAL_818;
  wire [3:0] _EVAL_819;
  wire [4:0] _EVAL_820;
  wire [2:0] _EVAL_821;
  wire [3:0] _EVAL_822;
  wire  _EVAL_823;
  wire [5:0] _EVAL_824;
  wire [2:0] _EVAL_825;
  wire [3:0] _EVAL_826;
  wire [32:0] _EVAL_828;
  wire [88:0] _EVAL_829;
  wire  _EVAL_830;
  wire [3:0] _EVAL_832;
  wire  _EVAL_833;
  wire [46:0] _EVAL_834;
  wire [5:0] _EVAL_835;
  wire [46:0] _EVAL_836;
  wire  _EVAL_837;
  reg  _EVAL_838;
  reg [31:0] _RAND_30;
  wire [88:0] _EVAL_839;
  wire  _EVAL_840;
  wire [4:0] _EVAL_841;
  wire  _EVAL_842;
  wire [5:0] _EVAL_843;
  wire [7:0] _EVAL_845;
  wire  _EVAL_846;
  reg  _EVAL_847;
  reg [31:0] _RAND_31;
  wire  _EVAL_848;
  wire [31:0] _EVAL_849;
  wire [32:0] _EVAL_850;
  wire [2:0] _EVAL_851;
  wire [5:0] _EVAL_852;
  wire [32:0] _EVAL_853;
  wire  _EVAL_854;
  wire  _EVAL_855;
  wire  _EVAL_857;
  wire [5:0] _EVAL_859;
  wire  _EVAL_860;
  wire  _EVAL_861;
  wire [5:0] _EVAL_862;
  wire [4:0] _EVAL_863;
  wire  _EVAL_865;
  wire  _EVAL_866;
  wire [88:0] _EVAL_868;
  wire  _EVAL_869;
  wire  _EVAL_870;
  wire  _EVAL_871;
  wire [2:0] _EVAL_872;
  wire [5:0] _EVAL_874;
  wire  _EVAL_876;
  wire [5:0] _EVAL_877;
  wire  _EVAL_878;
  wire  _EVAL_879;
  wire  _EVAL_881;
  wire  _EVAL_882;
  wire  _EVAL_883;
  wire [5:0] _EVAL_884;
  wire  _EVAL_885;
  wire  _EVAL_886;
  wire  _EVAL_887;
  wire  _EVAL_888;
  wire [2:0] _EVAL_889;
  wire  _EVAL_890;
  wire  _EVAL_891;
  wire  _EVAL_892;
  wire  _EVAL_893;
  wire [4:0] _EVAL_894;
  reg [5:0] _EVAL_895;
  reg [31:0] _RAND_32;
  wire  _EVAL_896;
  wire [7:0] _EVAL_898;
  wire [6:0] _EVAL_899;
  wire  _EVAL_900;
  wire [7:0] _EVAL_901;
  wire  _EVAL_903;
  wire  _EVAL_904;
  wire [5:0] _EVAL_905;
  wire [32:0] _EVAL_906;
  wire [7:0] _EVAL_907;
  wire [5:0] _EVAL_908;
  wire [2:0] _EVAL_909;
  wire [5:0] _EVAL_911;
  wire [5:0] _EVAL_912;
  wire [88:0] _EVAL_914;
  wire  _EVAL_915;
  wire [46:0] _EVAL_917;
  wire [7:0] _EVAL_918;
  wire [32:0] _EVAL_919;
  wire  _EVAL_921;
  wire [5:0] _EVAL_922;
  wire  _EVAL_923;
  wire  _EVAL_924;
  wire  _EVAL_925;
  wire  _EVAL_926;
  wire [32:0] _EVAL_927;
  wire  _EVAL_929;
  wire [32:0] _EVAL_931;
  wire [7:0] _EVAL_932;
  wire  _EVAL_934;
  wire  _EVAL_936;
  wire  _EVAL_937;
  wire [5:0] _EVAL_938;
  wire  _EVAL_939;
  wire  _EVAL_940;
  wire [40:0] _EVAL_941;
  wire [32:0] _EVAL_942;
  wire  _EVAL_943;
  wire [2:0] _EVAL_944;
  wire [6:0] _EVAL_945;
  wire [5:0] _EVAL_946;
  wire  _EVAL_947;
  wire  _EVAL_950;
  wire [31:0] _EVAL_951;
  wire [2:0] _EVAL_952;
  wire [5:0] _EVAL_953;
  wire  _EVAL_954;
  wire [3:0] _EVAL_955;
  wire  _EVAL_957;
  wire [7:0] _EVAL_958;
  wire  _EVAL_959;
  wire  _EVAL_960;
  reg [2:0] _EVAL_961;
  reg [31:0] _RAND_33;
  wire  _EVAL_962;
  wire  _EVAL_963;
  wire  _EVAL_964;
  wire [46:0] _EVAL_965;
  wire  _EVAL_966;
  wire  _EVAL_967;
  wire [5:0] _EVAL_968;
  wire [5:0] _EVAL_969;
  wire  _EVAL_971;
  wire  _EVAL_972;
  wire [31:0] _EVAL_973;
  reg  _EVAL_975;
  reg [31:0] _RAND_34;
  wire [32:0] _EVAL_976;
  wire  _EVAL_977;
  reg  _EVAL_978;
  reg [31:0] _RAND_35;
  wire [2:0] _EVAL_979;
  wire  _EVAL_981;
  wire  _EVAL_982;
  wire [4:0] _EVAL_983;
  wire  _EVAL_984;
  wire  _EVAL_985;
  wire  _EVAL_988;
  wire [46:0] _EVAL_989;
  wire  _EVAL_990;
  wire  _EVAL_991;
  wire [3:0] _EVAL_992;
  wire  _EVAL_993;
  wire  _EVAL_995;
  wire [3:0] _EVAL_996;
  wire [32:0] _EVAL_997;
  reg [5:0] _EVAL_998;
  reg [31:0] _RAND_36;
  wire  _EVAL_999;
  wire [7:0] _EVAL_1000;
  wire [7:0] _EVAL_1001;
  wire [5:0] _EVAL_1002;
  wire [7:0] _EVAL_1003;
  wire [7:0] _EVAL_1004;
  wire [31:0] _EVAL_1006;
  reg  _EVAL_1008;
  reg [31:0] _RAND_37;
  wire [5:0] _EVAL_1009;
  wire  _EVAL_1010;
  wire [5:0] _EVAL_1011;
  wire  _EVAL_1012;
  wire [46:0] _EVAL_1013;
  wire [5:0] _EVAL_1014;
  wire  _EVAL_1016;
  wire  _EVAL_1017;
  wire  _EVAL_1018;
  wire [31:0] _EVAL_1021;
  wire [6:0] _EVAL_1022;
  wire [32:0] _EVAL_1023;
  wire  _EVAL_1024;
  wire  _EVAL_1025;
  wire  _EVAL_1026;
  assign _EVAL_410 = _EVAL_554 | _EVAL_914;
  assign _EVAL_173 = _EVAL_857 ? _EVAL_388 : 89'h0;
  assign _EVAL_830 = _EVAL_171 ? _EVAL_403 : _EVAL_838;
  assign _EVAL_82 = _EVAL_528[1:0];
  assign _EVAL_912 = {_EVAL_192, 3'h0};
  assign _EVAL_1024 = _EVAL_869 | _EVAL_348;
  assign _EVAL_522 = $signed(_EVAL_224) & 33'shc0008000;
  assign _EVAL_288 = {1'b0,$signed(_EVAL_1021)};
  assign _EVAL_681 = _EVAL_559 | _EVAL_438;
  assign _EVAL_696 = _EVAL_660[2:0];
  assign _EVAL_190 = _EVAL_729[7:1];
  assign _EVAL_204 = _EVAL_613[5:2];
  assign _EVAL_755 = _EVAL_273 & _EVAL_179;
  assign _EVAL_924 = _EVAL_74 & _EVAL_830;
  assign _EVAL_915 = _EVAL_355 & _EVAL_876;
  assign _EVAL_327 = _EVAL_814 & _EVAL_345;
  assign _EVAL_503 = {_EVAL_813, 1'h0};
  assign _EVAL_268 = _EVAL_375[1];
  assign _EVAL_144 = _EVAL_485 | _EVAL_937;
  assign _EVAL_694 = {{1'd0}, _EVAL_241};
  assign _EVAL_276 = _EVAL_1012 & _EVAL_962;
  assign _EVAL_278 = _EVAL_249 ? _EVAL_614 : 6'h0;
  assign _EVAL_808 = _EVAL_555 & _EVAL_460;
  assign _EVAL_888 = _EVAL_96 & _EVAL_892;
  assign _EVAL_675 = _EVAL_122 & _EVAL_1012;
  assign _EVAL_624 = _EVAL_518 & _EVAL_982;
  assign _EVAL_991 = _EVAL_195 | _EVAL_479;
  assign _EVAL_464 = _EVAL_690 == 2'h1;
  assign _EVAL_592 = _EVAL_785 & _EVAL_458;
  assign _EVAL_292 = _EVAL_279 & _EVAL_888;
  assign _EVAL_859 = _EVAL_583 | _EVAL_682;
  assign _EVAL_49 = _EVAL_462[38];
  assign _EVAL_416 = $signed(_EVAL_804) & 33'shc0008000;
  assign _EVAL_450 = _EVAL_23 & _EVAL_371;
  assign _EVAL_408 = _EVAL_480 & _EVAL_855;
  assign _EVAL_632 = _EVAL_940 ? _EVAL_378 : _EVAL_480;
  assign _EVAL_367 = {_EVAL_245,_EVAL_179,_EVAL_532,_EVAL_250};
  assign _EVAL_892 = _EVAL_472 ? _EVAL_749 : _EVAL_679;
  assign _EVAL_338 = _EVAL_472 ? _EVAL_768 : _EVAL_275;
  assign _EVAL_499 = {_EVAL_422, 1'h0};
  assign _EVAL_211 = _EVAL & _EVAL_543;
  assign _EVAL_939 = _EVAL_1016 & _EVAL_277;
  assign _EVAL_382 = _EVAL_967 & _EVAL_344;
  assign _EVAL_644 = {_EVAL_460,_EVAL_754,_EVAL_675};
  assign _EVAL_502 = _EVAL_476 & _EVAL_675;
  assign _EVAL_571 = _EVAL_975 & _EVAL_876;
  assign _EVAL_187 = _EVAL_452 != 3'h0;
  assign _EVAL_596 = _EVAL_208[5:0];
  assign _EVAL_452 = {_EVAL_890,_EVAL_348,_EVAL_869};
  assign _EVAL_997 = _EVAL_500;
  assign _EVAL_457 = _EVAL_577 ? _EVAL_198 : 6'h0;
  assign _EVAL_785 = _EVAL_969[5:3];
  assign _EVAL_371 = _EVAL_93 == 3'h4;
  assign _EVAL_341 = {_EVAL_22,2'h0,_EVAL_369,_EVAL_25,2'h0,_EVAL_132,1'h0};
  assign _EVAL_886 = _EVAL_903 ? _EVAL_915 : _EVAL_975;
  assign _EVAL_374 = _EVAL_15 == 3'h4;
  assign _EVAL_626 = _EVAL_434 ? _EVAL_798 : 89'h0;
  assign _EVAL_375 = ~_EVAL_539;
  assign _EVAL_799 = _EVAL_28 & _EVAL_448;
  assign _EVAL_602 = _EVAL_23 & _EVAL_212;
  assign _EVAL_98 = _EVAL_691[33];
  assign _EVAL_684 = _EVAL_983[3:0];
  assign _EVAL_552 = _EVAL_112[0];
  assign _EVAL_587 = _EVAL_811[5:0];
  assign _EVAL_515 = $signed(_EVAL_504) == 33'sh0;
  assign _EVAL_41 = _EVAL_498[36:33];
  assign _EVAL_299 = _EVAL_762 & _EVAL_640;
  assign _EVAL_251 = _EVAL_613 | _EVAL_746;
  assign _EVAL_100 = _EVAL_321[75:44];
  assign _EVAL_470 = _EVAL_96 & _EVAL_837;
  assign _EVAL_230 = _EVAL_414 | _EVAL_357;
  assign _EVAL_277 = _EVAL_274 != 3'h0;
  assign _EVAL_524 = _EVAL_435 | _EVAL_467;
  assign _EVAL_922 = _EVAL_330[5:0];
  assign _EVAL_206 = _EVAL_269 & _EVAL_197;
  assign _EVAL_769 = {{1'd0}, _EVAL_550};
  assign _EVAL_66 = _EVAL_462[0];
  assign _EVAL_687 = _EVAL_440 & _EVAL_707;
  assign _EVAL_946 = _EVAL_768 ? _EVAL_614 : 6'h0;
  assign _EVAL_566 = _EVAL_408 | _EVAL_377;
  assign _EVAL_809 = _EVAL_125 & _EVAL_943;
  assign _EVAL_837 = _EVAL_472 ? _EVAL_226 : _EVAL_777;
  assign _EVAL_720 = _EVAL_160 & _EVAL_394;
  assign _EVAL_435 = _EVAL_813 | _EVAL_203;
  assign _EVAL_348 = _EVAL_0 & _EVAL_638;
  assign _EVAL_92 = _EVAL_462[82:79];
  assign _EVAL_730 = _EVAL_852[5:2];
  assign _EVAL_127 = _EVAL_882 | _EVAL_481;
  assign _EVAL_164 = _EVAL_111 & _EVAL_990;
  assign _EVAL_955 = _EVAL_282 & _EVAL_424;
  assign _EVAL_628 = _EVAL_751[7:2];
  assign _EVAL_791 = _EVAL_578[5:1];
  assign _EVAL_313 = _EVAL_497 ? _EVAL_866 : _EVAL_1008;
  assign _EVAL_761 = _EVAL_496 | _EVAL_178;
  assign _EVAL_574 = _EVAL_523[5:2];
  assign _EVAL_424 = _EVAL_235[3:0];
  assign _EVAL_1009 = _EVAL_765 | _EVAL_678;
  assign _EVAL_420 = _EVAL_356;
  assign _EVAL_768 = _EVAL_324 & _EVAL_869;
  assign _EVAL_917 = _EVAL_368 | _EVAL_421;
  assign _EVAL_174 = _EVAL_171 ? _EVAL_220 : _EVAL_373;
  assign _EVAL_765 = {{2'd0}, _EVAL_256};
  assign _EVAL_31 = _EVAL_462[39];
  assign _EVAL_869 = _EVAL_122 & _EVAL_878;
  assign _EVAL_147 = _EVAL_291 ? _EVAL_900 : _EVAL_988;
  assign _EVAL_985 = _EVAL_291 ? _EVAL_176 : _EVAL_771;
  assign _EVAL_311 = _EVAL_167;
  assign _EVAL_762 = _EVAL_497 & _EVAL_45;
  assign _EVAL_541 = _EVAL_921 | _EVAL_788;
  assign _EVAL_947 = _EVAL_111 & _EVAL_981;
  assign _EVAL_107 = _EVAL_462[43];
  assign _EVAL_84 = _EVAL_655[0];
  assign _EVAL_784 = _EVAL_367 | _EVAL_1014;
  assign _EVAL_976 = _EVAL_180;
  assign _EVAL_252 = _EVAL_903 ? _EVAL_268 : _EVAL_847;
  assign _EVAL_564 = _EVAL_331 ? _EVAL_577 : _EVAL_334;
  assign _EVAL_384 = _EVAL_661[0];
  assign _EVAL_131 = _EVAL_466[41:38];
  assign _EVAL_487 = _EVAL_332 & _EVAL_675;
  assign _EVAL_671 = _EVAL_898[7:2];
  assign _EVAL_473 = _EVAL_268 & _EVAL_307;
  assign _EVAL_324 = _EVAL_362[0];
  assign _EVAL_488 = {1'b0,$signed(_EVAL_456)};
  assign _EVAL_908 = {{2'd0}, _EVAL_406};
  assign _EVAL_386 = _EVAL_784 | _EVAL_824;
  assign _EVAL_64 = _EVAL_883 | _EVAL_363;
  assign _EVAL_220 = _EVAL_440[0];
  assign _EVAL_175 = _EVAL_513[2];
  assign _EVAL_963 = _EVAL_661[1];
  assign _EVAL_474 = _EVAL_846 ? _EVAL_538 : 6'h0;
  assign _EVAL_306 = ~_EVAL_501;
  assign _EVAL_778 = ~_EVAL_958;
  assign _EVAL_678 = _EVAL_636 ? _EVAL_538 : 6'h0;
  assign _EVAL_598 = _EVAL_907[7:2];
  assign _EVAL_32 = _EVAL_331 ? _EVAL_802 : _EVAL_861;
  assign _EVAL_236 = $signed(_EVAL_906) == 33'sh0;
  assign _EVAL_622 = _EVAL_242 | _EVAL_677;
  assign _EVAL_459 = _EVAL_531 | _EVAL_471;
  assign _EVAL_872 = _EVAL_375 & _EVAL_274;
  assign _EVAL_905 = {{2'd0}, _EVAL_730};
  assign _EVAL_879 = _EVAL_513[1];
  assign _EVAL_38 = _EVAL_691[43:42];
  assign _EVAL_467 = _EVAL_820[2:0];
  assign _EVAL_233 = _EVAL_121[0];
  assign _EVAL_776 = _EVAL_593 & _EVAL_950;
  assign _EVAL_806 = _EVAL_331 ? _EVAL_881 : _EVAL_555;
  assign _EVAL_437 = _EVAL_313 ? _EVAL_341 : 47'h0;
  assign _EVAL_682 = {_EVAL_652, 3'h0};
  assign _EVAL_763 = _EVAL_291 & _EVAL_125;
  assign _EVAL_510 = _EVAL_125 & _EVAL_893;
  assign _EVAL_721 = _EVAL_877[2:0];
  assign _EVAL_99 = _EVAL_462[32:1];
  assign _EVAL_634 = _EVAL_23 & _EVAL_967;
  assign _EVAL_330 = _EVAL_642 - _EVAL_409;
  assign _EVAL_340 = _EVAL_735[5:0];
  assign _EVAL_243 = $signed(_EVAL_415) & 33'shc0008000;
  assign _EVAL_612 = _EVAL_847 & _EVAL_307;
  assign _EVAL_451 = {_EVAL_430,_EVAL_634,_EVAL_380,_EVAL_259,_EVAL_855};
  assign _EVAL_355 = _EVAL_375[0];
  assign _EVAL_757 = _EVAL_687 | _EVAL_381;
  assign _EVAL_640 = _EVAL_557 != 4'h0;
  assign _EVAL_988 = _EVAL_681 | _EVAL_959;
  assign _EVAL_804 = {1'b0,$signed(_EVAL_601)};
  assign _EVAL_283 = _EVAL_940 ? _EVAL_636 : _EVAL_610;
  assign _EVAL_256 = _EVAL_803 ? _EVAL_186 : 4'h0;
  assign _EVAL_195 = _EVAL_515 & _EVAL_211;
  assign _EVAL_767 = _EVAL_366 | _EVAL_319;
  assign _EVAL_828 = {1'b0,$signed(_EVAL_136)};
  assign _EVAL_773 = _EVAL_1022[5:0];
  assign _EVAL_188 = _EVAL_639[0];
  assign _EVAL_493 = _EVAL_45 & _EVAL_1018;
  assign _EVAL_898 = ~_EVAL_627;
  assign _EVAL_142 = _EVAL_321[36:33];
  assign _EVAL_811 = _EVAL_998 - _EVAL_447;
  assign _EVAL_817 = {_EVAL_611, 4'h0};
  assign _EVAL_909 = ~_EVAL_961;
  assign _EVAL_995 = _EVAL_276 | _EVAL_848;
  assign _EVAL_794 = _EVAL_497 ? _EVAL_846 : _EVAL_453;
  assign _EVAL_520 = _EVAL_125 & _EVAL_392;
  assign _EVAL_267 = _EVAL_28 & _EVAL_772;
  assign _EVAL_601 = _EVAL_136 ^ 32'h40000000;
  assign _EVAL_802 = _EVAL_398 | _EVAL_460;
  assign _EVAL_1004 = _EVAL_585 | _EVAL_1001;
  assign _EVAL_406 = _EVAL_617 ? _EVAL_186 : 4'h0;
  assign _EVAL_983 = {_EVAL_783, 1'h0};
  assign _EVAL_700 = _EVAL_451 | _EVAL_901;
  assign _EVAL_389 = _EVAL_706 != 4'h0;
  assign _EVAL_760 = _EVAL_443 == 2'h0;
  assign _EVAL_546 = _EVAL_855 | _EVAL_259;
  assign _EVAL_739 = _EVAL_784[5:2];
  assign _EVAL_594 = _EVAL_580[7:1];
  assign _EVAL_896 = $signed(_EVAL_976) == 33'sh0;
  assign _EVAL_439 = _EVAL_915 ? _EVAL_614 : 6'h0;
  assign _EVAL_196 = $signed(_EVAL_828) & 33'shc0008000;
  assign _EVAL_322 = _EVAL_96 & _EVAL_379;
  assign _EVAL_543 = _EVAL_331 ? _EVAL_879 : _EVAL_334;
  assign _EVAL_984 = _EVAL_291 ? _EVAL_271 : _EVAL_342;
  assign _EVAL_495 = _EVAL_938 | _EVAL_1011;
  assign _EVAL_216 = _EVAL_422 | _EVAL_889;
  assign _EVAL_981 = _EVAL_903 ? _EVAL_258 : _EVAL_656;
  assign _EVAL_870 = _EVAL_610 & _EVAL_634;
  assign _EVAL_889 = _EVAL_499[2:0];
  assign _EVAL_658 = _EVAL_940 ? _EVAL_803 : _EVAL_454;
  assign _EVAL_573 = _EVAL_871 | _EVAL_199;
  assign _EVAL_941 = {_EVAL_71,_EVAL_150,_EVAL_104,_EVAL_33,_EVAL_115,_EVAL_110,_EVAL_155};
  assign _EVAL_343 = _EVAL_569;
  assign _EVAL_943 = _EVAL_291 ? _EVAL_285 : _EVAL_771;
  assign _EVAL_509 = _EVAL_234 | _EVAL_179;
  assign _EVAL_781 = {{5'd0}, _EVAL_842};
  assign _EVAL_298 = {_EVAL_216, 2'h0};
  assign _EVAL_954 = _EVAL_707 != 3'h0;
  assign _EVAL_570 = $signed(_EVAL_927) == 33'sh0;
  assign _EVAL_212 = _EVAL_575 == 2'h0;
  assign _EVAL_562 = {_EVAL_744, 1'h0};
  assign _EVAL_519 = _EVAL_639 & _EVAL_826;
  assign _EVAL_388 = {_EVAL_86,_EVAL_135,_EVAL_120,_EVAL_222,_EVAL_136,_EVAL_13,_EVAL_1,_EVAL_73,_EVAL_364};
  assign _EVAL_409 = {{5'd0}, _EVAL_657};
  assign _EVAL_881 = _EVAL_175 & _EVAL_460;
  assign _EVAL_193 = _EVAL_373 & _EVAL_250;
  assign _EVAL_241 = _EVAL_793[5:1];
  assign _EVAL_1021 = _EVAL_58 ^ 32'h80008000;
  assign _EVAL_882 = _EVAL_1017 | _EVAL_534;
  assign _EVAL_312 = _EVAL_946 | _EVAL_968;
  assign _EVAL_633 = _EVAL_374 & _EVAL_1026;
  assign _EVAL_979 = _EVAL_216 | _EVAL_529;
  assign _EVAL_792 = _EVAL_236 | _EVAL_202;
  assign _EVAL_349 = {{1'd0}, _EVAL_69};
  assign _EVAL_250 = _EVAL_122 & _EVAL_761;
  assign _EVAL_661 = ~_EVAL_955;
  assign _EVAL_146 = _EVAL_643 | _EVAL_633;
  assign _EVAL_641 = _EVAL_717[2:0];
  assign _EVAL_965 = _EVAL_283 ? _EVAL_483 : 47'h0;
  assign _EVAL_705 = _EVAL_148 & _EVAL_860;
  assign _EVAL_248 = {{2'd0}, _EVAL_14};
  assign _EVAL_990 = _EVAL_903 ? _EVAL_672 : _EVAL_518;
  assign _EVAL_542 = _EVAL_851 & _EVAL_387;
  assign _EVAL_280 = _EVAL_760 & _EVAL_168;
  assign _EVAL_796 = {1'b0,$signed(_EVAL_262)};
  assign _EVAL_315 = ~_EVAL_999;
  assign _EVAL_821 = _EVAL_757 | _EVAL_527;
  assign _EVAL_362 = ~_EVAL_490;
  assign _EVAL_456 = _EVAL_136 ^ 32'h80008000;
  assign _EVAL_271 = _EVAL_963 & _EVAL_316;
  assign _EVAL_310 = _EVAL_171 & _EVAL_74;
  assign _EVAL_1018 = _EVAL_497 ? _EVAL_718 : _EVAL_453;
  assign _EVAL_88 = _EVAL_655[42];
  assign _EVAL_689 = _EVAL_945[5:0];
  assign _EVAL_385 = _EVAL_274 & _EVAL_944;
  assign _EVAL_848 = _EVAL_878 & _EVAL_322;
  assign _EVAL_982 = _EVAL_97 & _EVAL_295;
  assign _EVAL_4 = _EVAL_545 | _EVAL_358;
  assign _EVAL_723 = _EVAL_443 == 2'h1;
  assign _EVAL_525 = ~_EVAL_957;
  assign _EVAL_938 = _EVAL_702 | _EVAL_457;
  assign _EVAL_344 = _EVAL_28 & _EVAL_548;
  assign _EVAL_959 = _EVAL_771 & _EVAL_450;
  assign _EVAL_960 = _EVAL_310 & _EVAL_954;
  assign _EVAL_996 = _EVAL_414[5:2];
  assign _EVAL_228 = _EVAL_477[3:0];
  assign _EVAL_477 = {_EVAL_519, 1'h0};
  assign _EVAL_558 = _EVAL_291 ? _EVAL_384 : _EVAL_600;
  assign _EVAL_865 = _EVAL_639[3];
  assign _EVAL_329 = _EVAL_331 ? _EVAL_802 : _EVAL_861;
  assign _EVAL_356 = $signed(_EVAL_396) & 33'shc0008000;
  assign _EVAL_966 = _EVAL_212 & _EVAL_493;
  assign _EVAL_819 = _EVAL_714[7:4];
  assign _EVAL_551 = _EVAL_442 | _EVAL_989;
  assign _EVAL_890 = _EVAL_97 & _EVAL_279;
  assign _EVAL_683 = _EVAL_171 ? _EVAL_509 : _EVAL_169;
  assign _EVAL_526 = _EVAL_371 & _EVAL_809;
  assign _EVAL_746 = {{2'd0}, _EVAL_204};
  assign _EVAL_320 = {{1'd0}, _EVAL_894};
  assign _EVAL_609 = {_EVAL_242, 2'h0};
  assign _EVAL_925 = _EVAL & _EVAL_214;
  assign _EVAL_637 = _EVAL_349 | 2'h2;
  assign _EVAL_899 = _EVAL_895 - _EVAL_433;
  assign _EVAL_972 = _EVAL_325 | _EVAL_854;
  assign _EVAL_911 = {{5'd0}, _EVAL_833};
  assign _EVAL_62 = _EVAL_836[0];
  assign _EVAL_829 = _EVAL_353 | _EVAL_868;
  assign _EVAL_934 = _EVAL_384 & _EVAL_705;
  assign _EVAL_185 = {1'b0,$signed(_EVAL_50)};
  assign _EVAL_673 = _EVAL_708[3:0];
  assign _EVAL_787 = _EVAL_331 & _EVAL;
  assign _EVAL_208 = 21'h3f << _EVAL_284;
  assign _EVAL_754 = _EVAL_0 & _EVAL_515;
  assign _EVAL_537 = {{1'd0}, _EVAL_621};
  assign _EVAL_358 = _EVAL_418 & _EVAL_924;
  assign _EVAL_76 = _EVAL_462[41];
  assign _EVAL_404 = _EVAL_832 | _EVAL_673;
  assign _EVAL_106 = _EVAL_691[46:44];
  assign _EVAL_716 = 23'hff << _EVAL_6;
  assign _EVAL_621 = _EVAL_703[7:1];
  assign _EVAL_481 = _EVAL_792 & _EVAL_607;
  assign _EVAL_26 = _EVAL_462[40];
  assign _EVAL_623 = _EVAL_564 ? _EVAL_798 : 89'h0;
  assign _EVAL_171 = _EVAL_213 == 6'h0;
  assign _EVAL_539 = _EVAL_952 & _EVAL_641;
  assign _EVAL_289 = _EVAL_896 & _EVAL_925;
  assign _EVAL_932 = ~_EVAL_659;
  assign _EVAL_253 = _EVAL_261 ? _EVAL_388 : 89'h0;
  assign _EVAL_532 = _EVAL_0 & _EVAL_418;
  assign _EVAL_659 = _EVAL_402[7:0];
  assign _EVAL_370 = _EVAL_562[3:0];
  assign _EVAL_590 = _EVAL_1002[5:1];
  assign _EVAL_224 = {1'b0,$signed(_EVAL_973)};
  assign _EVAL_210 = _EVAL_661[2];
  assign _EVAL_648 = _EVAL_644 & _EVAL_232;
  assign _EVAL_309 = _EVAL_923 ? _EVAL_186 : 4'h0;
  assign _EVAL_432 = _EVAL_822[1];
  assign _EVAL_851 = _EVAL_859[5:3];
  assign _EVAL_971 = _EVAL_290 & _EVAL_651;
  assign _EVAL_1013 = _EVAL_632 ? _EVAL_341 : 47'h0;
  assign _EVAL_818 = _EVAL_608[7:1];
  assign _EVAL_638 = $signed(_EVAL_789) == 33'sh0;
  assign _EVAL_77 = _EVAL_498[32:1];
  assign _EVAL_693 = _EVAL_321[82:79];
  assign _EVAL_738 = _EVAL_15[2:1];
  assign _EVAL_63 = _EVAL_691[0];
  assign _EVAL_442 = _EVAL_437 | _EVAL_347;
  assign _EVAL_803 = _EVAL_770 & _EVAL_380;
  assign _EVAL_664 = _EVAL_399 | _EVAL_474;
  assign _EVAL_545 = _EVAL_991 | _EVAL_206;
  assign _EVAL_398 = _EVAL_675 | _EVAL_754;
  assign _EVAL_625 = {{2'd0}, _EVAL_163};
  assign _EVAL_261 = _EVAL_331 ? _EVAL_487 : _EVAL_476;
  assign _EVAL_429 = _EVAL_148 & _EVAL_645;
  assign _EVAL_258 = _EVAL_1010 | _EVAL_982;
  assign _EVAL_651 = _EVAL_28 & _EVAL_553;
  assign _EVAL_383 = _EVAL_1008 & _EVAL_429;
  assign _EVAL_209 = _EVAL_486 ? _EVAL_839 : 89'h0;
  assign _EVAL_290 = _EVAL_738 == 2'h1;
  assign _EVAL_363 = _EVAL_761 & _EVAL_615;
  assign _EVAL_402 = 23'hff << _EVAL_141;
  assign _EVAL_314 = _EVAL_567 | _EVAL_992;
  assign _EVAL_707 = {_EVAL_179,_EVAL_532,_EVAL_250};
  assign _EVAL_70 = _EVAL_498[88:86];
  assign _EVAL_993 = $signed(_EVAL_997) == 33'sh0;
  assign _EVAL_489 = _EVAL_899[5:0];
  assign _EVAL_876 = _EVAL_122 & _EVAL_200;
  assign _EVAL_394 = _EVAL_101 == 3'h4;
  assign _EVAL_319 = _EVAL_658 ? _EVAL_728 : 47'h0;
  assign _EVAL_198 = _EVAL_315 ? _EVAL_628 : 6'h0;
  assign _EVAL_618 = _EVAL_819 & _EVAL_397;
  assign _EVAL_153 = _EVAL_680[2:0];
  assign _EVAL_835 = _EVAL_263 ? _EVAL_635 : 6'h0;
  assign _EVAL_605 = _EVAL_571 | _EVAL_612;
  assign _EVAL_300 = _EVAL_672 & _EVAL_982;
  assign _EVAL_430 = _EVAL_826 & _EVAL_530;
  assign _EVAL_871 = _EVAL_464 & _EVAL_799;
  assign _EVAL_620 = _EVAL_806 ? _EVAL_839 : 89'h0;
  assign _EVAL_273 = _EVAL_440[2];
  assign _EVAL_657 = _EVAL_28 & _EVAL_257;
  assign _EVAL_904 = _EVAL_763 & _EVAL_389;
  assign _EVAL_878 = $signed(_EVAL_853) == 33'sh0;
  assign _EVAL_465 = _EVAL_497 ? _EVAL_183 : _EVAL_1008;
  assign _EVAL_704 = {{2'd0}, _EVAL_598};
  assign _EVAL_440 = ~_EVAL_592;
  assign _EVAL_380 = _EVAL_160 & _EVAL_723;
  assign _EVAL_67 = _EVAL_836[34];
  assign _EVAL_1016 = _EVAL_903 & _EVAL_111;
  assign _EVAL_223 = _EVAL_667 ? _EVAL_184 : 47'h0;
  assign _EVAL_887 = _EVAL_565 | _EVAL_727;
  assign _EVAL_43 = _EVAL_462[88:86];
  assign _EVAL_528 = _EVAL_498[82:79];
  assign _EVAL_1022 = _EVAL_494 - _EVAL_731;
  assign _EVAL_392 = _EVAL_291 ? _EVAL_900 : _EVAL_988;
  assign _EVAL_269 = $signed(_EVAL_343) == 33'sh0;
  assign _EVAL_184 = {_EVAL_30,2'h0,_EVAL_726,_EVAL_15,2'h0,_EVAL_72,1'h0};
  assign _EVAL_790 = 23'hff << _EVAL_120;
  assign _EVAL_726 = {{2'd0}, _EVAL_95};
  assign _EVAL_868 = _EVAL_318 ? _EVAL_798 : 89'h0;
  assign _EVAL_257 = _EVAL_940 ? _EVAL_205 : _EVAL_964;
  assign _EVAL_214 = _EVAL_331 ? _EVAL_175 : _EVAL_555;
  assign _EVAL_842 = _EVAL_74 & _EVAL_683;
  assign _EVAL_1025 = _EVAL_403 & _EVAL_532;
  assign _EVAL_861 = _EVAL_797 | _EVAL_808;
  assign _EVAL_733 = _EVAL_171 ? _EVAL_755 : _EVAL_563;
  assign _EVAL_507 = _EVAL_491[7:1];
  assign _EVAL_914 = _EVAL_427 ? _EVAL_798 : 89'h0;
  assign _EVAL_65 = _EVAL_655[36:33];
  assign _EVAL_919 = $signed(_EVAL_185) & 33'shc0000000;
  assign _EVAL_397 = _EVAL_714[3:0];
  assign _EVAL_751 = ~_EVAL_469;
  assign _EVAL_662 = _EVAL_600 & _EVAL_705;
  assign _EVAL_849 = _EVAL_462[75:44];
  assign _EVAL_710 = _EVAL_860 & _EVAL_413;
  assign _EVAL_207 = _EVAL_291 ? _EVAL_617 : _EVAL_737;
  assign _EVAL_743 = _EVAL_903 ? _EVAL_355 : _EVAL_975;
  assign _EVAL_786 = ~_EVAL_376;
  assign _EVAL_222 = {{1'd0}, _EVAL_637};
  assign _EVAL_202 = $signed(_EVAL_240) == 33'sh0;
  assign _EVAL_498 = _EVAL_516 | _EVAL_620;
  assign _EVAL_1001 = {_EVAL_361, 4'h0};
  assign _EVAL_926 = _EVAL_822[2];
  assign _EVAL_433 = {{5'd0}, _EVAL_470};
  assign _EVAL_462 = _EVAL_712 | _EVAL_722;
  assign _EVAL_712 = _EVAL_173 | _EVAL_626;
  assign _EVAL_323 = $signed(_EVAL_488) & 33'shc0008000;
  assign _EVAL_834 = _EVAL_917 | _EVAL_670;
  assign _EVAL_157 = _EVAL_466[0];
  assign _EVAL_833 = _EVAL_45 & _EVAL_653;
  assign _EVAL_414 = _EVAL_391 | _EVAL_769;
  assign _EVAL_81 = _EVAL_472 ? _EVAL_226 : _EVAL_777;
  assign _EVAL_391 = {_EVAL_385,_EVAL_982,_EVAL_307,_EVAL_876};
  assign _EVAL_742 = _EVAL_872 | _EVAL_696;
  assign _EVAL_1000 = {{2'd0}, _EVAL_441};
  assign _EVAL_964 = _EVAL_823 | _EVAL_870;
  assign _EVAL_39 = _EVAL_691[32:1];
  assign _EVAL_284 = {{1'd0}, _EVAL_34};
  assign _EVAL_708 = {_EVAL_832, 2'h0};
  assign _EVAL_78 = _EVAL_655[85:83];
  assign _EVAL_485 = _EVAL_685 | _EVAL_280;
  assign _EVAL_744 = _EVAL_822 & _EVAL_557;
  assign _EVAL_989 = _EVAL_753 ? _EVAL_728 : 47'h0;
  assign _EVAL_114 = _EVAL_321[88:86];
  assign _EVAL_568 = _EVAL_331 ? _EVAL_332 : _EVAL_476;
  assign _EVAL_307 = _EVAL_0 & _EVAL_269;
  assign _EVAL_860 = _EVAL_25 == 3'h4;
  assign _EVAL_653 = _EVAL_497 ? _EVAL_701 : _EVAL_541;
  assign _EVAL_264 = _EVAL_193 | _EVAL_514;
  assign _EVAL_643 = _EVAL_971 | _EVAL_425;
  assign _EVAL_295 = $signed(_EVAL_758) == 33'sh0;
  assign _EVAL_11 = _EVAL_691[41:38];
  assign _EVAL_585 = {{1'd0}, _EVAL_818};
  assign _EVAL_219 = _EVAL_111 & _EVAL_743;
  assign _EVAL_303 = _EVAL_497 ? _EVAL_432 : _EVAL_492;
  assign _EVAL_44 = _EVAL_655[37];
  assign _EVAL_285 = _EVAL_661[3];
  assign _EVAL_357 = {{2'd0}, _EVAL_996};
  assign _EVAL_281 = _EVAL_451[7:1];
  assign _EVAL_1006 = _EVAL_58 ^ 32'h40000000;
  assign _EVAL_347 = _EVAL_511 ? _EVAL_184 : 47'h0;
  assign _EVAL_852 = _EVAL_793 | _EVAL_694;
  assign _EVAL_126 = _EVAL_466[34];
  assign _EVAL_316 = _EVAL_37 & _EVAL_374;
  assign _EVAL_753 = _EVAL_497 ? _EVAL_923 : _EVAL_665;
  assign _EVAL_180 = $signed(_EVAL_796) & 33'shc0008000;
  assign _EVAL_460 = _EVAL_97 & _EVAL_896;
  assign _EVAL_506 = _EVAL_45 & _EVAL_465;
  assign _EVAL_378 = _EVAL_188 & _EVAL_855;
  assign _EVAL_181 = {{1'd0}, _EVAL_297};
  assign _EVAL_10 = _EVAL_655[78:76];
  assign _EVAL_893 = _EVAL_291 ? _EVAL_210 : _EVAL_737;
  assign _EVAL_479 = _EVAL_638 & _EVAL_177;
  assign _EVAL_282 = _EVAL_235[7:4];
  assign _EVAL_850 = {1'b0,$signed(_EVAL_58)};
  assign _EVAL_254 = _EVAL_87[2];
  assign _EVAL_366 = _EVAL_1013 | _EVAL_223;
  assign _EVAL_205 = _EVAL_885 | _EVAL_634;
  assign _EVAL_443 = _EVAL_101[2:1];
  assign _EVAL_513 = ~_EVAL_542;
  assign _EVAL_855 = _EVAL_148 & _EVAL_464;
  assign _EVAL_550 = _EVAL_391[5:1];
  assign _EVAL_772 = _EVAL_940 ? _EVAL_770 : _EVAL_454;
  assign _EVAL_992 = _EVAL_711[3:0];
  assign _EVAL_645 = _EVAL_690 == 2'h0;
  assign _EVAL_950 = _EVAL_826 != 4'h0;
  assign _EVAL_270 = _EVAL_742 | _EVAL_393;
  assign _EVAL_544 = _EVAL_37 & _EVAL_227;
  assign _EVAL_575 = _EVAL_93[2:1];
  assign _EVAL_654 = _EVAL_639[1];
  assign _EVAL_714 = _EVAL_918 | _EVAL_817;
  assign _EVAL_952 = _EVAL_717[5:3];
  assign _EVAL_614 = _EVAL_525 ? _EVAL_671 : 6'h0;
  assign _EVAL_393 = _EVAL_595[2:0];
  assign _EVAL_244 = _EVAL_492 & _EVAL_544;
  assign _EVAL_577 = _EVAL_879 & _EVAL_754;
  assign _EVAL_379 = _EVAL_472 ? _EVAL_324 : _EVAL_275;
  assign _EVAL_103 = _EVAL_321[0];
  assign _EVAL_1026 = _EVAL_125 & _EVAL_165;
  assign _EVAL_608 = _EVAL_907 | _EVAL_704;
  assign _EVAL_491 = _EVAL_700 | _EVAL_1003;
  assign _EVAL_381 = _EVAL_560[2:0];
  assign _EVAL_297 = _EVAL_251[5:1];
  assign _EVAL_291 = _EVAL_998 == 6'h0;
  assign _EVAL_422 = _EVAL_513 & _EVAL_644;
  assign _EVAL_158 = _EVAL_466[33];
  assign _EVAL_534 = _EVAL_295 & _EVAL_164;
  assign _EVAL_583 = {{1'd0}, _EVAL_791};
  assign _EVAL_567 = _EVAL_744 | _EVAL_370;
  assign _EVAL_201 = {1'b0,$signed(_EVAL_1006)};
  assign _EVAL_885 = _EVAL_546 | _EVAL_380;
  assign _EVAL_247 = _EVAL_50 ^ 32'h80008000;
  assign _EVAL_123 = _EVAL_466[32:1];
  assign _EVAL_504 = _EVAL_536;
  assign _EVAL_668 = _EVAL_557 & _EVAL_586;
  assign _EVAL_527 = _EVAL_863[2:0];
  assign _EVAL_617 = _EVAL_210 & _EVAL_720;
  assign _EVAL_672 = _EVAL_375[2];
  assign _EVAL_701 = _EVAL_972 | _EVAL_602;
  assign _EVAL_536 = $signed(_EVAL_260) & 33'shc0008000;
  assign _EVAL_530 = ~_EVAL_611;
  assign _EVAL_170 = 23'hff << _EVAL_52;
  assign _EVAL_42 = _EVAL_655[39];
  assign _EVAL_242 = _EVAL_783 | _EVAL_684;
  assign _EVAL_927 = _EVAL_942;
  assign _EVAL_874 = {{1'd0}, _EVAL_841};
  assign _EVAL_732 = _EVAL_213 - _EVAL_781;
  assign _EVAL_516 = _EVAL_253 | _EVAL_623;
  assign _EVAL_19 = _EVAL_466[43:42];
  assign _EVAL_798 = {_EVAL_128,_EVAL_79,_EVAL_52,_EVAL_248,_EVAL_58,_EVAL_149,_EVAL_46,_EVAL_94,_EVAL_941};
  assign _EVAL_788 = _EVAL_453 & _EVAL_602;
  assign _EVAL_907 = _EVAL_729 | _EVAL_619;
  assign _EVAL_53 = _EVAL_655[88:86];
  assign _EVAL_441 = _EVAL_296[7:2];
  assign _EVAL_572 = _EVAL_629 ? _EVAL_839 : 89'h0;
  assign _EVAL_937 = _EVAL_394 & _EVAL_510;
  assign _EVAL_711 = {_EVAL_567, 2'h0};
  assign _EVAL_747 = _EVAL_473 ? _EVAL_198 : 6'h0;
  assign _EVAL_923 = _EVAL_926 & _EVAL_854;
  assign _EVAL_548 = _EVAL_940 ? _EVAL_865 : _EVAL_610;
  assign _EVAL_325 = _EVAL_429 | _EVAL_544;
  assign _EVAL_354 = _EVAL_654 & _EVAL_259;
  assign _EVAL_529 = _EVAL_298[2:0];
  assign _EVAL_2 = _EVAL_498[85:83];
  assign _EVAL_129 = _EVAL_466[46:44];
  assign _EVAL_421 = _EVAL_984 ? _EVAL_184 : 47'h0;
  assign _EVAL_752 = _EVAL_985 ? _EVAL_483 : 47'h0;
  assign _EVAL_627 = _EVAL_790[7:0];
  assign _EVAL_836 = _EVAL_551 | _EVAL_606;
  assign _EVAL_396 = {1'b0,$signed(_EVAL_247)};
  assign _EVAL_666 = _EVAL_383 | _EVAL_244;
  assign _EVAL_579 = _EVAL_200 & _EVAL_219;
  assign _EVAL_246 = _EVAL_439 | _EVAL_747;
  assign _EVAL_359 = _EVAL_405 & _EVAL_348;
  assign _EVAL_942 = $signed(_EVAL_850) & 33'shc0000000;
  assign _EVAL_54 = _EVAL_655[43];
  assign _EVAL_232 = ~_EVAL_652;
  assign _EVAL_973 = _EVAL_50 ^ 32'h40000000;
  assign _EVAL_944 = ~_EVAL_192;
  assign _EVAL_165 = _EVAL_291 ? _EVAL_963 : _EVAL_342;
  assign _EVAL_900 = _EVAL_649 | _EVAL_450;
  assign _EVAL_703 = {_EVAL_401,_EVAL_450,_EVAL_720,_EVAL_316,_EVAL_705};
  assign _EVAL_500 = $signed(_EVAL_850) & 33'shc0008000;
  assign _EVAL_722 = _EVAL_733 ? _EVAL_839 : 89'h0;
  assign _EVAL_403 = _EVAL_440[1];
  assign _EVAL_364 = {_EVAL_55,_EVAL_12,_EVAL_20,_EVAL_133,_EVAL_7,_EVAL_83,_EVAL_48};
  assign _EVAL_677 = _EVAL_609[3:0];
  assign _EVAL_810 = _EVAL_625 | 3'h4;
  assign _EVAL_231 = _EVAL_644 != 3'h0;
  assign _EVAL_296 = _EVAL_703 | _EVAL_537;
  assign _EVAL_301 = _EVAL_342 & _EVAL_316;
  assign _EVAL_512 = _EVAL_432 & _EVAL_544;
  assign _EVAL_80 = _EVAL_498[0];
  assign _EVAL_824 = {{2'd0}, _EVAL_739};
  assign _EVAL_5 = _EVAL_462[42];
  assign _EVAL_929 = _EVAL & _EVAL_329;
  assign _EVAL_667 = _EVAL_940 ? _EVAL_354 : _EVAL_978;
  assign _EVAL_199 = _EVAL_645 & _EVAL_506;
  assign _EVAL_631 = _EVAL_472 & _EVAL_96;
  assign _EVAL_649 = _EVAL_540 | _EVAL_720;
  assign _EVAL_669 = _EVAL_367[5:1];
  assign _EVAL_262 = _EVAL_50 ^ 32'h80000000;
  assign _EVAL_630 = _EVAL_778[7:2];
  assign _EVAL_369 = {{2'd0}, _EVAL_8};
  assign _EVAL_438 = _EVAL_737 & _EVAL_720;
  assign _EVAL_1002 = {_EVAL_346,_EVAL_890,_EVAL_348,_EVAL_869};
  assign _EVAL_877 = _EVAL_181 | _EVAL_843;
  assign _EVAL_822 = ~_EVAL_327;
  assign _EVAL_448 = _EVAL_940 ? _EVAL_188 : _EVAL_480;
  assign _EVAL_999 = _EVAL_128[2];
  assign _EVAL_9 = _EVAL_171 ? _EVAL_509 : _EVAL_169;
  assign _EVAL_235 = _EVAL_845 | _EVAL_724;
  assign _EVAL_255 = _EVAL_563 & _EVAL_179;
  assign _EVAL_578 = _EVAL_852 | _EVAL_905;
  assign _EVAL_603 = {_EVAL_138,_EVAL_108,_EVAL_90,_EVAL_119,_EVAL_61,_EVAL_85,_EVAL_91};
  assign _EVAL_514 = _EVAL_838 & _EVAL_532;
  assign _EVAL_279 = $signed(_EVAL_420) == 33'sh0;
  assign _EVAL_168 = _EVAL_45 & _EVAL_779;
  assign _EVAL_346 = _EVAL_452 & _EVAL_909;
  assign _EVAL_770 = _EVAL_639[2];
  assign _EVAL_425 = _EVAL_227 & _EVAL_756;
  assign _EVAL_130 = _EVAL_462[36:33];
  assign _EVAL_735 = _EVAL_674 - _EVAL_953;
  assign _EVAL_977 = _EVAL_382 | _EVAL_966;
  assign _EVAL_249 = _EVAL_220 & _EVAL_250;
  assign _EVAL_294 = _EVAL_787 & _EVAL_231;
  assign _EVAL_203 = _EVAL_503[2:0];
  assign _EVAL_695 = _EVAL_732[5:0];
  assign _EVAL_234 = _EVAL_250 | _EVAL_532;
  assign _EVAL_846 = _EVAL_718 & _EVAL_602;
  assign _EVAL_866 = _EVAL_183 & _EVAL_429;
  assign _EVAL_461 = _EVAL_454 & _EVAL_380;
  assign _EVAL_557 = {_EVAL_602,_EVAL_854,_EVAL_544,_EVAL_429};
  assign _EVAL_145 = _EVAL_286[0];
  assign _EVAL_401 = _EVAL_706 & _EVAL_786;
  assign _EVAL_21 = _EVAL_462[37];
  assign _EVAL_599 = _EVAL_709 ? _EVAL_835 : 6'h0;
  assign _EVAL_727 = _EVAL_646 & _EVAL_348;
  assign _EVAL_724 = {_EVAL_376, 4'h0};
  assign _EVAL_565 = _EVAL_275 & _EVAL_869;
  assign _EVAL_820 = {_EVAL_435, 2'h0};
  assign _EVAL_777 = _EVAL_887 | _EVAL_239;
  assign _EVAL_517 = _EVAL_665 & _EVAL_854;
  assign _EVAL_580 = _EVAL_296 | _EVAL_1000;
  assign _EVAL_156 = _EVAL_940 ? _EVAL_205 : _EVAL_964;
  assign _EVAL_482 = $signed(_EVAL_288) & 33'shc0008000;
  assign _EVAL_616 = _EVAL_176 ? _EVAL_538 : 6'h0;
  assign _EVAL_1023 = $signed(_EVAL_185) & 33'shc0008000;
  assign _EVAL_940 = _EVAL_642 == 6'h0;
  assign _EVAL_472 = _EVAL_895 == 6'h0;
  assign _EVAL_756 = _EVAL_45 & _EVAL_303;
  assign _EVAL_921 = _EVAL_666 | _EVAL_517;
  assign _EVAL_1017 = _EVAL_289 | _EVAL_292;
  assign _EVAL_840 = _EVAL_334 & _EVAL_754;
  assign _EVAL_967 = _EVAL_575 == 2'h1;
  assign _EVAL_759 = _EVAL_836[37:35];
  assign _EVAL_717 = _EVAL_874 | _EVAL_912;
  assign _EVAL_918 = {{1'd0}, _EVAL_507};
  assign _EVAL_540 = _EVAL_705 | _EVAL_316;
  assign _EVAL_706 = {_EVAL_450,_EVAL_720,_EVAL_316,_EVAL_705};
  assign _EVAL_353 = _EVAL_886 ? _EVAL_388 : 89'h0;
  assign _EVAL_511 = _EVAL_497 ? _EVAL_512 : _EVAL_492;
  assign _EVAL_35 = _EVAL_321[78:76];
  assign _EVAL_789 = _EVAL_482;
  assign _EVAL_331 = _EVAL_674 == 6'h0;
  assign _EVAL_227 = _EVAL_738 == 2'h0;
  assign _EVAL_857 = _EVAL_171 ? _EVAL_249 : _EVAL_373;
  assign _EVAL_418 = _EVAL_993 | _EVAL_570;
  assign _EVAL_854 = _EVAL_160 & _EVAL_760;
  assign _EVAL_655 = _EVAL_829 | _EVAL_209;
  assign _EVAL_415 = {1'b0,$signed(_EVAL_951)};
  assign _EVAL_906 = _EVAL_1023;
  assign _EVAL_197 = _EVAL_111 & _EVAL_252;
  assign _EVAL_538 = _EVAL_552 ? _EVAL_630 : 6'h0;
  assign _EVAL_434 = _EVAL_171 ? _EVAL_1025 : _EVAL_838;
  assign _EVAL_731 = {{5'd0}, _EVAL_947};
  assign _EVAL_102 = _EVAL_498[75:44];
  assign _EVAL_613 = _EVAL_1002 | _EVAL_328;
  assign _EVAL_709 = _EVAL_749 & _EVAL_890;
  assign _EVAL_1012 = $signed(_EVAL_931) == 33'sh0;
  assign _EVAL_427 = _EVAL_472 ? _EVAL_359 : _EVAL_646;
  assign _EVAL_894 = _EVAL_386[5:1];
  assign _EVAL_179 = _EVAL_97 & _EVAL_792;
  assign _EVAL_161 = _EVAL_977 | _EVAL_526;
  assign _EVAL_715 = _EVAL_312 | _EVAL_599;
  assign _EVAL_328 = {{1'd0}, _EVAL_590};
  assign _EVAL_584 = _EVAL_196;
  assign _EVAL_595 = {_EVAL_742, 2'h0};
  assign _EVAL_478 = _EVAL_58 ^ 32'h80000000;
  assign _EVAL_200 = $signed(_EVAL_750) == 33'sh0;
  assign _EVAL_68 = _EVAL_698[30:0];
  assign _EVAL_962 = _EVAL & _EVAL_568;
  assign _EVAL_656 = _EVAL_605 | _EVAL_624;
  assign _EVAL_891 = _EVAL_171 ? _EVAL_273 : _EVAL_563;
  assign _EVAL_286 = _EVAL_691[37:35];
  assign _EVAL_405 = _EVAL_362[1];
  assign _EVAL_483 = {_EVAL_112,_EVAL_143,_EVAL_6,_EVAL_93,_EVAL_152,_EVAL_36,_EVAL_117,_EVAL_109};
  assign _EVAL_670 = _EVAL_207 ? _EVAL_728 : 47'h0;
  assign _EVAL_814 = _EVAL_1004[7:4];
  assign _EVAL_377 = _EVAL_978 & _EVAL_259;
  assign _EVAL_629 = _EVAL_472 ? _EVAL_709 : _EVAL_679;
  assign _EVAL_1010 = _EVAL_876 | _EVAL_307;
  assign _EVAL_51 = _EVAL_462[78:76];
  assign _EVAL_718 = _EVAL_822[3];
  assign _EVAL_458 = _EVAL_969[2:0];
  assign _EVAL_901 = {{1'd0}, _EVAL_281};
  assign _EVAL_554 = _EVAL_338 ? _EVAL_388 : 89'h0;
  assign _EVAL_447 = {{5'd0}, _EVAL_520};
  assign _EVAL_783 = _EVAL_661 & _EVAL_706;
  assign _EVAL_615 = _EVAL_74 & _EVAL_174;
  assign _EVAL_903 = _EVAL_494 == 6'h0;
  assign _EVAL_118 = _EVAL_498[78:76];
  assign _EVAL_569 = $signed(_EVAL_201) & 33'shc0008000;
  assign _EVAL_559 = _EVAL_662 | _EVAL_301;
  assign _EVAL_593 = _EVAL_940 & _EVAL_28;
  assign _EVAL_843 = {_EVAL_961, 3'h0};
  assign _EVAL_1014 = {{1'd0}, _EVAL_669};
  assign _EVAL_969 = _EVAL_320 | _EVAL_884;
  assign _EVAL_27 = _EVAL_321[85:83];
  assign _EVAL_239 = _EVAL_679 & _EVAL_890;
  assign _EVAL_497 = _EVAL_351 == 6'h0;
  assign _EVAL_560 = {_EVAL_687, 1'h0};
  assign _EVAL_496 = $signed(_EVAL_584) == 33'sh0;
  assign _EVAL_690 = _EVAL_25[2:1];
  assign _EVAL_116 = _EVAL_573 | _EVAL_710;
  assign _EVAL_931 = _EVAL_243;
  assign _EVAL_56 = _EVAL_903 ? _EVAL_258 : _EVAL_656;
  assign _EVAL_863 = {_EVAL_757, 2'h0};
  assign _EVAL_169 = _EVAL_264 | _EVAL_255;
  assign _EVAL_740 = _EVAL_246 | _EVAL_862;
  assign _EVAL_466 = _EVAL_834 | _EVAL_752;
  assign _EVAL_240 = _EVAL_919;
  assign _EVAL_167 = $signed(_EVAL_828) & 33'shc0000000;
  assign _EVAL_749 = _EVAL_362[2];
  assign _EVAL_691 = _EVAL_767 | _EVAL_965;
  assign _EVAL_24 = _EVAL_691[34];
  assign _EVAL_685 = _EVAL_723 & _EVAL_267;
  assign _EVAL_660 = {_EVAL_872, 1'h0};
  assign _EVAL_702 = _EVAL_487 ? _EVAL_614 : 6'h0;
  assign _EVAL_826 = {_EVAL_634,_EVAL_380,_EVAL_259,_EVAL_855};
  assign _EVAL_825 = _EVAL_877[5:3];
  assign _EVAL_936 = _EVAL_291 ? _EVAL_934 : _EVAL_600;
  assign _EVAL_318 = _EVAL_903 ? _EVAL_473 : _EVAL_847;
  assign _EVAL_140 = _EVAL_836[46:44];
  assign _EVAL_531 = _EVAL_278 | _EVAL_225;
  assign _EVAL_953 = {{5'd0}, _EVAL_929};
  assign _EVAL_387 = _EVAL_859[2:0];
  assign _EVAL_57 = _EVAL_655[32:1];
  assign _EVAL_957 = _EVAL_86[2];
  assign _EVAL_845 = {{1'd0}, _EVAL_594};
  assign _EVAL_636 = _EVAL_865 & _EVAL_634;
  assign _EVAL_274 = {_EVAL_982,_EVAL_307,_EVAL_876};
  assign _EVAL_841 = _EVAL_230[5:1];
  assign _EVAL_1011 = _EVAL_881 ? _EVAL_835 : 6'h0;
  assign _EVAL_945 = _EVAL_351 - _EVAL_911;
  assign _EVAL_968 = _EVAL_359 ? _EVAL_198 : 6'h0;
  assign _EVAL_883 = _EVAL_995 | _EVAL_579;
  assign _EVAL_823 = _EVAL_566 | _EVAL_461;
  assign _EVAL_226 = _EVAL_1024 | _EVAL_890;
  assign _EVAL_698 = _EVAL_655[75:44];
  assign _EVAL_1003 = {{2'd0}, _EVAL_221};
  assign _EVAL_606 = _EVAL_794 ? _EVAL_483 : 47'h0;
  assign _EVAL_221 = _EVAL_700[7:2];
  assign _EVAL_178 = $signed(_EVAL_311) == 33'sh0;
  assign _EVAL_413 = _EVAL_125 & _EVAL_558;
  assign _EVAL_29 = _EVAL_693[1:0];
  assign _EVAL_779 = _EVAL_497 ? _EVAL_926 : _EVAL_665;
  assign _EVAL_750 = _EVAL_416;
  assign _EVAL_586 = ~_EVAL_361;
  assign _EVAL_18 = _EVAL_497 ? _EVAL_701 : _EVAL_541;
  assign _EVAL_177 = _EVAL_96 & _EVAL_597;
  assign _EVAL_832 = _EVAL_519 | _EVAL_228;
  assign _EVAL_884 = {_EVAL_501, 3'h0};
  assign _EVAL_105 = _EVAL_836[41:38];
  assign _EVAL_728 = {_EVAL_121,_EVAL_59,_EVAL_284,_EVAL_101,_EVAL_47,_EVAL_124,_EVAL_134,_EVAL_40};
  assign _EVAL_619 = {{1'd0}, _EVAL_190};
  assign _EVAL_729 = {_EVAL_668,_EVAL_602,_EVAL_854,_EVAL_544,_EVAL_429};
  assign _EVAL_259 = _EVAL_37 & _EVAL_290;
  assign _EVAL_260 = {1'b0,$signed(_EVAL_478)};
  assign _EVAL_183 = _EVAL_822[0];
  assign _EVAL_862 = _EVAL_300 ? _EVAL_835 : 6'h0;
  assign _EVAL_463 = _EVAL_908 | _EVAL_616;
  assign _EVAL_469 = _EVAL_170[7:0];
  assign _EVAL_839 = {_EVAL_87,_EVAL_89,_EVAL_141,_EVAL_810,_EVAL_50,_EVAL_75,_EVAL_139,_EVAL_113,_EVAL_603};
  assign _EVAL_151 = _EVAL_836[33];
  assign _EVAL_597 = _EVAL_472 ? _EVAL_405 : _EVAL_646;
  assign _EVAL_176 = _EVAL_285 & _EVAL_450;
  assign _EVAL_345 = _EVAL_1004[3:0];
  assign _EVAL_607 = _EVAL_74 & _EVAL_891;
  assign _EVAL_635 = _EVAL_932[7:2];
  assign _EVAL_523 = ~_EVAL_596;
  assign _EVAL_951 = _EVAL_136 ^ 32'h80000000;
  assign _EVAL_263 = ~_EVAL_254;
  assign _EVAL_639 = ~_EVAL_618;
  assign _EVAL_853 = _EVAL_323;
  assign _EVAL_225 = _EVAL_1025 ? _EVAL_198 : 6'h0;
  assign _EVAL_17 = _EVAL_836[43:42];
  assign _EVAL_60 = _EVAL_836[32:1];
  assign _EVAL_471 = _EVAL_755 ? _EVAL_835 : 6'h0;
  assign _EVAL_793 = {_EVAL_648,_EVAL_460,_EVAL_754,_EVAL_675};
  assign _EVAL_332 = _EVAL_513[0];
  assign _EVAL_321 = _EVAL_410 | _EVAL_572;
  assign _EVAL_676 = _EVAL_631 & _EVAL_187;
  assign _EVAL_399 = {{2'd0}, _EVAL_309};
  assign _EVAL_159 = _EVAL_759[0];
  assign _EVAL_797 = _EVAL_502 | _EVAL_840;
  assign _EVAL_486 = _EVAL_903 ? _EVAL_300 : _EVAL_518;
  assign _EVAL_758 = _EVAL_522;
  assign _EVAL_490 = _EVAL_825 & _EVAL_721;
  assign _EVAL_680 = _EVAL_655[82:79];
  assign _EVAL_16 = _EVAL_321[32:1];
  assign _EVAL_186 = _EVAL_233 ? _EVAL_574 : 4'h0;
  assign _EVAL_553 = _EVAL_940 ? _EVAL_654 : _EVAL_978;
  assign _EVAL_813 = _EVAL_362 & _EVAL_452;
  assign _EVAL_3 = _EVAL_849[29:0];
  assign _EVAL_137 = _EVAL_462[85:83];
  assign _EVAL_958 = _EVAL_716[7:0];
  assign _EVAL_245 = _EVAL_707 & _EVAL_306;
  assign _EVAL_368 = _EVAL_936 ? _EVAL_341 : 47'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_192 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_213 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_275 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_334 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_342 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_351 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_361 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_373 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_376 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_453 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_454 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_476 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_480 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_492 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_494 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_501 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_518 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_555 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_563 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_600 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_610 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_611 = _RAND_21[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_642 = _RAND_22[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_646 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_652 = _RAND_24[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_665 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_674 = _RAND_26[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_679 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_737 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_771 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_838 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_847 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_895 = _RAND_32[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_961 = _RAND_33[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_975 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_978 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_998 = _RAND_36[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_1008 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_162) begin
    if (_EVAL_154) begin
      _EVAL_192 <= 3'h7;
    end else if (_EVAL_939) begin
      _EVAL_192 <= _EVAL_270;
    end
    if (_EVAL_154) begin
      _EVAL_213 <= 6'h0;
    end else if (_EVAL_310) begin
      _EVAL_213 <= _EVAL_459;
    end else begin
      _EVAL_213 <= _EVAL_695;
    end
    if (_EVAL_154) begin
      _EVAL_275 <= 1'h0;
    end else if (_EVAL_472) begin
      _EVAL_275 <= _EVAL_768;
    end
    if (_EVAL_154) begin
      _EVAL_334 <= 1'h0;
    end else if (_EVAL_331) begin
      _EVAL_334 <= _EVAL_577;
    end
    if (_EVAL_154) begin
      _EVAL_342 <= 1'h0;
    end else if (_EVAL_291) begin
      _EVAL_342 <= _EVAL_271;
    end
    if (_EVAL_154) begin
      _EVAL_351 <= 6'h0;
    end else if (_EVAL_762) begin
      _EVAL_351 <= _EVAL_664;
    end else begin
      _EVAL_351 <= _EVAL_689;
    end
    if (_EVAL_154) begin
      _EVAL_361 <= 4'hf;
    end else if (_EVAL_299) begin
      _EVAL_361 <= _EVAL_314;
    end
    if (_EVAL_154) begin
      _EVAL_373 <= 1'h0;
    end else if (_EVAL_171) begin
      _EVAL_373 <= _EVAL_249;
    end
    if (_EVAL_154) begin
      _EVAL_376 <= 4'hf;
    end else if (_EVAL_904) begin
      _EVAL_376 <= _EVAL_622;
    end
    if (_EVAL_154) begin
      _EVAL_453 <= 1'h0;
    end else if (_EVAL_497) begin
      _EVAL_453 <= _EVAL_846;
    end
    if (_EVAL_154) begin
      _EVAL_454 <= 1'h0;
    end else if (_EVAL_940) begin
      _EVAL_454 <= _EVAL_803;
    end
    if (_EVAL_154) begin
      _EVAL_476 <= 1'h0;
    end else if (_EVAL_331) begin
      _EVAL_476 <= _EVAL_487;
    end
    if (_EVAL_154) begin
      _EVAL_480 <= 1'h0;
    end else if (_EVAL_940) begin
      _EVAL_480 <= _EVAL_378;
    end
    if (_EVAL_154) begin
      _EVAL_492 <= 1'h0;
    end else if (_EVAL_497) begin
      _EVAL_492 <= _EVAL_512;
    end
    if (_EVAL_154) begin
      _EVAL_494 <= 6'h0;
    end else if (_EVAL_1016) begin
      _EVAL_494 <= _EVAL_740;
    end else begin
      _EVAL_494 <= _EVAL_773;
    end
    if (_EVAL_154) begin
      _EVAL_501 <= 3'h7;
    end else if (_EVAL_960) begin
      _EVAL_501 <= _EVAL_821;
    end
    if (_EVAL_154) begin
      _EVAL_518 <= 1'h0;
    end else if (_EVAL_903) begin
      _EVAL_518 <= _EVAL_300;
    end
    if (_EVAL_154) begin
      _EVAL_555 <= 1'h0;
    end else if (_EVAL_331) begin
      _EVAL_555 <= _EVAL_881;
    end
    if (_EVAL_154) begin
      _EVAL_563 <= 1'h0;
    end else if (_EVAL_171) begin
      _EVAL_563 <= _EVAL_755;
    end
    if (_EVAL_154) begin
      _EVAL_600 <= 1'h0;
    end else if (_EVAL_291) begin
      _EVAL_600 <= _EVAL_934;
    end
    if (_EVAL_154) begin
      _EVAL_610 <= 1'h0;
    end else if (_EVAL_940) begin
      _EVAL_610 <= _EVAL_636;
    end
    if (_EVAL_154) begin
      _EVAL_611 <= 4'hf;
    end else if (_EVAL_776) begin
      _EVAL_611 <= _EVAL_404;
    end
    if (_EVAL_154) begin
      _EVAL_642 <= 6'h0;
    end else if (_EVAL_593) begin
      _EVAL_642 <= _EVAL_1009;
    end else begin
      _EVAL_642 <= _EVAL_922;
    end
    if (_EVAL_154) begin
      _EVAL_646 <= 1'h0;
    end else if (_EVAL_472) begin
      _EVAL_646 <= _EVAL_359;
    end
    if (_EVAL_154) begin
      _EVAL_652 <= 3'h7;
    end else if (_EVAL_294) begin
      _EVAL_652 <= _EVAL_979;
    end
    if (_EVAL_154) begin
      _EVAL_665 <= 1'h0;
    end else if (_EVAL_497) begin
      _EVAL_665 <= _EVAL_923;
    end
    if (_EVAL_154) begin
      _EVAL_674 <= 6'h0;
    end else if (_EVAL_787) begin
      _EVAL_674 <= _EVAL_495;
    end else begin
      _EVAL_674 <= _EVAL_340;
    end
    if (_EVAL_154) begin
      _EVAL_679 <= 1'h0;
    end else if (_EVAL_472) begin
      _EVAL_679 <= _EVAL_709;
    end
    if (_EVAL_154) begin
      _EVAL_737 <= 1'h0;
    end else if (_EVAL_291) begin
      _EVAL_737 <= _EVAL_617;
    end
    if (_EVAL_154) begin
      _EVAL_771 <= 1'h0;
    end else if (_EVAL_291) begin
      _EVAL_771 <= _EVAL_176;
    end
    if (_EVAL_154) begin
      _EVAL_838 <= 1'h0;
    end else if (_EVAL_171) begin
      _EVAL_838 <= _EVAL_1025;
    end
    if (_EVAL_154) begin
      _EVAL_847 <= 1'h0;
    end else if (_EVAL_903) begin
      _EVAL_847 <= _EVAL_473;
    end
    if (_EVAL_154) begin
      _EVAL_895 <= 6'h0;
    end else if (_EVAL_631) begin
      _EVAL_895 <= _EVAL_715;
    end else begin
      _EVAL_895 <= _EVAL_489;
    end
    if (_EVAL_154) begin
      _EVAL_961 <= 3'h7;
    end else if (_EVAL_676) begin
      _EVAL_961 <= _EVAL_524;
    end
    if (_EVAL_154) begin
      _EVAL_975 <= 1'h0;
    end else if (_EVAL_903) begin
      _EVAL_975 <= _EVAL_915;
    end
    if (_EVAL_154) begin
      _EVAL_978 <= 1'h0;
    end else if (_EVAL_940) begin
      _EVAL_978 <= _EVAL_354;
    end
    if (_EVAL_154) begin
      _EVAL_998 <= 6'h0;
    end else if (_EVAL_763) begin
      _EVAL_998 <= _EVAL_463;
    end else begin
      _EVAL_998 <= _EVAL_587;
    end
    if (_EVAL_154) begin
      _EVAL_1008 <= 1'h0;
    end else if (_EVAL_497) begin
      _EVAL_1008 <= _EVAL_866;
    end
  end
endmodule
