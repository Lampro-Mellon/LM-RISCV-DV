//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_95(
  output [1:0]  _EVAL,
  output        _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  output        _EVAL_3,
  input         _EVAL_4,
  output [3:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  input  [31:0] _EVAL_7,
  output [31:0] _EVAL_8,
  input         _EVAL_9,
  output [2:0]  _EVAL_10,
  output        _EVAL_11,
  input         _EVAL_12,
  input  [29:0] _EVAL_13,
  output [1:0]  _EVAL_14,
  output        _EVAL_15,
  output [2:0]  _EVAL_16,
  input         _EVAL_17,
  output [29:0] _EVAL_18,
  output        _EVAL_19,
  input  [2:0]  _EVAL_20,
  input  [1:0]  _EVAL_21,
  output [2:0]  _EVAL_22,
  output        _EVAL_23,
  input  [3:0]  _EVAL_24,
  output        _EVAL_25,
  input         _EVAL_26,
  input  [31:0] _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input  [2:0]  _EVAL_32,
  output        _EVAL_33,
  input         _EVAL_34,
  input  [2:0]  _EVAL_35,
  output        _EVAL_36,
  output [1:0]  _EVAL_37,
  output [2:0]  _EVAL_38,
  input         _EVAL_39,
  input  [1:0]  _EVAL_40,
  input  [1:0]  _EVAL_41,
  output        _EVAL_42,
  input         _EVAL_43,
  output        _EVAL_44,
  output [2:0]  _EVAL_45,
  output [31:0] _EVAL_46,
  input  [2:0]  _EVAL_47,
  output        _EVAL_48
);
  assign _EVAL_8 = _EVAL_7;
  assign _EVAL_16 = _EVAL_32;
  assign _EVAL_22 = _EVAL_35;
  assign _EVAL_14 = _EVAL_41;
  assign _EVAL_45 = _EVAL_6;
  assign _EVAL_37 = _EVAL_40;
  assign _EVAL_11 = _EVAL_39;
  assign _EVAL_18 = _EVAL_13;
  assign _EVAL_33 = _EVAL_43;
  assign _EVAL_36 = _EVAL_2;
  assign _EVAL_25 = _EVAL_26;
  assign _EVAL_48 = _EVAL_4;
  assign _EVAL_15 = _EVAL_9;
  assign _EVAL_5 = _EVAL_24;
  assign _EVAL_46 = _EVAL_27;
  assign _EVAL_19 = _EVAL_29;
  assign _EVAL_10 = _EVAL_47;
  assign _EVAL_23 = _EVAL_34;
  assign _EVAL_0 = _EVAL_28;
  assign _EVAL_44 = _EVAL_31;
  assign _EVAL_42 = _EVAL_12;
  assign _EVAL_38 = _EVAL_20;
  assign _EVAL = _EVAL_21;
  assign _EVAL_3 = _EVAL_30;
endmodule
