//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_149(
  output [2:0]  _EVAL,
  input         _EVAL_0,
  input  [6:0]  _EVAL_1,
  input  [31:0] _EVAL_2,
  output        _EVAL_3,
  input  [11:0] _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [1:0]  _EVAL_7,
  input         _EVAL_8,
  output        _EVAL_9,
  input  [3:0]  _EVAL_10,
  output [31:0] _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  output        _EVAL_14,
  output [2:0]  _EVAL_15,
  output [31:0] _EVAL_16,
  input  [1:0]  _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  output [1:0]  _EVAL_20,
  output        _EVAL_21,
  input         _EVAL_22,
  output        _EVAL_23,
  output        _EVAL_24,
  input  [2:0]  _EVAL_25,
  output [1:0]  _EVAL_26,
  output        _EVAL_27,
  input  [31:0] _EVAL_28,
  input  [2:0]  _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32
);
  wire  dmOuter__EVAL;
  wire [8:0] dmOuter__EVAL_0;
  wire [6:0] dmOuter__EVAL_1;
  wire [31:0] dmOuter__EVAL_2;
  wire  dmOuter__EVAL_3;
  wire  dmOuter__EVAL_4;
  wire [2:0] dmOuter__EVAL_5;
  wire  dmOuter__EVAL_6;
  wire  dmOuter__EVAL_7;
  wire  dmOuter__EVAL_8;
  wire  dmOuter__EVAL_9;
  wire  dmOuter__EVAL_10;
  wire [2:0] dmOuter__EVAL_11;
  wire  dmOuter__EVAL_12;
  wire [31:0] dmOuter__EVAL_13;
  wire  dmOuter__EVAL_14;
  wire  dmOuter__EVAL_15;
  wire  dmOuter__EVAL_16;
  wire [1:0] dmOuter__EVAL_17;
  wire  dmOuter__EVAL_18;
  wire  dmOuter__EVAL_19;
  wire  dmOuter__EVAL_20;
  wire [3:0] dmOuter__EVAL_21;
  wire  dmOuter__EVAL_22;
  wire  dmOuter__EVAL_23;
  wire  dmOuter__EVAL_24;
  wire [1:0] dmOuter__EVAL_25;
  wire  dmOuter__EVAL_26;
  wire  dmOuter__EVAL_27;
  wire [31:0] dmOuter__EVAL_28;
  wire [1:0] dmOuter__EVAL_29;
  wire [31:0] dmOuter__EVAL_30;
  wire  dmOuter__EVAL_31;
  wire  dmInner__EVAL;
  wire  dmInner__EVAL_0;
  wire  dmInner__EVAL_1;
  wire  dmInner__EVAL_2;
  wire  dmInner__EVAL_3;
  wire [11:0] dmInner__EVAL_4;
  wire  dmInner__EVAL_5;
  wire  dmInner__EVAL_6;
  wire  dmInner__EVAL_7;
  wire [2:0] dmInner__EVAL_8;
  wire [31:0] dmInner__EVAL_9;
  wire [2:0] dmInner__EVAL_10;
  wire  dmInner__EVAL_11;
  wire  dmInner__EVAL_12;
  wire [31:0] dmInner__EVAL_13;
  wire  dmInner__EVAL_14;
  wire [3:0] dmInner__EVAL_15;
  wire  dmInner__EVAL_16;
  wire [3:0] dmInner__EVAL_17;
  wire [2:0] dmInner__EVAL_18;
  wire [31:0] dmInner__EVAL_19;
  wire  dmInner__EVAL_20;
  wire [31:0] dmInner__EVAL_21;
  wire  dmInner__EVAL_22;
  wire  dmInner__EVAL_23;
  wire [1:0] dmInner__EVAL_24;
  wire [2:0] dmInner__EVAL_25;
  wire [2:0] dmInner__EVAL_26;
  wire [8:0] dmInner__EVAL_27;
  wire  dmInner__EVAL_28;
  wire  dmInner__EVAL_29;
  wire [1:0] dmInner__EVAL_30;
  wire  dmInner__EVAL_31;
  wire [2:0] dmInner__EVAL_32;
  wire  dmInner__EVAL_33;
  wire  dmInner__EVAL_34;
  wire [1:0] dmInner__EVAL_35;
  wire [2:0] dmInner__EVAL_36;
  _EVAL_136 dmOuter (
    ._EVAL(dmOuter__EVAL),
    ._EVAL_0(dmOuter__EVAL_0),
    ._EVAL_1(dmOuter__EVAL_1),
    ._EVAL_2(dmOuter__EVAL_2),
    ._EVAL_3(dmOuter__EVAL_3),
    ._EVAL_4(dmOuter__EVAL_4),
    ._EVAL_5(dmOuter__EVAL_5),
    ._EVAL_6(dmOuter__EVAL_6),
    ._EVAL_7(dmOuter__EVAL_7),
    ._EVAL_8(dmOuter__EVAL_8),
    ._EVAL_9(dmOuter__EVAL_9),
    ._EVAL_10(dmOuter__EVAL_10),
    ._EVAL_11(dmOuter__EVAL_11),
    ._EVAL_12(dmOuter__EVAL_12),
    ._EVAL_13(dmOuter__EVAL_13),
    ._EVAL_14(dmOuter__EVAL_14),
    ._EVAL_15(dmOuter__EVAL_15),
    ._EVAL_16(dmOuter__EVAL_16),
    ._EVAL_17(dmOuter__EVAL_17),
    ._EVAL_18(dmOuter__EVAL_18),
    ._EVAL_19(dmOuter__EVAL_19),
    ._EVAL_20(dmOuter__EVAL_20),
    ._EVAL_21(dmOuter__EVAL_21),
    ._EVAL_22(dmOuter__EVAL_22),
    ._EVAL_23(dmOuter__EVAL_23),
    ._EVAL_24(dmOuter__EVAL_24),
    ._EVAL_25(dmOuter__EVAL_25),
    ._EVAL_26(dmOuter__EVAL_26),
    ._EVAL_27(dmOuter__EVAL_27),
    ._EVAL_28(dmOuter__EVAL_28),
    ._EVAL_29(dmOuter__EVAL_29),
    ._EVAL_30(dmOuter__EVAL_30),
    ._EVAL_31(dmOuter__EVAL_31)
  );
  _EVAL_148 dmInner (
    ._EVAL(dmInner__EVAL),
    ._EVAL_0(dmInner__EVAL_0),
    ._EVAL_1(dmInner__EVAL_1),
    ._EVAL_2(dmInner__EVAL_2),
    ._EVAL_3(dmInner__EVAL_3),
    ._EVAL_4(dmInner__EVAL_4),
    ._EVAL_5(dmInner__EVAL_5),
    ._EVAL_6(dmInner__EVAL_6),
    ._EVAL_7(dmInner__EVAL_7),
    ._EVAL_8(dmInner__EVAL_8),
    ._EVAL_9(dmInner__EVAL_9),
    ._EVAL_10(dmInner__EVAL_10),
    ._EVAL_11(dmInner__EVAL_11),
    ._EVAL_12(dmInner__EVAL_12),
    ._EVAL_13(dmInner__EVAL_13),
    ._EVAL_14(dmInner__EVAL_14),
    ._EVAL_15(dmInner__EVAL_15),
    ._EVAL_16(dmInner__EVAL_16),
    ._EVAL_17(dmInner__EVAL_17),
    ._EVAL_18(dmInner__EVAL_18),
    ._EVAL_19(dmInner__EVAL_19),
    ._EVAL_20(dmInner__EVAL_20),
    ._EVAL_21(dmInner__EVAL_21),
    ._EVAL_22(dmInner__EVAL_22),
    ._EVAL_23(dmInner__EVAL_23),
    ._EVAL_24(dmInner__EVAL_24),
    ._EVAL_25(dmInner__EVAL_25),
    ._EVAL_26(dmInner__EVAL_26),
    ._EVAL_27(dmInner__EVAL_27),
    ._EVAL_28(dmInner__EVAL_28),
    ._EVAL_29(dmInner__EVAL_29),
    ._EVAL_30(dmInner__EVAL_30),
    ._EVAL_31(dmInner__EVAL_31),
    ._EVAL_32(dmInner__EVAL_32),
    ._EVAL_33(dmInner__EVAL_33),
    ._EVAL_34(dmInner__EVAL_34),
    ._EVAL_35(dmInner__EVAL_35),
    ._EVAL_36(dmInner__EVAL_36)
  );
  assign dmInner__EVAL_23 = _EVAL_5;
  assign dmInner__EVAL_20 = _EVAL_18;
  assign dmInner__EVAL_10 = _EVAL_25;
  assign dmOuter__EVAL_17 = dmInner__EVAL_24;
  assign _EVAL_3 = dmOuter__EVAL_12;
  assign dmInner__EVAL_31 = _EVAL_19;
  assign dmInner__EVAL_33 = _EVAL_30;
  assign dmOuter__EVAL_8 = _EVAL_31;
  assign dmOuter__EVAL_1 = _EVAL_1;
  assign dmOuter__EVAL_2 = _EVAL_28;
  assign dmInner__EVAL_22 = dmOuter__EVAL_18;
  assign dmInner__EVAL_27 = dmOuter__EVAL_0;
  assign dmOuter__EVAL_27 = _EVAL_32;
  assign _EVAL_9 = dmInner__EVAL_6;
  assign dmOuter__EVAL_19 = dmInner__EVAL_7;
  assign _EVAL_20 = dmOuter__EVAL_25;
  assign dmOuter__EVAL_29 = _EVAL_17;
  assign _EVAL_21 = dmOuter__EVAL_14;
  assign dmOuter__EVAL_24 = _EVAL_8;
  assign _EVAL_27 = dmOuter__EVAL_15;
  assign dmOuter__EVAL_10 = dmInner__EVAL;
  assign _EVAL = dmInner__EVAL_8;
  assign dmOuter__EVAL_4 = _EVAL_13;
  assign dmInner__EVAL_18 = dmOuter__EVAL_5;
  assign dmInner__EVAL_11 = _EVAL_6;
  assign _EVAL_24 = dmInner__EVAL_12;
  assign dmInner__EVAL_2 = _EVAL_0;
  assign dmInner__EVAL_25 = _EVAL_29;
  assign _EVAL_16 = dmOuter__EVAL_30;
  assign dmOuter__EVAL_13 = dmInner__EVAL_21;
  assign _EVAL_11 = dmInner__EVAL_9;
  assign dmInner__EVAL_1 = dmOuter__EVAL_16;
  assign dmOuter__EVAL_3 = _EVAL_22;
  assign dmInner__EVAL_19 = dmOuter__EVAL_28;
  assign dmOuter__EVAL_9 = dmInner__EVAL_5;
  assign _EVAL_14 = dmOuter__EVAL_26;
  assign dmOuter__EVAL_11 = dmInner__EVAL_26;
  assign dmOuter__EVAL_7 = dmInner__EVAL_16;
  assign _EVAL_15 = dmInner__EVAL_36;
  assign dmInner__EVAL_0 = dmOuter__EVAL_22;
  assign dmInner__EVAL_15 = dmOuter__EVAL_21;
  assign dmInner__EVAL_14 = dmOuter__EVAL;
  assign dmInner__EVAL_32 = _EVAL_12;
  assign dmOuter__EVAL_31 = dmInner__EVAL_34;
  assign dmInner__EVAL_35 = _EVAL_7;
  assign _EVAL_23 = dmOuter__EVAL;
  assign dmInner__EVAL_29 = dmOuter__EVAL_20;
  assign dmInner__EVAL_3 = dmOuter__EVAL_23;
  assign _EVAL_26 = dmInner__EVAL_30;
  assign dmInner__EVAL_4 = _EVAL_4;
  assign dmInner__EVAL_17 = _EVAL_10;
  assign dmInner__EVAL_28 = dmOuter__EVAL_6;
  assign dmInner__EVAL_13 = _EVAL_2;
endmodule
