//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_5_assert(
  input         _EVAL,
  input  [3:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [3:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [3:0]  _EVAL_7,
  input  [2:0]  _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [1:0]  _EVAL_14,
  input  [31:0] _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input  [2:0]  _EVAL_18
);
  wire [32:0] _EVAL_20;
  wire  _EVAL_22;
  wire  _EVAL_23;
  reg [31:0] _EVAL_24;
  reg [31:0] _RAND_0;
  wire [32:0] _EVAL_25;
  reg  _EVAL_26;
  reg [31:0] _RAND_1;
  reg [5:0] _EVAL_27;
  reg [31:0] _RAND_2;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire [1:0] _EVAL_37;
  wire  _EVAL_38;
  wire [1:0] _EVAL_39;
  wire  _EVAL_41;
  wire [32:0] _EVAL_42;
  wire  _EVAL_43;
  wire [32:0] _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire [1:0] _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire [32:0] _EVAL_59;
  wire [7:0] _EVAL_60;
  wire [3:0] _EVAL_61;
  wire  _EVAL_62;
  wire [3:0] _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  reg [2:0] _EVAL_66;
  reg [31:0] _RAND_3;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  reg [5:0] _EVAL_71;
  reg [31:0] _RAND_4;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire [32:0] _EVAL_74;
  wire  _EVAL_75;
  wire [7:0] _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire [6:0] _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire [22:0] _EVAL_87;
  wire  _EVAL_88;
  wire [7:0] _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire [32:0] _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire [5:0] _EVAL_108;
  wire  _EVAL_109;
  wire [32:0] _EVAL_110;
  wire  _EVAL_112;
  wire [31:0] _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire [31:0] _EVAL_116;
  wire [1:0] _EVAL_117;
  wire  _EVAL_118;
  wire [31:0] plusarg_reader_out;
  reg [1:0] _EVAL_120;
  reg [31:0] _RAND_5;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire [5:0] _EVAL_123;
  wire  _EVAL_124;
  wire [32:0] _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_128;
  wire  _EVAL_129;
  reg  _EVAL_130;
  reg [31:0] _RAND_6;
  wire  _EVAL_131;
  wire [1:0] _EVAL_132;
  wire  _EVAL_133;
  wire [32:0] _EVAL_134;
  wire [32:0] _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire [31:0] _EVAL_140;
  wire [32:0] _EVAL_141;
  wire  _EVAL_142;
  wire [1:0] _EVAL_143;
  wire  _EVAL_144;
  wire [32:0] _EVAL_145;
  wire [6:0] _EVAL_146;
  wire [31:0] _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire [7:0] _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire [6:0] _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire [31:0] _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  reg [5:0] _EVAL_180;
  reg [31:0] _RAND_7;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire [32:0] _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire [31:0] _EVAL_193;
  reg [2:0] _EVAL_194;
  reg [31:0] _RAND_8;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire [1:0] _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire [3:0] _EVAL_200;
  wire  _EVAL_201;
  wire [31:0] _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_206;
  wire [1:0] _EVAL_207;
  wire [1:0] _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire [22:0] _EVAL_211;
  wire [1:0] _EVAL_212;
  reg [2:0] _EVAL_213;
  reg [31:0] _RAND_9;
  wire [3:0] _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire [6:0] _EVAL_223;
  wire [5:0] _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  reg  _EVAL_236;
  reg [31:0] _RAND_10;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire [32:0] _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  reg [3:0] _EVAL_243;
  reg [31:0] _RAND_11;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  reg [3:0] _EVAL_252;
  reg [31:0] _RAND_12;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire [32:0] _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire [5:0] _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire [5:0] _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire [32:0] _EVAL_275;
  wire [1:0] _EVAL_276;
  wire  _EVAL_277;
  wire [5:0] _EVAL_278;
  reg [31:0] _EVAL_279;
  reg [31:0] _RAND_13;
  wire  _EVAL_280;
  wire  _EVAL_281;
  reg [5:0] _EVAL_282;
  reg [31:0] _RAND_14;
  wire  _EVAL_283;
  wire [32:0] _EVAL_284;
  wire [1:0] _EVAL_285;
  wire  _EVAL_286;
  reg [1:0] _EVAL_287;
  reg [31:0] _RAND_15;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  reg  _EVAL_304;
  reg [31:0] _RAND_16;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire [31:0] _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire [32:0] _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire  _EVAL_321;
  wire  _EVAL_322;
  wire  _EVAL_323;
  wire  _EVAL_324;
  wire  _EVAL_325;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_250 = _EVAL_174 | _EVAL_172;
  assign _EVAL_125 = $signed(_EVAL_141) & -33'sh2000;
  assign _EVAL_291 = _EVAL_18 == 3'h4;
  assign _EVAL_63 = {_EVAL_283,_EVAL_99,_EVAL_38,_EVAL_221};
  assign _EVAL_25 = $signed(_EVAL_59) & -33'sh1000000;
  assign _EVAL_69 = ~_EVAL_254;
  assign _EVAL_81 = _EVAL_27 - 6'h1;
  assign _EVAL_165 = _EVAL_271 | _EVAL_260;
  assign _EVAL_216 = $signed(_EVAL_42) == 33'sh0;
  assign _EVAL_83 = _EVAL_129 | _EVAL_12;
  assign _EVAL_301 = _EVAL_29 & _EVAL_245;
  assign _EVAL_195 = _EVAL_18 == 3'h1;
  assign _EVAL_210 = _EVAL_154 | _EVAL_12;
  assign _EVAL_39 = _EVAL_117 | _EVAL_120;
  assign _EVAL_325 = _EVAL_324 | _EVAL_12;
  assign _EVAL_84 = _EVAL_78 | _EVAL_12;
  assign _EVAL_146 = _EVAL_180 - 6'h1;
  assign _EVAL_220 = ~_EVAL_45;
  assign _EVAL_90 = _EVAL_185 & _EVAL_308;
  assign _EVAL_23 = _EVAL_18 == 3'h0;
  assign _EVAL_323 = _EVAL_200 == 4'h0;
  assign _EVAL_273 = _EVAL_295 | _EVAL_12;
  assign _EVAL_260 = _EVAL_49 & _EVAL_183;
  assign _EVAL_110 = _EVAL_24 + 32'h1;
  assign _EVAL_312 = _EVAL_198 | _EVAL_12;
  assign _EVAL_86 = _EVAL_271 | _EVAL_103;
  assign _EVAL_263 = _EVAL_143[0];
  assign _EVAL_308 = _EVAL_27 == 6'h0;
  assign _EVAL_191 = ~_EVAL_253;
  assign _EVAL_253 = _EVAL_160 | _EVAL_12;
  assign _EVAL_85 = _EVAL_138 & _EVAL_226;
  assign _EVAL_284 = $signed(_EVAL_92) & -33'sh5000;
  assign _EVAL_197 = ~_EVAL_207;
  assign _EVAL_142 = _EVAL_46 | _EVAL_264;
  assign _EVAL_215 = ~_EVAL_288;
  assign _EVAL_199 = _EVAL_9 & _EVAL_196;
  assign _EVAL_202 = {{24'd0}, _EVAL_89};
  assign _EVAL_53 = _EVAL_232 | _EVAL_12;
  assign _EVAL_173 = _EVAL_71 - 6'h1;
  assign _EVAL_310 = ~_EVAL_281;
  assign _EVAL_59 = {1'b0,$signed(_EVAL_313)};
  assign _EVAL_160 = _EVAL_113 == 32'h0;
  assign _EVAL_133 = _EVAL_8 == 3'h5;
  assign _EVAL_75 = _EVAL_117 != _EVAL_207;
  assign _EVAL_256 = _EVAL_74;
  assign _EVAL_314 = _EVAL_15 == _EVAL_279;
  assign _EVAL_233 = _EVAL_13 == _EVAL_304;
  assign _EVAL_235 = _EVAL_14 == 2'h0;
  assign _EVAL_116 = _EVAL_15 ^ 32'h80000000;
  assign _EVAL_229 = _EVAL_9 & _EVAL_259;
  assign _EVAL_155 = _EVAL_29 | _EVAL_185;
  assign _EVAL_186 = _EVAL_91 | _EVAL_12;
  assign _EVAL_305 = ~_EVAL_17;
  assign _EVAL_122 = $signed(_EVAL_275) == 33'sh0;
  assign _EVAL_153 = _EVAL_208[0];
  assign _EVAL_277 = _EVAL_4 == _EVAL_243;
  assign _EVAL_298 = _EVAL_18 == _EVAL_194;
  assign _EVAL_211 = 23'hff << _EVAL_4;
  assign _EVAL_281 = _EVAL_306 | _EVAL_12;
  assign _EVAL_37 = 2'h1 << _EVAL_2;
  assign _EVAL_232 = _EVAL_18 <= 3'h6;
  assign _EVAL_237 = _EVAL_271 | _EVAL_12;
  assign _EVAL_65 = _EVAL_9 & _EVAL_190;
  assign _EVAL_185 = _EVAL & _EVAL_6;
  assign _EVAL_196 = _EVAL_8 == 3'h3;
  assign _EVAL_105 = ~_EVAL_325;
  assign _EVAL_55 = _EVAL_217 | _EVAL_12;
  assign _EVAL_60 = _EVAL_87[7:0];
  assign _EVAL_248 = ~_EVAL_1;
  assign _EVAL_80 = _EVAL_247 | _EVAL_12;
  assign _EVAL_188 = _EVAL_29 & _EVAL_121;
  assign _EVAL_139 = _EVAL_226 | _EVAL_122;
  assign _EVAL_20 = $signed(_EVAL_134) & -33'sh1000;
  assign _EVAL_152 = _EVAL_9 & _EVAL_31;
  assign _EVAL_274 = _EVAL_178 & _EVAL_220;
  assign _EVAL_168 = _EVAL_15[1];
  assign _EVAL_82 = ~_EVAL_255;
  assign _EVAL_31 = _EVAL_8 == 3'h7;
  assign _EVAL_313 = _EVAL_15 ^ 32'h2000000;
  assign _EVAL_68 = ~_EVAL_210;
  assign _EVAL_140 = _EVAL_15 ^ 32'h40000000;
  assign _EVAL_200 = ~_EVAL_7;
  assign _EVAL_275 = _EVAL_44;
  assign _EVAL_192 = _EVAL_183 & _EVAL_286;
  assign _EVAL_62 = ~_EVAL_58;
  assign _EVAL_299 = ~_EVAL_296;
  assign _EVAL_316 = _EVAL_0 == _EVAL_252;
  assign _EVAL_57 = _EVAL_10 == _EVAL_236;
  assign _EVAL_148 = _EVAL_2 == _EVAL_26;
  assign _EVAL_296 = _EVAL_170 | _EVAL_12;
  assign _EVAL_226 = _EVAL_289 | _EVAL_179;
  assign _EVAL_183 = ~_EVAL_168;
  assign _EVAL_280 = _EVAL_319 | _EVAL_12;
  assign _EVAL_150 = _EVAL_211[7:0];
  assign _EVAL_70 = _EVAL_298 | _EVAL_12;
  assign _EVAL_269 = ~_EVAL_157;
  assign _EVAL_242 = ~_EVAL_102;
  assign _EVAL_241 = _EVAL_323 | _EVAL_12;
  assign _EVAL_157 = _EVAL_30 | _EVAL_12;
  assign _EVAL_293 = _EVAL_251 | _EVAL_12;
  assign _EVAL_100 = ~_EVAL_79;
  assign _EVAL_261 = _EVAL_173[5:0];
  assign _EVAL_245 = _EVAL_282 == 6'h0;
  assign _EVAL_102 = _EVAL_34 | _EVAL_12;
  assign _EVAL_112 = _EVAL_138 & _EVAL_139;
  assign _EVAL_322 = ~_EVAL_237;
  assign _EVAL_257 = _EVAL_3 <= 3'h3;
  assign _EVAL_108 = _EVAL_76[7:2];
  assign _EVAL_249 = ~_EVAL_245;
  assign _EVAL_30 = _EVAL_214 == 4'h0;
  assign _EVAL_124 = ~_EVAL_228;
  assign _EVAL_129 = _EVAL_142 | _EVAL_114;
  assign _EVAL_41 = ~_EVAL_151;
  assign _EVAL_204 = ~_EVAL_309;
  assign _EVAL_162 = ~_EVAL_234;
  assign _EVAL_251 = _EVAL_3 == 3'h0;
  assign _EVAL_272 = ~_EVAL_175;
  assign _EVAL_35 = _EVAL_6 & _EVAL_176;
  assign _EVAL_42 = _EVAL_125;
  assign _EVAL_221 = _EVAL_165 | _EVAL_77;
  assign _EVAL_46 = _EVAL_93 & _EVAL_216;
  assign _EVAL_300 = _EVAL_168 & _EVAL_286;
  assign _EVAL_163 = _EVAL_8 == _EVAL_213;
  assign _EVAL_203 = _EVAL_15[0];
  assign _EVAL_56 = _EVAL_98 & _EVAL_300;
  assign _EVAL_207 = _EVAL_274 ? _EVAL_132 : 2'h0;
  assign _EVAL_136 = _EVAL_263 | _EVAL_12;
  assign _EVAL_38 = _EVAL_165 | _EVAL_51;
  assign _EVAL_218 = ~_EVAL_53;
  assign _EVAL_164 = _EVAL_94 | _EVAL_12;
  assign _EVAL_306 = _EVAL_3 <= 3'h4;
  assign _EVAL_319 = _EVAL_75 | _EVAL_72;
  assign _EVAL_93 = _EVAL_0 <= 4'h6;
  assign _EVAL_52 = _EVAL_6 & _EVAL_45;
  assign _EVAL_115 = _EVAL_6 & _EVAL_291;
  assign _EVAL_172 = _EVAL_24 < plusarg_reader_out;
  assign _EVAL_228 = _EVAL_290 | _EVAL_12;
  assign _EVAL_113 = _EVAL_15 & _EVAL_202;
  assign _EVAL_266 = ~_EVAL_80;
  assign _EVAL_187 = _EVAL_0[0];
  assign _EVAL_159 = _EVAL_9 & _EVAL_219;
  assign _EVAL_255 = _EVAL_257 | _EVAL_12;
  assign _EVAL_309 = _EVAL_8[2];
  assign _EVAL_51 = _EVAL_98 & _EVAL_167;
  assign _EVAL_106 = _EVAL_314 | _EVAL_12;
  assign _EVAL_126 = _EVAL_262 | _EVAL_122;
  assign _EVAL_43 = _EVAL_97 | _EVAL_264;
  assign _EVAL_145 = _EVAL_25;
  assign _EVAL_175 = _EVAL_148 | _EVAL_12;
  assign _EVAL_258 = _EVAL_316 | _EVAL_12;
  assign _EVAL_88 = ~_EVAL_16;
  assign _EVAL_178 = _EVAL_185 & _EVAL_230;
  assign _EVAL_201 = $signed(_EVAL_256) == 33'sh0;
  assign _EVAL_307 = _EVAL_57 | _EVAL_12;
  assign _EVAL_78 = _EVAL_3 <= 3'h1;
  assign _EVAL_123 = _EVAL_81[5:0];
  assign _EVAL_154 = _EVAL_14 != 2'h2;
  assign _EVAL_297 = _EVAL_18 == 3'h5;
  assign _EVAL_107 = _EVAL_235 | _EVAL_12;
  assign _EVAL_166 = _EVAL_6 & _EVAL_195;
  assign _EVAL_176 = _EVAL_18 == 3'h2;
  assign _EVAL_104 = $signed(_EVAL_145) == 33'sh0;
  assign _EVAL_135 = {1'b0,$signed(_EVAL_116)};
  assign _EVAL_217 = _EVAL_3 <= 3'h2;
  assign _EVAL_321 = ~_EVAL_308;
  assign _EVAL_97 = _EVAL_112 | _EVAL_46;
  assign _EVAL_230 = _EVAL_180 == 6'h0;
  assign _EVAL_222 = ~_EVAL_317;
  assign _EVAL_92 = {1'b0,$signed(_EVAL_15)};
  assign _EVAL_303 = ~_EVAL_293;
  assign _EVAL_324 = _EVAL_17 == _EVAL_130;
  assign _EVAL_134 = {1'b0,$signed(_EVAL_147)};
  assign _EVAL_77 = _EVAL_98 & _EVAL_192;
  assign _EVAL_95 = _EVAL_9 & _EVAL_133;
  assign _EVAL_209 = _EVAL_117 != 2'h0;
  assign _EVAL_198 = _EVAL_138 & _EVAL_126;
  assign _EVAL_285 = _EVAL_212 & _EVAL_197;
  assign _EVAL_158 = _EVAL_6 & _EVAL_23;
  assign _EVAL_238 = _EVAL_18[0];
  assign _EVAL_118 = ~_EVAL_315;
  assign _EVAL_61 = ~_EVAL_63;
  assign _EVAL_311 = ~_EVAL_186;
  assign _EVAL_288 = _EVAL_248 | _EVAL_12;
  assign _EVAL_98 = _EVAL_276[0];
  assign _EVAL_144 = ~_EVAL_128;
  assign _EVAL_96 = ~_EVAL_106;
  assign _EVAL_234 = _EVAL_43 | _EVAL_12;
  assign _EVAL_76 = ~_EVAL_150;
  assign _EVAL_302 = _EVAL_9 & _EVAL_137;
  assign _EVAL_184 = _EVAL_8 == 3'h2;
  assign _EVAL_32 = _EVAL_3 != 3'h0;
  assign _EVAL_182 = ~_EVAL_107;
  assign _EVAL_219 = _EVAL_8 == 3'h1;
  assign _EVAL_174 = _EVAL_41 | _EVAL_292;
  assign _EVAL_206 = _EVAL_6 & _EVAL_321;
  assign _EVAL_99 = _EVAL_86 | _EVAL_56;
  assign _EVAL_22 = _EVAL_163 | _EVAL_12;
  assign _EVAL_91 = _EVAL_305 | _EVAL_1;
  assign _EVAL_318 = {1'b0,$signed(_EVAL_177)};
  assign _EVAL_290 = _EVAL_14 == _EVAL_287;
  assign _EVAL_147 = _EVAL_15 ^ 32'h3000;
  assign _EVAL_262 = _EVAL_48 | _EVAL_179;
  assign _EVAL_224 = _EVAL_146[5:0];
  assign _EVAL_161 = ~_EVAL_136;
  assign _EVAL_190 = _EVAL_8 == 3'h0;
  assign _EVAL_79 = _EVAL_233 | _EVAL_12;
  assign _EVAL_317 = _EVAL_250 | _EVAL_12;
  assign _EVAL_286 = ~_EVAL_203;
  assign _EVAL_54 = 2'h1 << _EVAL_187;
  assign _EVAL_189 = _EVAL_20;
  assign _EVAL_292 = plusarg_reader_out == 32'h0;
  assign _EVAL_101 = _EVAL_98 & _EVAL_131;
  assign _EVAL_94 = _EVAL_4 >= 4'h2;
  assign _EVAL_295 = _EVAL_7 == _EVAL_63;
  assign _EVAL_315 = _EVAL_28 | _EVAL_12;
  assign _EVAL_47 = ~_EVAL_240;
  assign _EVAL_171 = ~_EVAL_12;
  assign _EVAL_276 = _EVAL_54 | 2'h1;
  assign _EVAL_227 = ~_EVAL_280;
  assign _EVAL_131 = _EVAL_168 & _EVAL_203;
  assign _EVAL_44 = $signed(_EVAL_318) & -33'sh2000;
  assign _EVAL_45 = _EVAL_18 == 3'h6;
  assign _EVAL_34 = ~_EVAL_153;
  assign _EVAL_193 = _EVAL_110[31:0];
  assign _EVAL_254 = _EVAL_88 | _EVAL_12;
  assign _EVAL_239 = _EVAL_284;
  assign _EVAL_177 = _EVAL_15 ^ 32'h20000000;
  assign _EVAL_212 = _EVAL_120 | _EVAL_117;
  assign _EVAL_231 = ~_EVAL_241;
  assign _EVAL_167 = _EVAL_183 & _EVAL_203;
  assign _EVAL_170 = _EVAL_3 == _EVAL_66;
  assign _EVAL_169 = _EVAL_0 <= 4'h8;
  assign _EVAL_214 = _EVAL_7 & _EVAL_61;
  assign _EVAL_181 = _EVAL_9 & _EVAL_249;
  assign _EVAL_117 = _EVAL_188 ? _EVAL_37 : 2'h0;
  assign _EVAL_149 = ~_EVAL_55;
  assign _EVAL_87 = 23'hff << _EVAL_0;
  assign _EVAL_265 = _EVAL_223[5:0];
  assign _EVAL_264 = _EVAL_169 & _EVAL_50;
  assign _EVAL_179 = $signed(_EVAL_239) == 33'sh0;
  assign _EVAL_278 = _EVAL_89[7:2];
  assign _EVAL_48 = _EVAL_50 | _EVAL_104;
  assign _EVAL_28 = _EVAL_14 <= 2'h2;
  assign _EVAL_143 = _EVAL_39 >> _EVAL_13;
  assign _EVAL_49 = _EVAL_276[1];
  assign _EVAL_29 = _EVAL_11 & _EVAL_9;
  assign _EVAL_67 = ~_EVAL_273;
  assign _EVAL_244 = ~_EVAL_22;
  assign _EVAL_121 = _EVAL_71 == 6'h0;
  assign _EVAL_247 = _EVAL_85 | _EVAL_264;
  assign _EVAL_271 = _EVAL_0 >= 4'h2;
  assign _EVAL_89 = ~_EVAL_60;
  assign _EVAL_151 = _EVAL_120 != 2'h0;
  assign _EVAL_114 = _EVAL_138 & _EVAL_122;
  assign _EVAL_72 = ~_EVAL_209;
  assign _EVAL_109 = ~_EVAL_258;
  assign _EVAL_223 = _EVAL_282 - 6'h1;
  assign _EVAL_141 = {1'b0,$signed(_EVAL_140)};
  assign _EVAL_270 = ~_EVAL_164;
  assign _EVAL_50 = $signed(_EVAL_189) == 33'sh0;
  assign _EVAL_320 = _EVAL_6 & _EVAL_297;
  assign _EVAL_58 = _EVAL_277 | _EVAL_12;
  assign _EVAL_208 = _EVAL_120 >> _EVAL_2;
  assign _EVAL_137 = _EVAL_8 == 3'h6;
  assign _EVAL_103 = _EVAL_49 & _EVAL_168;
  assign _EVAL_138 = _EVAL_0 <= 4'h2;
  assign _EVAL_283 = _EVAL_86 | _EVAL_101;
  assign _EVAL_289 = _EVAL_201 | _EVAL_104;
  assign _EVAL_132 = 2'h1 << _EVAL_13;
  assign _EVAL_267 = ~_EVAL_70;
  assign _EVAL_246 = ~_EVAL_312;
  assign _EVAL_128 = _EVAL_305 | _EVAL_12;
  assign _EVAL_64 = ~_EVAL_83;
  assign _EVAL_33 = ~_EVAL_307;
  assign _EVAL_74 = $signed(_EVAL_135) & -33'shc000;
  assign _EVAL_225 = _EVAL_9 & _EVAL_184;
  assign _EVAL_240 = _EVAL_32 | _EVAL_12;
  assign _EVAL_259 = _EVAL_8 == 3'h4;
  assign _EVAL_73 = ~_EVAL_84;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_24 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_26 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_27 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_66 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_71 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_120 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_130 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_180 = _RAND_7[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_194 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_213 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_236 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_243 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_252 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_279 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_282 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_287 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_304 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_5) begin
    if (_EVAL_12) begin
      _EVAL_24 <= 32'h0;
    end else if (_EVAL_155) begin
      _EVAL_24 <= 32'h0;
    end else begin
      _EVAL_24 <= _EVAL_193;
    end
    if (_EVAL_301) begin
      _EVAL_26 <= _EVAL_2;
    end
    if (_EVAL_12) begin
      _EVAL_27 <= 6'h0;
    end else if (_EVAL_185) begin
      if (_EVAL_308) begin
        if (_EVAL_238) begin
          _EVAL_27 <= _EVAL_108;
        end else begin
          _EVAL_27 <= 6'h0;
        end
      end else begin
        _EVAL_27 <= _EVAL_123;
      end
    end
    if (_EVAL_301) begin
      _EVAL_66 <= _EVAL_3;
    end
    if (_EVAL_12) begin
      _EVAL_71 <= 6'h0;
    end else if (_EVAL_29) begin
      if (_EVAL_121) begin
        if (_EVAL_204) begin
          _EVAL_71 <= _EVAL_278;
        end else begin
          _EVAL_71 <= 6'h0;
        end
      end else begin
        _EVAL_71 <= _EVAL_261;
      end
    end
    if (_EVAL_12) begin
      _EVAL_120 <= 2'h0;
    end else begin
      _EVAL_120 <= _EVAL_285;
    end
    if (_EVAL_90) begin
      _EVAL_130 <= _EVAL_17;
    end
    if (_EVAL_12) begin
      _EVAL_180 <= 6'h0;
    end else if (_EVAL_185) begin
      if (_EVAL_230) begin
        if (_EVAL_238) begin
          _EVAL_180 <= _EVAL_108;
        end else begin
          _EVAL_180 <= 6'h0;
        end
      end else begin
        _EVAL_180 <= _EVAL_224;
      end
    end
    if (_EVAL_90) begin
      _EVAL_194 <= _EVAL_18;
    end
    if (_EVAL_301) begin
      _EVAL_213 <= _EVAL_8;
    end
    if (_EVAL_90) begin
      _EVAL_236 <= _EVAL_10;
    end
    if (_EVAL_90) begin
      _EVAL_243 <= _EVAL_4;
    end
    if (_EVAL_301) begin
      _EVAL_252 <= _EVAL_0;
    end
    if (_EVAL_301) begin
      _EVAL_279 <= _EVAL_15;
    end
    if (_EVAL_12) begin
      _EVAL_282 <= 6'h0;
    end else if (_EVAL_29) begin
      if (_EVAL_245) begin
        if (_EVAL_204) begin
          _EVAL_282 <= _EVAL_278;
        end else begin
          _EVAL_282 <= 6'h0;
        end
      end else begin
        _EVAL_282 <= _EVAL_265;
      end
    end
    if (_EVAL_90) begin
      _EVAL_287 <= _EVAL_14;
    end
    if (_EVAL_90) begin
      _EVAL_304 <= _EVAL_13;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afd189d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d50d3ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_303) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a2b1a9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cedbb2a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4a3ed6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_322) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a20aad11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(367ad8f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(532dfdd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_311) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3971dbe9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d909696)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_322) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d40214e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46589e9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47779b2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_310) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68b41c4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cea8e794)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fde0f62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95fc45ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5936f5cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93632caa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(193635c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adff85dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faf32356)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b851c92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_310) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62c6245)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(baaf203e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfcea3e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(108d6b68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95ec7fbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77031b21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3dde930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e836425e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b2559d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_299) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3e97ad3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9b9b984)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95f71f26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72f75509)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f96849e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(871837df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de9f22ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55f793fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74111759)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(700b6574)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_303) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a491891e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bbc0e4a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9925c76c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_311) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d754183f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f7927e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0fdd9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(939f55fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(274218bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_303) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e3e8422)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_311) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8474a01a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39675167)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_322) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38ba2189)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee89593e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb264eaa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(335dbdb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65a52e24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84cbd8e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94419b8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_311) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b387b855)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfee51f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4983bb91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ebd35bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b043aa43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f18b0eec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e557154)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d726ca7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_299) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd14be4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(952ac748)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0ef96d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97718c56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69a63f87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4e042e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_322) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e8f04c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6413ced3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a36777a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
