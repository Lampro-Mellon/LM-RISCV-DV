//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_85(
  input  [31:0] _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  output [2:0]  _EVAL_3,
  output        _EVAL_4,
  output        _EVAL_5,
  input  [29:0] _EVAL_6,
  output [2:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  output        _EVAL_10,
  output [31:0] _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input  [31:0] _EVAL_14,
  output        _EVAL_15,
  input  [3:0]  _EVAL_16,
  output [1:0]  _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19,
  input         _EVAL_20,
  input  [1:0]  _EVAL_21,
  output        _EVAL_22,
  input  [2:0]  _EVAL_23,
  input         _EVAL_24,
  output [31:0] _EVAL_25,
  input         _EVAL_26,
  output [29:0] _EVAL_27,
  output [1:0]  _EVAL_28,
  input         _EVAL_29,
  output [3:0]  _EVAL_30,
  output [2:0]  _EVAL_31,
  input         _EVAL_32,
  output [1:0]  _EVAL_33
);
  reg [29:0] _EVAL_34;
  reg [31:0] _RAND_0;
  wire  _EVAL_35;
  wire [30:0] _EVAL_36;
  wire  _EVAL_37;
  reg [2:0] _EVAL_38;
  reg [31:0] _RAND_1;
  wire  _EVAL_39;
  wire [1:0] _EVAL_40;
  reg  _EVAL_41;
  reg [31:0] _RAND_2;
  wire [2:0] _EVAL_43;
  reg [1:0] _EVAL_45;
  reg [31:0] _RAND_3;
  wire  _EVAL_46;
  reg [31:0] _EVAL_47;
  reg [31:0] _RAND_4;
  wire  _EVAL_48;
  wire [1:0] _EVAL_49;
  wire  _EVAL_51;
  reg  _EVAL_54;
  reg [31:0] _RAND_5;
  wire  _EVAL_55;
  wire [1:0] _EVAL_57;
  wire [30:0] _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_61;
  reg  _EVAL_62;
  reg [31:0] _RAND_6;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire [30:0] _EVAL_67;
  wire  _EVAL_68;
  reg [2:0] _EVAL_71;
  reg [31:0] _RAND_7;
  wire  _EVAL_72;
  wire [2:0] _EVAL_75;
  wire [1:0] _EVAL_77;
  reg  _EVAL_79;
  reg [31:0] _RAND_8;
  wire [29:0] _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  reg [2:0] _EVAL_87;
  reg [31:0] _RAND_9;
  wire  _EVAL_88;
  reg  _EVAL_89;
  reg [31:0] _RAND_10;
  wire [1:0] _EVAL_90;
  wire  _EVAL_92;
  wire  _EVAL_93;
  reg  _EVAL_94;
  reg [31:0] _RAND_11;
  wire  _EVAL_95;
  reg  _EVAL_96;
  reg [31:0] _RAND_12;
  wire  _EVAL_97;
  wire  Queue__EVAL;
  wire  Queue__EVAL_0;
  wire [31:0] Queue__EVAL_1;
  wire [31:0] Queue__EVAL_2;
  wire [1:0] Queue__EVAL_3;
  wire [2:0] Queue__EVAL_4;
  wire [2:0] Queue__EVAL_5;
  wire  Queue__EVAL_6;
  wire  Queue__EVAL_7;
  wire [2:0] Queue__EVAL_8;
  wire [2:0] Queue__EVAL_9;
  wire  Queue__EVAL_10;
  wire  Queue__EVAL_11;
  wire [1:0] Queue__EVAL_12;
  wire  Queue__EVAL_13;
  wire  Queue__EVAL_14;
  wire  Queue__EVAL_15;
  wire  Queue__EVAL_16;
  wire [1:0] Queue__EVAL_17;
  wire  Queue__EVAL_18;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  reg [1:0] _EVAL_104;
  reg [31:0] _RAND_13;
  reg [31:0] _EVAL_105;
  reg [31:0] _RAND_14;
  reg  _EVAL_106;
  reg [31:0] _RAND_15;
  wire  _EVAL_107;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_112;
  reg  _EVAL_113;
  reg [31:0] _RAND_16;
  wire  _EVAL_114;
  wire  _EVAL_116;
  wire  _EVAL_117;
  reg  _EVAL_118;
  reg [31:0] _RAND_17;
  wire [1:0] _EVAL_119;
  wire  _EVAL_124;
  reg [1:0] _EVAL_125;
  reg [31:0] _RAND_18;
  wire [1:0] _EVAL_126;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_134;
  wire  _EVAL_137;
  wire  _EVAL_139;
  wire  _EVAL_141;
  reg  _EVAL_142;
  reg [31:0] _RAND_19;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  _EVAL_84 Queue (
    ._EVAL(Queue__EVAL),
    ._EVAL_0(Queue__EVAL_0),
    ._EVAL_1(Queue__EVAL_1),
    ._EVAL_2(Queue__EVAL_2),
    ._EVAL_3(Queue__EVAL_3),
    ._EVAL_4(Queue__EVAL_4),
    ._EVAL_5(Queue__EVAL_5),
    ._EVAL_6(Queue__EVAL_6),
    ._EVAL_7(Queue__EVAL_7),
    ._EVAL_8(Queue__EVAL_8),
    ._EVAL_9(Queue__EVAL_9),
    ._EVAL_10(Queue__EVAL_10),
    ._EVAL_11(Queue__EVAL_11),
    ._EVAL_12(Queue__EVAL_12),
    ._EVAL_13(Queue__EVAL_13),
    ._EVAL_14(Queue__EVAL_14),
    ._EVAL_15(Queue__EVAL_15),
    ._EVAL_16(Queue__EVAL_16),
    ._EVAL_17(Queue__EVAL_17),
    ._EVAL_18(Queue__EVAL_18)
  );
  assign _EVAL_27 = _EVAL_34;
  assign _EVAL_116 = _EVAL_55 ? 1'h0 : _EVAL_46;
  assign _EVAL_134 = ~_EVAL_106;
  assign _EVAL_17 = Queue__EVAL_17;
  assign _EVAL_40 = {_EVAL_113,_EVAL_79};
  assign _EVAL_85 = _EVAL_55 | _EVAL_137;
  assign _EVAL_139 = ~_EVAL_142;
  assign _EVAL_25 = Queue__EVAL_1;
  assign _EVAL_75 = _EVAL_104 + _EVAL_119;
  assign _EVAL_3 = Queue__EVAL_5;
  assign _EVAL_55 = _EVAL_118 & _EVAL_93;
  assign _EVAL_130 = _EVAL_118 & _EVAL_112;
  assign _EVAL_59 = _EVAL_112 & _EVAL_118;
  assign _EVAL_100 = _EVAL_144 & _EVAL_131;
  assign _EVAL_97 = ~_EVAL_96;
  assign _EVAL_18 = Queue__EVAL_6;
  assign _EVAL_109 = _EVAL_2[2];
  assign _EVAL_117 = _EVAL_96 ? 1'h0 : 1'h1;
  assign Queue__EVAL_15 = _EVAL_20;
  assign Queue__EVAL_12 = _EVAL_125;
  assign _EVAL_95 = ~_EVAL_109;
  assign _EVAL_33 = _EVAL_98 ? 2'h2 : 2'h0;
  assign _EVAL_90 = _EVAL_75[1:0];
  assign _EVAL_67 = _EVAL_137 ? {{1'd0}, _EVAL_34} : _EVAL_58;
  assign _EVAL_46 = _EVAL_85 ? _EVAL_61 : _EVAL_124;
  assign Queue__EVAL_18 = _EVAL_29;
  assign _EVAL_36 = _EVAL_55 ? {{1'd0}, _EVAL_34} : _EVAL_67;
  assign _EVAL_43 = _EVAL_90 - _EVAL_57;
  assign _EVAL_57 = {{1'd0}, _EVAL_145};
  assign Queue__EVAL_4 = _EVAL_71;
  assign _EVAL_66 = _EVAL_144 & _EVAL_94;
  assign _EVAL_7 = _EVAL_87;
  assign _EVAL_77 = _EVAL_142 ? 2'h2 : {{1'd0}, _EVAL_117};
  assign _EVAL_49 = {_EVAL_41,_EVAL_88};
  assign _EVAL_5 = _EVAL_55 ? 1'h0 : _EVAL_48;
  assign Queue__EVAL_13 = _EVAL_106 & _EVAL_65;
  assign _EVAL_124 = _EVAL_37 & _EVAL_0;
  assign Queue__EVAL_7 = _EVAL_141 & _EVAL_139;
  assign _EVAL_37 = _EVAL_55 ? 1'h0 : _EVAL_48;
  assign _EVAL_15 = Queue__EVAL_10;
  assign _EVAL_112 = _EVAL_32 | _EVAL_68;
  assign _EVAL_58 = {{1'd0}, _EVAL_34};
  assign _EVAL_64 = _EVAL_2 == 3'h5;
  assign _EVAL_92 = ~_EVAL_118;
  assign _EVAL_99 = _EVAL_124 & _EVAL_35;
  assign _EVAL_4 = _EVAL_94;
  assign _EVAL_131 = _EVAL_72 | _EVAL_0;
  assign _EVAL_126 = _EVAL_43[1:0];
  assign _EVAL_144 = ~_EVAL_114;
  assign _EVAL_137 = _EVAL_89 & _EVAL_92;
  assign _EVAL_10 = Queue__EVAL_11;
  assign _EVAL_145 = _EVAL_20 & _EVAL_86;
  assign _EVAL_35 = ~_EVAL_64;
  assign _EVAL_141 = _EVAL_8 & _EVAL_96;
  assign _EVAL_93 = ~_EVAL_112;
  assign _EVAL_107 = ~_EVAL_54;
  assign _EVAL_39 = _EVAL_134 | _EVAL_142;
  assign _EVAL_98 = _EVAL_118 & _EVAL_107;
  assign _EVAL_28 = Queue__EVAL_3;
  assign _EVAL_84 = _EVAL_36[29:0];
  assign _EVAL_110 = _EVAL_8 & _EVAL_97;
  assign _EVAL_48 = _EVAL_85 ? _EVAL_66 : _EVAL_144;
  assign Queue__EVAL_2 = _EVAL;
  assign _EVAL_65 = _EVAL_32 | _EVAL_142;
  assign _EVAL_114 = _EVAL_104 >= 2'h3;
  assign _EVAL_11 = _EVAL_47;
  assign _EVAL_61 = _EVAL_144 & _EVAL_72;
  assign Queue__EVAL_14 = _EVAL_9;
  assign _EVAL_30 = {_EVAL_40,_EVAL_49};
  assign _EVAL_51 = _EVAL_124 | _EVAL_55;
  assign Queue__EVAL_9 = {{1'd0}, _EVAL_77};
  assign _EVAL_31 = Queue__EVAL_8;
  assign _EVAL_143 = _EVAL_124 | _EVAL_85;
  assign Queue__EVAL_16 = _EVAL_110 & _EVAL_139;
  assign _EVAL_22 = Queue__EVAL_0;
  assign _EVAL_72 = ~_EVAL_94;
  assign _EVAL_68 = _EVAL_54 & _EVAL_39;
  assign _EVAL_119 = {{1'd0}, _EVAL_116};
  assign _EVAL_88 = ~_EVAL_62;
  assign _EVAL_86 = Queue__EVAL_11;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_34 = _RAND_0[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_38 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_41 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_45 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_47 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_54 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_62 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_71 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_79 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_87 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_89 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_94 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_96 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_104 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_105 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_106 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_113 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_118 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_125 = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_142 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_9) begin
    if (_EVAL_29) begin
      _EVAL_34 <= 30'h0;
    end else if (_EVAL_55) begin
      _EVAL_34 <= _EVAL_84;
    end else if (_EVAL_85) begin
      _EVAL_34 <= _EVAL_84;
    end else if (_EVAL_99) begin
      _EVAL_34 <= _EVAL_6;
    end else begin
      _EVAL_34 <= _EVAL_84;
    end
    if (!(_EVAL_55)) begin
      if (!(_EVAL_85)) begin
        if (_EVAL_124) begin
          _EVAL_38 <= _EVAL_12;
        end
      end
    end
    if (!(_EVAL_55)) begin
      if (!(_EVAL_85)) begin
        if (_EVAL_124) begin
          _EVAL_41 <= _EVAL_26;
        end
      end
    end
    if (!(_EVAL_55)) begin
      if (!(_EVAL_85)) begin
        if (_EVAL_124) begin
          _EVAL_45 <= _EVAL_21;
        end
      end
    end
    if (_EVAL_112) begin
      _EVAL_47 <= _EVAL_105;
    end
    if (!(_EVAL_55)) begin
      if (!(_EVAL_85)) begin
        if (_EVAL_124) begin
          _EVAL_54 <= _EVAL_64;
        end
      end
    end
    if (!(_EVAL_55)) begin
      if (!(_EVAL_85)) begin
        if (_EVAL_124) begin
          _EVAL_62 <= _EVAL_24;
        end
      end
    end
    if (_EVAL_59) begin
      _EVAL_71 <= _EVAL_38;
    end
    if (!(_EVAL_55)) begin
      if (!(_EVAL_85)) begin
        if (_EVAL_124) begin
          _EVAL_79 <= _EVAL_19;
        end
      end
    end
    if (_EVAL_29) begin
      _EVAL_87 <= 3'h0;
    end else if (!(_EVAL_55)) begin
      if (!(_EVAL_85)) begin
        if (_EVAL_99) begin
          _EVAL_87 <= {{1'd0}, _EVAL_21};
        end
      end
    end
    if (_EVAL_29) begin
      _EVAL_89 <= 1'h0;
    end else if (_EVAL_55) begin
      _EVAL_89 <= _EVAL_85;
    end else if (_EVAL_85) begin
      _EVAL_89 <= _EVAL_85;
    end else begin
      _EVAL_89 <= _EVAL_143;
    end
    if (!(_EVAL_55)) begin
      if (!(_EVAL_85)) begin
        if (_EVAL_99) begin
          _EVAL_94 <= _EVAL_95;
        end
      end
    end
    if (_EVAL_59) begin
      _EVAL_96 <= _EVAL_94;
    end
    if (_EVAL_29) begin
      _EVAL_104 <= 2'h0;
    end else begin
      _EVAL_104 <= _EVAL_126;
    end
    if (!(_EVAL_55)) begin
      if (_EVAL_85) begin
        _EVAL_105 <= _EVAL_14;
      end else if (_EVAL_99) begin
        _EVAL_105 <= _EVAL_14;
      end
    end
    if (_EVAL_29) begin
      _EVAL_106 <= 1'h0;
    end else if (_EVAL_65) begin
      _EVAL_106 <= _EVAL_130;
    end
    if (!(_EVAL_55)) begin
      if (!(_EVAL_85)) begin
        if (_EVAL_124) begin
          _EVAL_113 <= _EVAL_13;
        end
      end
    end
    if (_EVAL_29) begin
      _EVAL_118 <= 1'h0;
    end else if (_EVAL_55) begin
      _EVAL_118 <= _EVAL_55;
    end else if (_EVAL_85) begin
      _EVAL_118 <= _EVAL_100;
    end else begin
      _EVAL_118 <= _EVAL_51;
    end
    if (_EVAL_59) begin
      _EVAL_125 <= _EVAL_45;
    end
    if (_EVAL_59) begin
      _EVAL_142 <= _EVAL_54;
    end
  end
endmodule
