//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_160(
  output        _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  output [3:0]  _EVAL_3,
  input         _EVAL_4,
  output        _EVAL_5,
  input         _EVAL_6,
  input  [31:0] _EVAL_7,
  input         _EVAL_8,
  output [1:0]  _EVAL_9,
  output [3:0]  _EVAL_10,
  input  [1:0]  _EVAL_11,
  output [31:0] _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  output        _EVAL_15,
  input         _EVAL_16,
  output        _EVAL_17,
  output        _EVAL_18,
  output [31:0] _EVAL_19,
  output        _EVAL_20,
  input  [3:0]  _EVAL_21,
  input  [3:0]  _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  output        _EVAL_25,
  output [2:0]  _EVAL_26,
  input         _EVAL_27,
  input  [2:0]  _EVAL_28,
  input  [3:0]  _EVAL_29,
  output [31:0] _EVAL_30,
  output        _EVAL_31,
  output        _EVAL_32,
  output        _EVAL_33,
  output [2:0]  _EVAL_34,
  output        _EVAL_35,
  input         _EVAL_36,
  input  [2:0]  _EVAL_37,
  input  [31:0] _EVAL_38,
  output        _EVAL_39,
  output        _EVAL_40,
  input         _EVAL_41,
  input         _EVAL_42,
  output        _EVAL_43,
  output [2:0]  _EVAL_44,
  input         _EVAL_45,
  output        _EVAL_46,
  input         _EVAL_47,
  output        _EVAL_48,
  input  [31:0] _EVAL_49,
  output        _EVAL_50,
  output [3:0]  _EVAL_51,
  input         _EVAL_52,
  input         _EVAL_53,
  input         _EVAL_54
);
  assign _EVAL_5 = _EVAL_47;
  assign _EVAL_26 = _EVAL_37;
  assign _EVAL_35 = _EVAL_36;
  assign _EVAL_43 = _EVAL_0;
  assign _EVAL_39 = _EVAL_4;
  assign _EVAL = _EVAL_52;
  assign _EVAL_9 = _EVAL_11;
  assign _EVAL_15 = _EVAL_45;
  assign _EVAL_33 = _EVAL_53;
  assign _EVAL_3 = _EVAL_21;
  assign _EVAL_46 = _EVAL_54;
  assign _EVAL_18 = _EVAL_24;
  assign _EVAL_20 = _EVAL_23;
  assign _EVAL_31 = _EVAL_16;
  assign _EVAL_50 = _EVAL_6;
  assign _EVAL_34 = _EVAL_28;
  assign _EVAL_17 = _EVAL_8;
  assign _EVAL_10 = _EVAL_22;
  assign _EVAL_19 = _EVAL_38;
  assign _EVAL_32 = _EVAL_41;
  assign _EVAL_44 = _EVAL_1;
  assign _EVAL_48 = _EVAL_13;
  assign _EVAL_30 = _EVAL_7;
  assign _EVAL_40 = _EVAL_14;
  assign _EVAL_12 = _EVAL_49;
  assign _EVAL_25 = _EVAL_42;
  assign _EVAL_51 = _EVAL_29;
endmodule
