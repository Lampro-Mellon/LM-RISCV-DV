//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_116(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  output [7:0]  _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19,
  input         _EVAL_20,
  input         _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  input  [2:0]  _EVAL_25,
  input  [1:0]  _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  input         _EVAL_38,
  input         _EVAL_39,
  input         _EVAL_40,
  input         _EVAL_41,
  input         _EVAL_42,
  input         _EVAL_43,
  input         _EVAL_44,
  input         _EVAL_45,
  input         _EVAL_46,
  output        _EVAL_47,
  input         _EVAL_48,
  output        _EVAL_49,
  input         _EVAL_50,
  input         _EVAL_51,
  input         _EVAL_52,
  input         _EVAL_53,
  input         _EVAL_54,
  input         _EVAL_55,
  input         _EVAL_56,
  input         _EVAL_57,
  input         _EVAL_58,
  input         _EVAL_59,
  input         _EVAL_60,
  input         _EVAL_61,
  input         _EVAL_62,
  input         _EVAL_63,
  input         _EVAL_64,
  input         _EVAL_65,
  input         _EVAL_66,
  output [31:0] _EVAL_67,
  output [2:0]  _EVAL_68,
  input         _EVAL_69,
  input         _EVAL_70,
  input         _EVAL_71,
  input         _EVAL_72,
  input         _EVAL_73,
  input         _EVAL_74,
  input         _EVAL_75,
  input         _EVAL_76,
  input  [2:0]  _EVAL_77,
  output        _EVAL_78,
  input         _EVAL_79,
  input         _EVAL_80,
  input         _EVAL_81,
  input         _EVAL_82,
  input         _EVAL_83,
  input         _EVAL_84,
  input         _EVAL_85,
  output [7:0]  _EVAL_86,
  input         _EVAL_87,
  input  [2:0]  _EVAL_88,
  input         _EVAL_89,
  input         _EVAL_90,
  input         _EVAL_91,
  input         _EVAL_92,
  input         _EVAL_93,
  input         _EVAL_94,
  input         _EVAL_95,
  input         _EVAL_96,
  input         _EVAL_97,
  input         _EVAL_98,
  input         _EVAL_99,
  input         _EVAL_100,
  input         _EVAL_101,
  input         _EVAL_102,
  input         _EVAL_103,
  input         _EVAL_104,
  input         _EVAL_105,
  input         _EVAL_106,
  input         _EVAL_107,
  input         _EVAL_108,
  input         _EVAL_109,
  input         _EVAL_110,
  input         _EVAL_111,
  input         _EVAL_112,
  output        _EVAL_113,
  input         _EVAL_114,
  input         _EVAL_115,
  input         _EVAL_116,
  input         _EVAL_117,
  input         _EVAL_118,
  input         _EVAL_119,
  output [1:0]  _EVAL_120,
  input         _EVAL_121,
  input         _EVAL_122,
  input         _EVAL_123,
  input  [3:0]  _EVAL_124,
  input         _EVAL_125,
  input         _EVAL_126,
  input         _EVAL_127,
  input         _EVAL_128,
  input         _EVAL_129,
  input         _EVAL_130,
  input  [25:0] _EVAL_131,
  input         _EVAL_132,
  input         _EVAL_133,
  input         _EVAL_134,
  input         _EVAL_135,
  input         _EVAL_136,
  input         _EVAL_137,
  output [2:0]  _EVAL_138,
  input         _EVAL_139,
  input  [31:0] _EVAL_140,
  input         _EVAL_141,
  output        _EVAL_142,
  input         _EVAL_143,
  input         _EVAL_144,
  output        _EVAL_145,
  input         _EVAL_146,
  input         _EVAL_147,
  input         _EVAL_148,
  input         _EVAL_149,
  input         _EVAL_150,
  input         _EVAL_151,
  input         _EVAL_152,
  input         _EVAL_153
);
  wire  _EVAL_156;
  wire  _EVAL_158;
  wire  _EVAL_160;
  wire [25:0] _EVAL_161;
  wire  _EVAL_163;
  reg [3:0] _EVAL_164;
  reg [31:0] _RAND_0;
  wire [7:0] _EVAL_165;
  wire [7:0] _EVAL_166;
  wire [1:0] _EVAL_167;
  wire [1:0] _EVAL_170;
  wire [31:0] _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_176;
  wire [7:0] _EVAL_178;
  wire [17:0] _EVAL_180;
  wire [15:0] _EVAL_182;
  wire  _EVAL_185;
  wire [9:0] _EVAL_186;
  wire [15:0] _EVAL_188;
  wire [4:0] _EVAL_189;
  wire [31:0] _EVAL_190;
  wire [4:0] _EVAL_192;
  wire  _EVAL_195;
  wire  _EVAL_197;
  wire [4:0] _EVAL_198;
  wire [7:0] _EVAL_199;
  wire  _EVAL_203;
  wire [23:0] _EVAL_211;
  reg  _EVAL_212;
  reg [31:0] _RAND_1;
  wire  _EVAL_215;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire [4:0] _EVAL_220;
  wire  _EVAL_226;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire [9:0] _EVAL_232;
  wire  _EVAL_234;
  reg  _EVAL_236;
  reg [31:0] _RAND_2;
  wire [4:0] _EVAL_238;
  wire [15:0] _EVAL_240;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire [25:0] _EVAL_250;
  wire [31:0] _EVAL_255;
  wire [31:0] _EVAL_261;
  wire [25:0] _EVAL_264;
  wire  _EVAL_267;
  wire  _EVAL_270;
  reg [3:0] _EVAL_272;
  reg [31:0] _RAND_3;
  wire [17:0] _EVAL_273;
  wire [2:0] _EVAL_274;
  wire [4:0] _EVAL_276;
  reg  _EVAL_277;
  reg [31:0] _RAND_4;
  wire  _EVAL_278;
  wire  _EVAL_281;
  wire  _EVAL_283;
  wire [4:0] _EVAL_285;
  wire [9:0] _EVAL_286;
  wire [23:0] _EVAL_288;
  wire  _EVAL_289;
  wire [15:0] _EVAL_291;
  wire [1:0] _EVAL_293;
  wire [31:0] _EVAL_294;
  wire [4:0] _EVAL_295;
  reg [3:0] _EVAL_296;
  reg [31:0] _RAND_5;
  wire  _EVAL_297;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire [25:0] _EVAL_304;
  wire [3:0] _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_308;
  wire  _EVAL_311;
  wire [9:0] _EVAL_312;
  wire [31:0] _EVAL_313;
  wire  _EVAL_315;
  wire  _EVAL_317;
  wire  _EVAL_320;
  wire [7:0] _EVAL_324;
  wire [21:0] _EVAL_325;
  wire [4:0] _EVAL_329;
  wire  _EVAL_333;
  wire  _EVAL_336;
  wire [17:0] _EVAL_337;
  wire  _EVAL_338;
  wire  _EVAL_340;
  wire  _EVAL_343;
  wire [23:0] _EVAL_344;
  wire [4:0] _EVAL_349;
  wire [7:0] _EVAL_350;
  wire  _EVAL_353;
  reg  _EVAL_355;
  reg [31:0] _RAND_6;
  reg  _EVAL_356;
  reg [31:0] _RAND_7;
  wire  _EVAL_359;
  wire [15:0] _EVAL_366;
  wire  _EVAL_367;
  wire [4:0] _EVAL_368;
  wire [31:0] _EVAL_371;
  wire [15:0] _EVAL_379;
  reg  _EVAL_381;
  reg [31:0] _RAND_8;
  wire [15:0] _EVAL_382;
  wire  _EVAL_384;
  wire  _EVAL_393;
  wire [7:0] _EVAL_394;
  wire  _EVAL_397;
  wire [15:0] _EVAL_399;
  wire [1:0] _EVAL_400;
  wire [31:0] _EVAL_401;
  wire [31:0] _EVAL_403;
  reg [7:0] _EVAL_404;
  reg [31:0] _RAND_9;
  wire [4:0] _EVAL_405;
  wire  _EVAL_406;
  wire [7:0] _EVAL_411;
  reg [3:0] _EVAL_412;
  reg [31:0] _RAND_10;
  wire [31:0] _EVAL_414;
  wire [31:0] _EVAL_416;
  wire  _EVAL_417;
  wire [1:0] _EVAL_419;
  wire [2:0] _EVAL_420;
  wire  _EVAL_423;
  wire [2:0] _EVAL_425;
  wire [1:0] _EVAL_426;
  wire  _EVAL_427;
  wire [4:0] _EVAL_430;
  wire [4:0] _EVAL_431;
  wire  _EVAL_432;
  wire  _EVAL_433;
  wire [9:0] _EVAL_436;
  wire [9:0] _EVAL_437;
  wire [31:0] _EVAL_438;
  wire [31:0] _EVAL_439;
  wire [25:0] _EVAL_443;
  wire  _EVAL_444;
  wire [4:0] _EVAL_445;
  wire [25:0] _EVAL_447;
  wire [2:0] _EVAL_448;
  wire [17:0] _EVAL_450;
  wire [1:0] _EVAL_452;
  reg  _EVAL_454;
  reg [31:0] _RAND_11;
  wire  _EVAL_455;
  wire [4:0] _EVAL_459;
  wire  _EVAL_463;
  wire  _EVAL_465;
  wire [4:0] _EVAL_466;
  wire  _EVAL_468;
  wire  _EVAL_471;
  wire  _EVAL_472;
  wire [4:0] _EVAL_483;
  reg  _EVAL_484;
  reg [31:0] _RAND_12;
  wire  _EVAL_485;
  reg  _EVAL_487;
  reg [31:0] _RAND_13;
  wire  _EVAL_488;
  wire  _EVAL_489;
  reg [3:0] _EVAL_493;
  reg [31:0] _RAND_14;
  wire [31:0] _EVAL_494;
  wire [4:0] _EVAL_495;
  wire [23:0] _EVAL_497;
  wire [31:0] _EVAL_498;
  wire [17:0] _EVAL_499;
  wire  _EVAL_500;
  wire  _EVAL_501;
  wire [1:0] _EVAL_502;
  wire [23:0] _EVAL_505;
  reg  _EVAL_506;
  reg [31:0] _RAND_15;
  reg  _EVAL_507;
  reg [31:0] _RAND_16;
  wire  _EVAL_511;
  wire [7:0] _EVAL_514;
  wire  _EVAL_516;
  wire  _EVAL_517;
  wire [31:0] _EVAL_518;
  wire  _EVAL_519;
  wire  _EVAL_520;
  wire [1:0] _EVAL_522;
  wire  _EVAL_524;
  wire [15:0] _EVAL_525;
  wire [15:0] _EVAL_526;
  wire  _EVAL_527;
  reg [3:0] _EVAL_531;
  reg [31:0] _RAND_17;
  wire  _EVAL_533;
  reg [3:0] _EVAL_542;
  reg [31:0] _RAND_18;
  wire  _EVAL_543;
  wire [7:0] _EVAL_545;
  reg  _EVAL_546;
  reg [31:0] _RAND_19;
  wire  _EVAL_547;
  wire [2:0] _EVAL_548;
  wire  _EVAL_550;
  wire  _EVAL_553;
  wire  _EVAL_556;
  wire  _EVAL_557;
  reg [3:0] _EVAL_558;
  reg [31:0] _RAND_20;
  wire  _EVAL_559;
  reg  _EVAL_560;
  reg [31:0] _RAND_21;
  reg [3:0] _EVAL_561;
  reg [31:0] _RAND_22;
  reg [3:0] _EVAL_563;
  reg [31:0] _RAND_23;
  wire [31:0] _EVAL_567;
  wire [4:0] _EVAL_569;
  wire  _EVAL_571;
  wire [7:0] _EVAL_575;
  wire  _EVAL_576;
  reg  _EVAL_582;
  reg [31:0] _RAND_24;
  wire [1:0] _EVAL_592;
  wire [23:0] _EVAL_593;
  wire  _EVAL_595;
  wire  _EVAL_597;
  wire [17:0] _EVAL_598;
  wire  _EVAL_601;
  wire [4:0] _EVAL_602;
  reg  _EVAL_603;
  reg [31:0] _RAND_25;
  wire [4:0] _EVAL_604;
  wire [23:0] _EVAL_605;
  wire  _EVAL_606;
  reg [3:0] _EVAL_607;
  reg [31:0] _RAND_26;
  wire [31:0] _EVAL_609;
  wire  _EVAL_611;
  wire [7:0] _EVAL_614;
  wire  _EVAL_615;
  reg  _EVAL_616;
  reg [31:0] _RAND_27;
  wire  _EVAL_618;
  wire  _EVAL_624;
  wire  _EVAL_628;
  wire [4:0] _EVAL_632;
  wire [4:0] _EVAL_634;
  wire  _EVAL_636;
  wire [9:0] _EVAL_639;
  wire  _EVAL_640;
  wire [4:0] _EVAL_642;
  reg  _EVAL_643;
  reg [31:0] _RAND_28;
  reg  _EVAL_644;
  reg [31:0] _RAND_29;
  wire [4:0] _EVAL_647;
  wire [1:0] _EVAL_648;
  wire  _EVAL_650;
  reg [3:0] _EVAL_653;
  reg [31:0] _RAND_30;
  wire [1:0] _EVAL_655;
  wire [9:0] _EVAL_657;
  wire  _EVAL_658;
  reg  _EVAL_661;
  reg [31:0] _RAND_31;
  wire [7:0] _EVAL_662;
  wire [4:0] _EVAL_664;
  wire [31:0] _EVAL_665;
  reg  _EVAL_666;
  reg [31:0] _RAND_32;
  wire [9:0] _EVAL_667;
  wire  _EVAL_669;
  wire  _EVAL_671;
  wire [4:0] _EVAL_672;
  wire  _EVAL_673;
  wire [4:0] _EVAL_674;
  wire  _EVAL_675;
  wire  _EVAL_676;
  wire [17:0] _EVAL_677;
  wire  _EVAL_678;
  wire [7:0] _EVAL_681;
  wire [25:0] _EVAL_683;
  wire [4:0] _EVAL_685;
  wire [4:0] _EVAL_687;
  wire  _EVAL_689;
  reg  _EVAL_690;
  reg [31:0] _RAND_33;
  wire  _EVAL_691;
  wire [9:0] _EVAL_693;
  wire  _EVAL_696;
  wire  _EVAL_697;
  wire [4:0] _EVAL_700;
  reg [3:0] _EVAL_702;
  reg [31:0] _RAND_34;
  reg [3:0] _EVAL_703;
  reg [31:0] _RAND_35;
  wire [31:0] _EVAL_705;
  wire [1:0] _EVAL_706;
  wire [31:0] _EVAL_707;
  wire [31:0] _EVAL_715;
  wire [23:0] _EVAL_716;
  wire [23:0] _EVAL_717;
  wire [31:0] _EVAL_718;
  wire [7:0] _EVAL_719;
  wire [4:0] _EVAL_720;
  wire  _EVAL_723;
  wire  _EVAL_724;
  reg  _EVAL_727;
  reg [31:0] _RAND_36;
  wire [1:0] _EVAL_728;
  wire [4:0] _EVAL_729;
  wire [4:0] _EVAL_730;
  wire [31:0] _EVAL_732;
  wire [4:0] _EVAL_733;
  wire [2:0] _EVAL_736;
  reg [3:0] _EVAL_737;
  reg [31:0] _RAND_37;
  wire [25:0] _EVAL_738;
  wire [23:0] _EVAL_741;
  wire  _EVAL_742;
  wire [4:0] _EVAL_743;
  wire  _EVAL_747;
  wire [1:0] _EVAL_749;
  wire [9:0] _EVAL_750;
  wire [7:0] _EVAL_753;
  wire  _EVAL_756;
  wire  _EVAL_759;
  wire  _EVAL_760;
  wire  _EVAL_762;
  wire [4:0] _EVAL_763;
  wire  _EVAL_765;
  wire [1:0] _EVAL_766;
  wire [4:0] _EVAL_772;
  reg [3:0] _EVAL_780;
  reg [31:0] _RAND_38;
  wire  _EVAL_782;
  reg  _EVAL_783;
  reg [31:0] _RAND_39;
  wire [31:0] _EVAL_784;
  wire  _EVAL_785;
  wire  _EVAL_786;
  wire  _EVAL_788;
  wire  _EVAL_791;
  wire [9:0] _EVAL_794;
  wire  _EVAL_795;
  wire  _EVAL_796;
  wire [3:0] _EVAL_805;
  wire [31:0] _EVAL_806;
  wire  _EVAL_810;
  wire [9:0] _EVAL_811;
  wire  _EVAL_812;
  wire  _EVAL_813;
  wire [23:0] _EVAL_815;
  wire  _EVAL_822;
  wire  _EVAL_823;
  wire  _EVAL_824;
  wire [23:0] _EVAL_833;
  reg [3:0] _EVAL_834;
  reg [31:0] _RAND_40;
  wire  _EVAL_835;
  wire [23:0] _EVAL_838;
  wire [1:0] _EVAL_840;
  wire  _EVAL_841;
  wire  _EVAL_844;
  wire  _EVAL_846;
  wire  _EVAL_847;
  wire [7:0] _EVAL_848;
  wire  _EVAL_850;
  wire [7:0] _EVAL_851;
  wire [2:0] _EVAL_852;
  wire [4:0] _EVAL_853;
  wire  _EVAL_855;
  wire [4:0] _EVAL_858;
  reg [3:0] _EVAL_861;
  reg [31:0] _RAND_41;
  wire [4:0] _EVAL_863;
  wire  _EVAL_864;
  wire [31:0] _EVAL_866;
  wire [4:0] _EVAL_872;
  wire  _EVAL_874;
  wire  _EVAL_879;
  reg  _EVAL_880;
  reg [31:0] _RAND_42;
  wire  _EVAL_881;
  wire [4:0] _EVAL_883;
  reg  _EVAL_887;
  reg [31:0] _RAND_43;
  wire  _EVAL_889;
  wire [1:0] _EVAL_890;
  reg  _EVAL_891;
  reg [31:0] _RAND_44;
  wire  _EVAL_892;
  wire  _EVAL_893;
  reg  _EVAL_896;
  reg [31:0] _RAND_45;
  wire  _EVAL_898;
  reg [3:0] _EVAL_899;
  reg [31:0] _RAND_46;
  wire [4:0] _EVAL_901;
  wire [3:0] _EVAL_902;
  wire [4:0] _EVAL_903;
  reg  _EVAL_906;
  reg [31:0] _RAND_47;
  wire  _EVAL_907;
  wire  _EVAL_912;
  wire  _EVAL_913;
  wire [31:0] _EVAL_915;
  wire  _EVAL_916;
  wire [9:0] _EVAL_918;
  wire [4:0] _EVAL_919;
  wire  _EVAL_923;
  wire [17:0] _EVAL_924;
  wire [31:0] _EVAL_929;
  wire  _EVAL_930;
  wire  _EVAL_934;
  wire  _EVAL_939;
  wire  _EVAL_942;
  reg  _EVAL_943;
  reg [31:0] _RAND_48;
  wire  _EVAL_945;
  wire  _EVAL_948;
  wire [31:0] _EVAL_953;
  wire [31:0] _EVAL_958;
  wire [31:0] _EVAL_959;
  wire  _EVAL_960;
  wire [17:0] _EVAL_962;
  wire [15:0] _EVAL_966;
  wire  _EVAL_968;
  wire [3:0] _EVAL_969;
  wire  _EVAL_970;
  wire [15:0] _EVAL_977;
  wire  _EVAL_978;
  wire [9:0] _EVAL_979;
  wire [31:0] _EVAL_980;
  wire [31:0] _EVAL_981;
  wire [31:0] _EVAL_986;
  wire  _EVAL_988;
  wire [3:0] _EVAL_990;
  wire [25:0] _EVAL_991;
  wire  _EVAL_992;
  wire [1:0] _EVAL_993;
  reg [3:0] _EVAL_994;
  reg [31:0] _RAND_49;
  wire [4:0] _EVAL_995;
  wire [9:0] _EVAL_999;
  wire  _EVAL_1002;
  wire  _EVAL_1005;
  wire [7:0] _EVAL_1011;
  wire [23:0] _EVAL_1013;
  wire  _EVAL_1018;
  wire  _EVAL_1020;
  wire [2:0] _EVAL_1021;
  wire [4:0] _EVAL_1023;
  wire  _EVAL_1024;
  wire [7:0] _EVAL_1026;
  reg [3:0] _EVAL_1028;
  reg [31:0] _RAND_50;
  wire  _EVAL_1030;
  wire  _EVAL_1031;
  wire  _EVAL_1032;
  wire [7:0] _EVAL_1035;
  reg  _EVAL_1040;
  reg [31:0] _RAND_51;
  reg  _EVAL_1041;
  reg [31:0] _RAND_52;
  wire  _EVAL_1042;
  wire [15:0] _EVAL_1048;
  reg [3:0] _EVAL_1052;
  reg [31:0] _RAND_53;
  wire  _EVAL_1054;
  wire [9:0] _EVAL_1056;
  reg  _EVAL_1057;
  reg [31:0] _RAND_54;
  wire [31:0] Queue__EVAL;
  wire [2:0] Queue__EVAL_0;
  wire [2:0] Queue__EVAL_1;
  wire  Queue__EVAL_2;
  wire  Queue__EVAL_3;
  wire [3:0] Queue__EVAL_4;
  wire [3:0] Queue__EVAL_5;
  wire  Queue__EVAL_6;
  wire  Queue__EVAL_7;
  wire [21:0] Queue__EVAL_8;
  wire  Queue__EVAL_9;
  wire  Queue__EVAL_10;
  wire [1:0] Queue__EVAL_11;
  wire [1:0] Queue__EVAL_12;
  wire  Queue__EVAL_13;
  wire  Queue__EVAL_14;
  wire [31:0] Queue__EVAL_15;
  wire [21:0] Queue__EVAL_16;
  wire  _EVAL_1059;
  wire [25:0] _EVAL_1060;
  wire  _EVAL_1066;
  wire  _EVAL_1072;
  wire  _EVAL_1073;
  wire [4:0] _EVAL_1074;
  wire  _EVAL_1075;
  wire [7:0] _EVAL_1080;
  wire  _EVAL_1087;
  wire  _EVAL_1089;
  wire [7:0] _EVAL_1091;
  wire [14:0] _EVAL_1092;
  wire  _EVAL_1093;
  wire  _EVAL_1098;
  wire  _EVAL_1100;
  wire [7:0] _EVAL_1101;
  wire [7:0] _EVAL_1106;
  wire [25:0] _EVAL_1110;
  wire  _EVAL_1111;
  wire  _EVAL_1112;
  wire [9:0] _EVAL_1113;
  wire [4:0] _EVAL_1114;
  wire  _EVAL_1115;
  wire  _EVAL_1117;
  wire [4:0] _EVAL_1119;
  wire [4:0] _EVAL_1120;
  reg  _EVAL_1121;
  reg [31:0] _RAND_55;
  wire [3:0] _EVAL_1123;
  wire [1:0] _EVAL_1124;
  wire [1:0] _EVAL_1128;
  wire [2:0] _EVAL_1129;
  wire [1:0] _EVAL_1130;
  reg  _EVAL_1131;
  reg [31:0] _RAND_56;
  wire  _EVAL_1132;
  wire  _EVAL_1135;
  wire  _EVAL_1138;
  wire  _EVAL_1140;
  wire [1:0] _EVAL_1141;
  wire [7:0] _EVAL_1143;
  reg  _EVAL_1147;
  reg [31:0] _RAND_57;
  wire  _EVAL_1148;
  wire  _EVAL_1150;
  wire  _EVAL_1153;
  wire  _EVAL_1154;
  wire  _EVAL_1156;
  wire [6:0] _EVAL_1157;
  wire [31:0] _EVAL_1159;
  wire [31:0] _EVAL_1160;
  wire  _EVAL_1163;
  wire [1:0] _EVAL_1164;
  reg  _EVAL_1166;
  reg [31:0] _RAND_58;
  wire  _EVAL_1168;
  wire [9:0] _EVAL_1172;
  wire [2:0] _EVAL_1174;
  wire [17:0] _EVAL_1177;
  wire  _EVAL_1178;
  wire [1:0] _EVAL_1181;
  wire [3:0] _EVAL_1184;
  reg [3:0] _EVAL_1186;
  reg [31:0] _RAND_59;
  reg  _EVAL_1187;
  reg [31:0] _RAND_60;
  reg  _EVAL_1188;
  reg [31:0] _RAND_61;
  wire [7:0] _EVAL_1190;
  wire  _EVAL_1191;
  wire [7:0] _EVAL_1192;
  wire  _EVAL_1200;
  wire [15:0] _EVAL_1204;
  wire [9:0] _EVAL_1205;
  reg  _EVAL_1206;
  reg [31:0] _RAND_62;
  wire [7:0] _EVAL_1208;
  reg  _EVAL_1211;
  reg [31:0] _RAND_63;
  wire  _EVAL_1215;
  wire [4:0] _EVAL_1216;
  wire  _EVAL_1217;
  wire  _EVAL_1218;
  wire  _EVAL_1219;
  wire [31:0] _EVAL_1220;
  wire [4:0] _EVAL_1221;
  wire [1:0] _EVAL_1222;
  wire  _EVAL_1225;
  wire  _EVAL_1228;
  reg  _EVAL_1229;
  reg [31:0] _RAND_64;
  wire [2:0] _EVAL_1230;
  wire [7:0] _EVAL_1232;
  reg  _EVAL_1235;
  reg [31:0] _RAND_65;
  wire  _EVAL_1236;
  wire  _EVAL_1237;
  wire [7:0] _EVAL_1238;
  wire [17:0] _EVAL_1239;
  reg  _EVAL_1240;
  reg [31:0] _RAND_66;
  reg  _EVAL_1245;
  reg [31:0] _RAND_67;
  wire  _EVAL_1247;
  wire  _EVAL_1248;
  wire [31:0] _EVAL_1249;
  wire  _EVAL_1250;
  wire  _EVAL_1251;
  wire  _EVAL_1252;
  wire [1:0] _EVAL_1253;
  wire  _EVAL_1255;
  wire  _EVAL_1257;
  wire [17:0] _EVAL_1258;
  wire [3:0] _EVAL_1260;
  wire  _EVAL_1261;
  wire [17:0] _EVAL_1263;
  wire [1:0] _EVAL_1264;
  wire [1:0] _EVAL_1265;
  wire [23:0] _EVAL_1267;
  wire [3:0] _EVAL_1271;
  reg [3:0] _EVAL_1273;
  reg [31:0] _RAND_68;
  wire [2:0] _EVAL_1275;
  wire [9:0] _EVAL_1276;
  wire  _EVAL_1278;
  wire [31:0] _EVAL_1279;
  wire [11:0] _EVAL_1280;
  wire [7:0] _EVAL_1282;
  wire [4:0] _EVAL_1284;
  reg [7:0] _EVAL_1286;
  reg [31:0] _RAND_69;
  reg  _EVAL_1287;
  reg [31:0] _RAND_70;
  reg [3:0] _EVAL_1288;
  reg [31:0] _RAND_71;
  reg [3:0] _EVAL_1289;
  reg [31:0] _RAND_72;
  wire  _EVAL_1292;
  reg  _EVAL_1293;
  reg [31:0] _RAND_73;
  wire [7:0] _EVAL_1295;
  wire [3:0] _EVAL_1298;
  reg  _EVAL_1301;
  reg [31:0] _RAND_74;
  wire [1:0] _EVAL_1303;
  wire [2:0] _EVAL_1304;
  wire [1:0] _EVAL_1306;
  wire  _EVAL_1307;
  wire [31:0] _EVAL_1308;
  wire  _EVAL_1309;
  reg  _EVAL_1311;
  reg [31:0] _RAND_75;
  reg  _EVAL_1314;
  reg [31:0] _RAND_76;
  wire [31:0] _EVAL_1315;
  reg [3:0] _EVAL_1318;
  reg [31:0] _RAND_77;
  wire  _EVAL_1320;
  wire  _EVAL_1321;
  wire  _EVAL_1323;
  wire  _EVAL_1325;
  wire [1:0] _EVAL_1330;
  reg  _EVAL_1331;
  reg [31:0] _RAND_78;
  wire  _EVAL_1333;
  wire [31:0] _EVAL_1335;
  wire [4:0] _EVAL_1336;
  wire [4:0] _EVAL_1337;
  wire [4:0] _EVAL_1339;
  reg  _EVAL_1342;
  reg [31:0] _RAND_79;
  wire [7:0] _EVAL_1345;
  wire  _EVAL_1347;
  reg [3:0] _EVAL_1351;
  reg [31:0] _RAND_80;
  wire  _EVAL_1352;
  wire [1:0] _EVAL_1353;
  wire [4:0] _EVAL_1354;
  reg [3:0] _EVAL_1356;
  reg [31:0] _RAND_81;
  wire [1:0] _EVAL_1357;
  wire [4:0] _EVAL_1359;
  wire [9:0] _EVAL_1362;
  wire  _EVAL_1367;
  wire [31:0] _EVAL_1368;
  wire [31:0] _EVAL_1372;
  wire  _EVAL_1374;
  wire  _EVAL_1377;
  wire  _EVAL_1378;
  wire [25:0] _EVAL_1379;
  wire  _EVAL_1381;
  wire  _EVAL_1382;
  reg  _EVAL_1383;
  reg [31:0] _RAND_82;
  reg  _EVAL_1388;
  reg [31:0] _RAND_83;
  wire [1:0] _EVAL_1390;
  reg  _EVAL_1396;
  reg [31:0] _RAND_84;
  wire [3:0] _EVAL_1397;
  wire [23:0] _EVAL_1398;
  wire [31:0] _EVAL_1400;
  wire  _EVAL_1403;
  reg  _EVAL_1407;
  reg [31:0] _RAND_85;
  reg  _EVAL_1408;
  reg [31:0] _RAND_86;
  wire  _EVAL_1409;
  wire  _EVAL_1410;
  wire [4:0] _EVAL_1414;
  wire  _EVAL_1415;
  wire [1:0] _EVAL_1416;
  wire [3:0] _EVAL_1417;
  wire [31:0] _EVAL_1422;
  wire  _EVAL_1423;
  wire [31:0] _EVAL_1425;
  reg [3:0] _EVAL_1427;
  reg [31:0] _RAND_87;
  wire [1:0] _EVAL_1429;
  wire  _EVAL_1430;
  wire  _EVAL_1431;
  wire [3:0] _EVAL_1433;
  wire [31:0] _EVAL_1435;
  wire  _EVAL_1436;
  wire  _EVAL_1437;
  wire  _EVAL_1438;
  reg [3:0] _EVAL_1440;
  reg [31:0] _RAND_88;
  wire [4:0] _EVAL_1441;
  reg [3:0] _EVAL_1442;
  reg [31:0] _RAND_89;
  wire  _EVAL_1444;
  wire [25:0] _EVAL_1445;
  wire  _EVAL_1451;
  wire  _EVAL_1454;
  wire [7:0] _EVAL_1456;
  wire [4:0] _EVAL_1457;
  wire [1:0] _EVAL_1460;
  wire [15:0] _EVAL_1461;
  wire  _EVAL_1462;
  wire  _EVAL_1464;
  wire  _EVAL_1465;
  wire [23:0] _EVAL_1466;
  wire [4:0] _EVAL_1469;
  wire [4:0] _EVAL_1472;
  wire [15:0] _EVAL_1473;
  wire [4:0] _EVAL_1474;
  wire  _EVAL_1476;
  wire  _EVAL_1477;
  wire [17:0] _EVAL_1481;
  reg [3:0] _EVAL_1484;
  reg [31:0] _RAND_90;
  wire  _EVAL_1486;
  wire  _EVAL_1492;
  reg  _EVAL_1493;
  reg [31:0] _RAND_91;
  wire [5:0] _EVAL_1495;
  wire [1:0] _EVAL_1496;
  wire [7:0] _EVAL_1497;
  wire  _EVAL_1498;
  wire  _EVAL_1502;
  wire [31:0] _EVAL_1503;
  wire [4:0] _EVAL_1504;
  reg  _EVAL_1506;
  reg [31:0] _RAND_92;
  wire  _EVAL_1507;
  wire [5:0] _EVAL_1508;
  reg  _EVAL_1510;
  reg [31:0] _RAND_93;
  reg [3:0] _EVAL_1515;
  reg [31:0] _RAND_94;
  wire [4:0] _EVAL_1517;
  wire [15:0] _EVAL_1519;
  wire [4:0] _EVAL_1520;
  wire [15:0] _EVAL_1522;
  wire  _EVAL_1524;
  wire [15:0] _EVAL_1527;
  wire  _EVAL_1531;
  wire  _EVAL_1532;
  wire [4:0] _EVAL_1534;
  wire  _EVAL_1537;
  wire [31:0] _EVAL_1540;
  reg  _EVAL_1544;
  reg [31:0] _RAND_95;
  wire [23:0] _EVAL_1549;
  wire [31:0] _EVAL_1550;
  wire  _EVAL_1551;
  wire [17:0] _EVAL_1552;
  wire  _EVAL_1554;
  wire [17:0] _EVAL_1556;
  wire [4:0] _EVAL_1560;
  wire [15:0] _EVAL_1564;
  wire  _EVAL_1565;
  wire [4:0] _EVAL_1566;
  wire  _EVAL_1569;
  wire [4:0] _EVAL_1571;
  wire [31:0] _EVAL_1572;
  wire [23:0] _EVAL_1573;
  wire  _EVAL_1575;
  wire [4:0] _EVAL_1576;
  wire [4:0] _EVAL_1577;
  reg  _EVAL_1581;
  reg [31:0] _RAND_96;
  wire [2:0] _EVAL_1583;
  wire [11:0] _EVAL_1587;
  wire  _EVAL_1589;
  wire  _EVAL_1592;
  reg  _EVAL_1593;
  reg [31:0] _RAND_97;
  wire  _EVAL_1595;
  wire [15:0] _EVAL_1597;
  wire  _EVAL_1598;
  reg  _EVAL_1602;
  reg [31:0] _RAND_98;
  wire  _EVAL_1608;
  wire [4:0] _EVAL_1609;
  reg [3:0] _EVAL_1610;
  reg [31:0] _RAND_99;
  wire  _EVAL_1613;
  wire  _EVAL_1614;
  wire [31:0] _EVAL_1617;
  reg  _EVAL_1618;
  reg [31:0] _RAND_100;
  wire  _EVAL_1621;
  wire [31:0] _EVAL_1623;
  wire  _EVAL_1626;
  reg [3:0] _EVAL_1629;
  reg [31:0] _RAND_101;
  wire  _EVAL_1630;
  wire [31:0] _EVAL_1632;
  wire  _EVAL_1637;
  reg  _EVAL_1641;
  reg [31:0] _RAND_102;
  wire [31:0] _EVAL_1643;
  wire [31:0] _EVAL_1644;
  reg  _EVAL_1645;
  reg [31:0] _RAND_103;
  wire [31:0] _EVAL_1646;
  wire [17:0] _EVAL_1648;
  wire  _EVAL_1654;
  wire  _EVAL_1656;
  wire  _EVAL_1659;
  wire [2:0] _EVAL_1662;
  reg  _EVAL_1664;
  reg [31:0] _RAND_104;
  wire  _EVAL_1665;
  wire  _EVAL_1666;
  wire  _EVAL_1668;
  wire  _EVAL_1669;
  reg  _EVAL_1670;
  reg [31:0] _RAND_105;
  reg  _EVAL_1671;
  reg [31:0] _RAND_106;
  reg [3:0] _EVAL_1672;
  reg [31:0] _RAND_107;
  wire [15:0] _EVAL_1674;
  reg [3:0] _EVAL_1676;
  reg [31:0] _RAND_108;
  wire [31:0] _EVAL_1678;
  wire [31:0] _EVAL_1680;
  wire  _EVAL_1681;
  wire  _EVAL_1682;
  wire  _EVAL_1683;
  reg [7:0] _EVAL_1686;
  reg [31:0] _RAND_109;
  wire [4:0] _EVAL_1688;
  wire [15:0] _EVAL_1690;
  wire [9:0] _EVAL_1693;
  wire [31:0] _EVAL_1698;
  wire  _EVAL_1699;
  wire  _EVAL_1704;
  wire  _EVAL_1705;
  wire  _EVAL_1706;
  wire [31:0] _EVAL_1710;
  wire [31:0] _EVAL_1712;
  wire  _EVAL_1713;
  wire  _EVAL_1714;
  reg [3:0] _EVAL_1720;
  reg [31:0] _RAND_110;
  wire  _EVAL_1726;
  reg  _EVAL_1730;
  reg [31:0] _RAND_111;
  wire  _EVAL_1732;
  wire  _EVAL_1737;
  wire [4:0] _EVAL_1738;
  wire [7:0] _EVAL_1740;
  wire [9:0] _EVAL_1744;
  reg [3:0] _EVAL_1746;
  reg [31:0] _RAND_112;
  wire  _EVAL_1748;
  wire  _EVAL_1749;
  wire  _EVAL_1751;
  wire  _EVAL_1753;
  wire  _EVAL_1758;
  wire [23:0] _EVAL_1759;
  wire [7:0] _EVAL_1760;
  wire  _EVAL_1761;
  wire  _EVAL_1762;
  wire [3:0] _EVAL_1763;
  reg  _EVAL_1765;
  reg [31:0] _RAND_113;
  wire  _EVAL_1766;
  wire  _EVAL_1768;
  wire  _EVAL_1770;
  wire [15:0] _EVAL_1771;
  reg [63:0] _EVAL_1775;
  reg [63:0] _RAND_114;
  reg  _EVAL_1777;
  reg [31:0] _RAND_115;
  wire  _EVAL_1779;
  wire  _EVAL_1780;
  wire [4:0] _EVAL_1785;
  wire [4:0] _EVAL_1787;
  wire  _EVAL_1788;
  wire  _EVAL_1790;
  wire [17:0] _EVAL_1791;
  wire [31:0] _EVAL_1796;
  reg [3:0] _EVAL_1797;
  reg [31:0] _RAND_116;
  wire [4:0] _EVAL_1799;
  wire [1:0] _EVAL_1803;
  wire  _EVAL_1805;
  wire  _EVAL_1806;
  wire  _EVAL_1809;
  wire [4:0] _EVAL_1812;
  wire [7:0] _EVAL_1813;
  wire  _EVAL_1815;
  wire [2:0] _EVAL_1817;
  reg  _EVAL_1820;
  reg [31:0] _RAND_117;
  wire [31:0] _EVAL_1821;
  reg [3:0] _EVAL_1822;
  reg [31:0] _RAND_118;
  wire [25:0] _EVAL_1823;
  wire  _EVAL_1825;
  reg  _EVAL_1826;
  reg [31:0] _RAND_119;
  wire [7:0] _EVAL_1827;
  reg [3:0] _EVAL_1828;
  reg [31:0] _RAND_120;
  wire [1:0] _EVAL_1829;
  reg  _EVAL_1831;
  reg [31:0] _RAND_121;
  wire  _EVAL_1834;
  wire  _EVAL_1842;
  wire  _EVAL_1843;
  wire  _EVAL_1844;
  wire  _EVAL_1848;
  wire [31:0] _EVAL_1849;
  wire  _EVAL_1851;
  wire [23:0] _EVAL_1855;
  wire [31:0] _EVAL_1857;
  wire [15:0] _EVAL_1859;
  wire  _EVAL_1860;
  reg [3:0] _EVAL_1863;
  reg [31:0] _RAND_122;
  wire  _EVAL_1864;
  wire  _EVAL_1866;
  wire [15:0] _EVAL_1868;
  wire  _EVAL_1871;
  wire [3:0] _EVAL_1872;
  wire [1:0] _EVAL_1874;
  reg  _EVAL_1875;
  reg [31:0] _RAND_123;
  wire  _EVAL_1877;
  reg  _EVAL_1880;
  reg [31:0] _RAND_124;
  reg [3:0] _EVAL_1882;
  reg [31:0] _RAND_125;
  wire [1:0] _EVAL_1883;
  wire  _EVAL_1885;
  wire [1:0] _EVAL_1886;
  wire  _EVAL_1890;
  reg [3:0] _EVAL_1891;
  reg [31:0] _RAND_126;
  wire [7:0] _EVAL_1892;
  wire [2:0] _EVAL_1898;
  wire [7:0] _EVAL_1899;
  wire  _EVAL_1900;
  wire  _EVAL_1901;
  wire  _EVAL_1903;
  wire [4:0] _EVAL_1904;
  wire  _EVAL_1907;
  wire  _EVAL_1908;
  wire [1:0] _EVAL_1912;
  wire [4:0] _EVAL_1914;
  reg  _EVAL_1917;
  reg [31:0] _RAND_127;
  wire [1:0] _EVAL_1918;
  wire  _EVAL_1922;
  wire [1:0] _EVAL_1923;
  wire [1:0] _EVAL_1925;
  wire [7:0] _EVAL_1927;
  reg  _EVAL_1929;
  reg [31:0] _RAND_128;
  wire [31:0] _EVAL_1930;
  wire  _EVAL_1934;
  wire  _EVAL_1935;
  wire  _EVAL_1937;
  wire [25:0] _EVAL_1939;
  reg  _EVAL_1942;
  reg [31:0] _RAND_129;
  wire [31:0] _EVAL_1943;
  wire  _EVAL_1949;
  wire [4:0] _EVAL_1950;
  wire [23:0] _EVAL_1952;
  wire [31:0] _EVAL_1953;
  wire  _EVAL_1956;
  wire [7:0] _EVAL_1959;
  wire [17:0] _EVAL_1961;
  wire [9:0] _EVAL_1963;
  wire [17:0] _EVAL_1964;
  wire  _EVAL_1967;
  wire [4:0] _EVAL_1968;
  wire [23:0] _EVAL_1969;
  wire [1:0] _EVAL_1970;
  wire [7:0] _EVAL_1976;
  wire  _EVAL_1979;
  wire  _EVAL_1982;
  wire [4:0] _EVAL_1983;
  wire [17:0] _EVAL_1987;
  wire  _EVAL_1990;
  wire [4:0] _EVAL_1997;
  wire [4:0] _EVAL_1998;
  wire  _EVAL_1999;
  wire [4:0] _EVAL_2003;
  wire [2:0] _EVAL_2004;
  reg  _EVAL_2009;
  reg [31:0] _RAND_130;
  wire [23:0] _EVAL_2010;
  wire  _EVAL_2013;
  wire [7:0] _EVAL_2016;
  wire [1:0] _EVAL_2017;
  wire  _EVAL_2018;
  wire  _EVAL_2020;
  wire  _EVAL_2022;
  wire [31:0] _EVAL_2024;
  wire  _EVAL_2025;
  wire [31:0] _EVAL_2026;
  wire [1:0] _EVAL_2029;
  reg [3:0] _EVAL_2030;
  reg [31:0] _RAND_131;
  wire  _EVAL_2034;
  wire  _EVAL_2036;
  wire  _EVAL_2042;
  wire  _EVAL_2046;
  wire [1:0] _EVAL_2047;
  wire  _EVAL_2048;
  wire  _EVAL_2050;
  wire  _EVAL_2052;
  wire [1:0] _EVAL_2053;
  wire [4:0] _EVAL_2054;
  wire [4:0] _EVAL_2055;
  wire [31:0] _EVAL_2056;
  wire  _EVAL_2057;
  wire  _EVAL_2058;
  wire [15:0] _EVAL_2061;
  wire  _EVAL_2063;
  reg  _EVAL_2065;
  reg [31:0] _RAND_132;
  wire  _EVAL_2070;
  wire  _EVAL_2074;
  wire  _EVAL_2077;
  wire [4:0] _EVAL_2080;
  wire  _EVAL_2081;
  wire [23:0] _EVAL_2085;
  reg  _EVAL_2086;
  reg [31:0] _RAND_133;
  wire [1:0] _EVAL_2090;
  wire  _EVAL_2091;
  wire  _EVAL_2092;
  wire [15:0] _EVAL_2094;
  reg  _EVAL_2096;
  reg [31:0] _RAND_134;
  wire  _EVAL_2098;
  wire [31:0] _EVAL_2099;
  wire  _EVAL_2101;
  wire [9:0] _EVAL_2102;
  wire  _EVAL_2104;
  wire  _EVAL_2105;
  wire  _EVAL_2108;
  wire [1:0] _EVAL_2109;
  wire  _EVAL_2111;
  wire  _EVAL_2112;
  wire [25:0] _EVAL_2113;
  wire [5:0] _EVAL_2114;
  wire [4:0] _EVAL_2115;
  wire  _EVAL_2119;
  wire [1:0] _EVAL_2120;
  wire [23:0] _EVAL_2122;
  wire  _EVAL_2128;
  wire  _EVAL_2130;
  wire [9:0] _EVAL_2132;
  wire [2:0] _EVAL_2136;
  wire [25:0] _EVAL_2137;
  wire [1:0] _EVAL_2138;
  wire [1:0] _EVAL_2139;
  wire  _EVAL_2141;
  wire [31:0] _EVAL_2143;
  wire [4:0] _EVAL_2146;
  wire [31:0] _EVAL_2147;
  reg  _EVAL_2148;
  reg [31:0] _RAND_135;
  wire [23:0] _EVAL_2152;
  reg  _EVAL_2154;
  reg [31:0] _RAND_136;
  wire  _EVAL_2155;
  wire [17:0] _EVAL_2156;
  wire [15:0] _EVAL_2157;
  wire [7:0] _EVAL_2158;
  wire [4:0] _EVAL_2159;
  wire  _EVAL_2160;
  wire  _EVAL_2161;
  reg  _EVAL_2162;
  reg [31:0] _RAND_137;
  wire [31:0] _EVAL_2164;
  wire  _EVAL_2166;
  wire  _EVAL_2168;
  wire  _EVAL_2173;
  wire  _EVAL_2176;
  reg  _EVAL_2177;
  reg [31:0] _RAND_138;
  wire [31:0] _EVAL_2178;
  wire  _EVAL_2180;
  wire [1:0] _EVAL_2182;
  reg [3:0] _EVAL_2183;
  reg [31:0] _RAND_139;
  wire [2:0] _EVAL_2185;
  wire [31:0] _EVAL_2186;
  wire [4:0] _EVAL_2188;
  wire  _EVAL_2189;
  wire  _EVAL_2190;
  wire [25:0] _EVAL_2196;
  wire  _EVAL_2197;
  wire  _EVAL_2198;
  wire  _EVAL_2199;
  wire  _EVAL_2201;
  wire  _EVAL_2202;
  reg  _EVAL_2203;
  reg [31:0] _RAND_140;
  wire [31:0] _EVAL_2206;
  wire [23:0] _EVAL_2211;
  wire  _EVAL_2212;
  reg  _EVAL_2215;
  reg [31:0] _RAND_141;
  wire  _EVAL_2216;
  reg [63:0] _EVAL_2218;
  reg [63:0] _RAND_142;
  wire  _EVAL_2225;
  wire [25:0] _EVAL_2226;
  wire [4:0] _EVAL_2227;
  wire [4:0] _EVAL_2228;
  reg  _EVAL_2229;
  reg [31:0] _RAND_143;
  wire [3:0] _EVAL_2231;
  reg  _EVAL_2233;
  reg [31:0] _RAND_144;
  wire [31:0] _EVAL_2234;
  wire [63:0] _EVAL_2237;
  wire  _EVAL_2239;
  wire [25:0] _EVAL_2240;
  wire  _EVAL_2244;
  reg  _EVAL_2247;
  reg [31:0] _RAND_145;
  wire [31:0] _EVAL_2248;
  wire  _EVAL_2249;
  wire [23:0] _EVAL_2257;
  wire  _EVAL_2259;
  wire [4:0] _EVAL_2261;
  wire [31:0] _EVAL_2263;
  wire [25:0] _EVAL_2264;
  wire  _EVAL_2265;
  wire [1:0] _EVAL_2267;
  wire [1:0] _EVAL_2276;
  reg  _EVAL_2277;
  reg [31:0] _RAND_146;
  wire [31:0] _EVAL_2279;
  wire  _EVAL_2281;
  wire [23:0] _EVAL_2282;
  wire [9:0] _EVAL_2283;
  wire  _EVAL_2286;
  wire  _EVAL_2287;
  wire  _EVAL_2289;
  reg  _EVAL_2291;
  reg [31:0] _RAND_147;
  reg [3:0] _EVAL_2293;
  reg [31:0] _RAND_148;
  wire  _EVAL_2300;
  reg  _EVAL_2301;
  reg [31:0] _RAND_149;
  wire [9:0] _EVAL_2303;
  reg [3:0] _EVAL_2307;
  reg [31:0] _RAND_150;
  reg  _EVAL_2308;
  reg [31:0] _RAND_151;
  wire [25:0] _EVAL_2309;
  wire  _EVAL_2311;
  reg  _EVAL_2312;
  reg [31:0] _RAND_152;
  wire [4:0] _EVAL_2315;
  wire  _EVAL_2316;
  wire [31:0] _EVAL_2319;
  wire  _EVAL_2322;
  wire  _EVAL_2324;
  wire [25:0] _EVAL_2330;
  wire  _EVAL_2331;
  wire [4:0] _EVAL_2332;
  wire [25:0] _EVAL_2336;
  wire [23:0] _EVAL_2337;
  reg  _EVAL_2339;
  reg [31:0] _RAND_153;
  reg  _EVAL_2341;
  reg [31:0] _RAND_154;
  wire  _EVAL_2342;
  wire  _EVAL_2343;
  wire  _EVAL_2346;
  wire [4:0] _EVAL_2348;
  wire  _EVAL_2350;
  wire  _EVAL_2351;
  wire  _EVAL_2352;
  wire [17:0] _EVAL_2353;
  reg  _EVAL_2357;
  reg [31:0] _RAND_155;
  wire [4:0] _EVAL_2359;
  reg  _EVAL_2360;
  reg [31:0] _RAND_156;
  wire [31:0] _EVAL_2365;
  reg  _EVAL_2366;
  reg [31:0] _RAND_157;
  wire  _EVAL_2369;
  wire  _EVAL_2372;
  wire  _EVAL_2374;
  wire  _EVAL_2377;
  wire  _EVAL_2380;
  reg  _EVAL_2381;
  reg [31:0] _RAND_158;
  wire [4:0] _EVAL_2385;
  wire [7:0] _EVAL_2389;
  wire [31:0] _EVAL_2391;
  wire  _EVAL_2392;
  reg [3:0] _EVAL_2393;
  reg [31:0] _RAND_159;
  wire  _EVAL_2394;
  wire [25:0] _EVAL_2396;
  wire  _EVAL_2398;
  wire  _EVAL_2400;
  wire  _EVAL_2406;
  wire  _EVAL_2407;
  wire [23:0] _EVAL_2408;
  wire [17:0] _EVAL_2410;
  wire  _EVAL_2413;
  wire [23:0] _EVAL_2415;
  wire  _EVAL_2417;
  wire [25:0] _EVAL_2418;
  wire  _EVAL_2421;
  reg  _EVAL_2422;
  reg [31:0] _RAND_160;
  wire  _EVAL_2428;
  wire [1:0] _EVAL_2429;
  wire [17:0] _EVAL_2434;
  wire [31:0] _EVAL_2435;
  wire [23:0] _EVAL_2439;
  reg  _EVAL_2444;
  reg [31:0] _RAND_161;
  wire  _EVAL_2446;
  wire [31:0] _EVAL_2447;
  wire [9:0] _EVAL_2448;
  wire [31:0] _EVAL_2450;
  wire  _EVAL_2457;
  wire  _EVAL_2461;
  reg [3:0] _EVAL_2462;
  reg [31:0] _RAND_162;
  wire [1:0] _EVAL_2463;
  wire [4:0] _EVAL_2467;
  wire  _EVAL_2470;
  wire  _EVAL_2473;
  wire  _EVAL_2474;
  wire  _EVAL_2477;
  wire  _EVAL_2481;
  reg  _EVAL_2484;
  reg [31:0] _RAND_163;
  wire  _EVAL_2486;
  wire [15:0] _EVAL_2487;
  wire [15:0] _EVAL_2488;
  wire  _EVAL_2489;
  reg [3:0] _EVAL_2490;
  reg [31:0] _RAND_164;
  wire [31:0] _EVAL_2491;
  wire [7:0] _EVAL_2492;
  reg [3:0] _EVAL_2493;
  reg [31:0] _RAND_165;
  wire  _EVAL_2495;
  wire  _EVAL_2499;
  wire [31:0] _EVAL_2501;
  wire  _EVAL_2503;
  wire [15:0] _EVAL_2508;
  wire  _EVAL_2510;
  wire [31:0] _EVAL_2512;
  wire  _EVAL_2515;
  reg  _EVAL_2516;
  reg [31:0] _RAND_166;
  wire  _EVAL_2519;
  wire  _EVAL_2520;
  wire  _EVAL_2521;
  wire [4:0] _EVAL_2522;
  wire  _EVAL_2523;
  wire  _EVAL_2527;
  wire  _EVAL_2528;
  wire  _EVAL_2530;
  wire [1:0] _EVAL_2532;
  wire [25:0] _EVAL_2534;
  wire [31:0] _EVAL_2535;
  reg [3:0] _EVAL_2537;
  reg [31:0] _RAND_167;
  wire  _EVAL_2541;
  wire [31:0] _EVAL_2543;
  wire [31:0] _EVAL_2544;
  reg [3:0] _EVAL_2546;
  reg [31:0] _RAND_168;
  wire [15:0] _EVAL_2547;
  wire [23:0] _EVAL_2549;
  reg [3:0] _EVAL_2557;
  reg [31:0] _RAND_169;
  wire [1:0] _EVAL_2559;
  reg [3:0] _EVAL_2561;
  reg [31:0] _RAND_170;
  wire [25:0] _EVAL_2563;
  wire  _EVAL_2566;
  wire  _EVAL_2568;
  wire  _EVAL_2575;
  wire  _EVAL_2577;
  wire  _EVAL_2578;
  wire [23:0] _EVAL_2579;
  reg  _EVAL_2580;
  reg [31:0] _RAND_171;
  reg  _EVAL_2583;
  reg [31:0] _RAND_172;
  wire [23:0] _EVAL_2586;
  wire  _EVAL_2587;
  reg  _EVAL_2589;
  reg [31:0] _RAND_173;
  wire [1:0] _EVAL_2590;
  wire [1:0] _EVAL_2591;
  wire  _EVAL_2595;
  wire  _EVAL_2596;
  wire  _EVAL_2598;
  wire [15:0] _EVAL_2600;
  wire  _EVAL_2603;
  wire  _EVAL_2605;
  wire [4:0] _EVAL_2610;
  wire  _EVAL_2611;
  reg  _EVAL_2616;
  reg [31:0] _RAND_174;
  wire [31:0] _EVAL_2618;
  wire  _EVAL_2621;
  wire  _EVAL_2622;
  wire [9:0] _EVAL_2623;
  reg [3:0] _EVAL_2626;
  reg [31:0] _RAND_175;
  reg [3:0] _EVAL_2629;
  reg [31:0] _RAND_176;
  wire  _EVAL_2630;
  wire  _EVAL_2633;
  wire  _EVAL_2635;
  wire [4:0] _EVAL_2636;
  wire [15:0] _EVAL_2637;
  wire  _EVAL_2638;
  wire [2:0] _EVAL_2639;
  wire [23:0] _EVAL_2641;
  wire [3:0] _EVAL_2642;
  wire  _EVAL_2648;
  wire [31:0] _EVAL_2654;
  wire  _EVAL_2660;
  wire  _EVAL_2661;
  wire [31:0] _EVAL_2664;
  wire  _EVAL_2666;
  reg  _EVAL_2667;
  reg [31:0] _RAND_177;
  wire  _EVAL_2668;
  reg  _EVAL_2669;
  reg [31:0] _RAND_178;
  wire [1:0] _EVAL_2671;
  wire  _EVAL_2674;
  wire [15:0] _EVAL_2681;
  wire  _EVAL_2683;
  reg  _EVAL_2690;
  reg [31:0] _RAND_179;
  wire  _EVAL_2691;
  wire [1:0] _EVAL_2692;
  wire  _EVAL_2693;
  wire [17:0] _EVAL_2694;
  wire [2:0] _EVAL_2696;
  wire [31:0] _EVAL_2697;
  wire  _EVAL_2701;
  wire  _EVAL_2703;
  wire  _EVAL_2706;
  wire  _EVAL_2707;
  wire [1:0] _EVAL_2709;
  wire  _EVAL_2711;
  wire  _EVAL_2714;
  wire [15:0] _EVAL_2716;
  reg  _EVAL_2717;
  reg [31:0] _RAND_180;
  wire  _EVAL_2719;
  wire [25:0] _EVAL_2722;
  wire [31:0] _EVAL_2727;
  wire  _EVAL_2728;
  wire  _EVAL_2737;
  wire [1:0] _EVAL_2739;
  wire  _EVAL_2740;
  wire  _EVAL_2741;
  wire  _EVAL_2743;
  wire [31:0] _EVAL_2747;
  wire [1:0] _EVAL_2749;
  wire [4:0] _EVAL_2751;
  wire [4:0] _EVAL_2752;
  wire  _EVAL_2755;
  wire  _EVAL_2756;
  wire  _EVAL_2757;
  wire  _EVAL_2758;
  wire  _EVAL_2760;
  wire [4:0] _EVAL_2761;
  wire  _EVAL_2764;
  wire [1:0] _EVAL_2765;
  reg  _EVAL_2766;
  reg [31:0] _RAND_181;
  wire [9:0] _EVAL_2767;
  wire [4:0] _EVAL_2774;
  wire [9:0] _EVAL_2776;
  wire [9:0] _EVAL_2777;
  reg  _EVAL_2778;
  reg [31:0] _RAND_182;
  wire  _EVAL_2779;
  wire [31:0] _EVAL_2780;
  reg [3:0] _EVAL_2781;
  reg [31:0] _RAND_183;
  reg  _EVAL_2782;
  reg [31:0] _RAND_184;
  wire  _EVAL_2784;
  wire [1:0] _EVAL_2786;
  wire [4:0] _EVAL_2787;
  wire [4:0] _EVAL_2788;
  wire [7:0] _EVAL_2794;
  wire [15:0] _EVAL_2797;
  wire  _EVAL_2800;
  wire [31:0] _EVAL_2801;
  wire [31:0] _EVAL_2802;
  wire  _EVAL_2804;
  wire [4:0] _EVAL_2805;
  reg [3:0] _EVAL_2806;
  reg [31:0] _RAND_185;
  wire [31:0] _EVAL_2811;
  wire [31:0] _EVAL_2812;
  wire  _EVAL_2813;
  wire  _EVAL_2815;
  wire [4:0] _EVAL_2819;
  wire [2:0] _EVAL_2820;
  wire  _EVAL_2823;
  wire [4:0] _EVAL_2824;
  reg  _EVAL_2825;
  reg [31:0] _RAND_186;
  reg [3:0] _EVAL_2827;
  reg [31:0] _RAND_187;
  reg  _EVAL_2828;
  reg [31:0] _RAND_188;
  wire  _EVAL_2829;
  wire [17:0] _EVAL_2832;
  reg  _EVAL_2837;
  reg [31:0] _RAND_189;
  wire  _EVAL_2838;
  wire [31:0] _EVAL_2840;
  wire  _EVAL_2841;
  wire [1:0] _EVAL_2843;
  wire [17:0] _EVAL_2845;
  reg  _EVAL_2847;
  reg [31:0] _RAND_190;
  wire [4:0] _EVAL_2848;
  wire  _EVAL_2851;
  wire  _EVAL_2852;
  wire [31:0] _EVAL_2853;
  wire [9:0] _EVAL_2854;
  wire  _EVAL_2855;
  wire [2:0] _EVAL_2856;
  wire  _EVAL_2857;
  wire  _EVAL_2861;
  wire  _EVAL_2862;
  wire  _EVAL_2864;
  wire [7:0] _EVAL_2865;
  wire [25:0] _EVAL_2866;
  wire  _EVAL_2867;
  wire [4:0] _EVAL_2869;
  wire [31:0] _EVAL_2874;
  reg  _EVAL_2876;
  reg [31:0] _RAND_191;
  wire [17:0] _EVAL_2878;
  wire  _EVAL_2880;
  wire [31:0] _EVAL_2882;
  wire [4:0] _EVAL_2883;
  wire  _EVAL_2884;
  wire [1:0] _EVAL_2887;
  reg [3:0] _EVAL_2889;
  reg [31:0] _RAND_192;
  wire [9:0] _EVAL_2894;
  wire  _EVAL_2895;
  wire [31:0] _EVAL_2896;
  wire  _EVAL_2898;
  wire [17:0] _EVAL_2901;
  reg  _EVAL_2905;
  reg [31:0] _RAND_193;
  reg  _EVAL_2910;
  reg [31:0] _RAND_194;
  wire  _EVAL_2912;
  wire  _EVAL_2914;
  wire  _EVAL_2915;
  reg  _EVAL_2918;
  reg [31:0] _RAND_195;
  reg [3:0] _EVAL_2920;
  reg [31:0] _RAND_196;
  wire  _EVAL_2922;
  wire [2:0] _EVAL_2928;
  wire  _EVAL_2929;
  wire [31:0] _EVAL_2932;
  wire  _EVAL_2933;
  wire  _EVAL_2935;
  wire  _EVAL_2936;
  wire  _EVAL_2938;
  wire [7:0] _EVAL_2940;
  wire  _EVAL_2943;
  wire [31:0] _EVAL_2944;
  wire [3:0] _EVAL_2948;
  wire [31:0] _EVAL_2949;
  wire [7:0] _EVAL_2951;
  wire  _EVAL_2952;
  wire  _EVAL_2954;
  wire  _EVAL_2958;
  wire [1:0] _EVAL_2959;
  wire  _EVAL_2961;
  wire [7:0] _EVAL_2964;
  wire [4:0] _EVAL_2967;
  wire  _EVAL_2968;
  wire [7:0] _EVAL_2970;
  wire [1:0] _EVAL_2971;
  wire [3:0] _EVAL_2978;
  wire  _EVAL_2979;
  wire  _EVAL_2980;
  wire [23:0] _EVAL_2981;
  reg [3:0] _EVAL_2984;
  reg [31:0] _RAND_197;
  reg  _EVAL_2988;
  reg [31:0] _RAND_198;
  wire [15:0] _EVAL_2989;
  reg  _EVAL_2993;
  reg [31:0] _RAND_199;
  wire [4:0] _EVAL_2994;
  wire [9:0] _EVAL_2995;
  wire [15:0] _EVAL_2996;
  wire [1:0] _EVAL_2997;
  reg  _EVAL_3001;
  reg [31:0] _RAND_200;
  wire [7:0] _EVAL_3003;
  reg [3:0] _EVAL_3005;
  reg [31:0] _RAND_201;
  wire [25:0] _EVAL_3011;
  wire [1:0] _EVAL_3012;
  wire  _EVAL_3016;
  wire [25:0] _EVAL_3017;
  wire [1:0] _EVAL_3018;
  wire [17:0] _EVAL_3019;
  wire [23:0] _EVAL_3020;
  wire [9:0] _EVAL_3022;
  wire [4:0] _EVAL_3023;
  wire [7:0] _EVAL_3024;
  wire [2:0] _EVAL_3027;
  wire  _EVAL_3030;
  wire  _EVAL_3031;
  wire [4:0] _EVAL_3035;
  wire  _EVAL_3036;
  wire [4:0] _EVAL_3037;
  wire  _EVAL_3039;
  reg [3:0] _EVAL_3040;
  reg [31:0] _RAND_202;
  wire [1:0] _EVAL_3042;
  wire  _EVAL_3043;
  wire  _EVAL_3044;
  wire [31:0] _EVAL_3045;
  wire [4:0] _EVAL_3046;
  wire [3:0] _EVAL_3047;
  wire [7:0] _EVAL_3048;
  wire  _EVAL_3051;
  wire  _EVAL_3053;
  wire  _EVAL_3056;
  wire [7:0] _EVAL_3058;
  wire [31:0] _EVAL_3059;
  reg [3:0] _EVAL_3062;
  reg [31:0] _RAND_203;
  wire [2:0] _EVAL_3064;
  wire [4:0] _EVAL_3067;
  wire  _EVAL_3080;
  wire  _EVAL_3083;
  wire  _EVAL_3086;
  wire  _EVAL_3087;
  wire  _EVAL_3088;
  wire  _EVAL_3090;
  wire  _EVAL_3092;
  wire  _EVAL_3093;
  wire  _EVAL_3094;
  wire [1:0] _EVAL_3096;
  wire [17:0] _EVAL_3098;
  wire  _EVAL_3099;
  wire  _EVAL_3100;
  wire [7:0] _EVAL_3102;
  wire  _EVAL_3104;
  wire  _EVAL_3105;
  reg [3:0] _EVAL_3108;
  reg [31:0] _RAND_204;
  wire  _EVAL_3110;
  wire [1:0] _EVAL_3111;
  wire [1:0] _EVAL_3114;
  wire [31:0] _EVAL_3115;
  wire [4:0] _EVAL_3119;
  wire [1:0] _EVAL_3120;
  wire [23:0] _EVAL_3123;
  wire [2:0] _EVAL_3125;
  wire [4:0] _EVAL_3126;
  wire [7:0] _EVAL_3127;
  wire [4:0] _EVAL_3128;
  reg  _EVAL_3129;
  reg [31:0] _RAND_205;
  wire [4:0] _EVAL_3131;
  reg  _EVAL_3133;
  reg [31:0] _RAND_206;
  wire  _EVAL_3140;
  wire [23:0] _EVAL_3141;
  wire [4:0] _EVAL_3144;
  wire  _EVAL_3145;
  wire  _EVAL_3146;
  wire [31:0] _EVAL_3148;
  wire [15:0] _EVAL_3149;
  wire  _EVAL_3150;
  reg  _EVAL_3152;
  reg [31:0] _RAND_207;
  wire  _EVAL_3154;
  wire  _EVAL_3158;
  wire  _EVAL_3164;
  wire [25:0] _EVAL_3168;
  wire  _EVAL_3169;
  reg  _EVAL_3171;
  reg [31:0] _RAND_208;
  reg [3:0] _EVAL_3172;
  reg [31:0] _RAND_209;
  reg [3:0] _EVAL_3173;
  reg [31:0] _RAND_210;
  reg  _EVAL_3181;
  reg [31:0] _RAND_211;
  wire  _EVAL_3189;
  wire [7:0] _EVAL_3190;
  wire [4:0] _EVAL_3191;
  wire  _EVAL_3193;
  reg  _EVAL_3194;
  reg [31:0] _RAND_212;
  reg  _EVAL_3196;
  reg [31:0] _RAND_213;
  reg  _EVAL_3197;
  reg [31:0] _RAND_214;
  wire  _EVAL_3200;
  reg  _EVAL_3203;
  reg [31:0] _RAND_215;
  wire [31:0] _EVAL_3204;
  wire  _EVAL_3205;
  wire  _EVAL_3207;
  wire  _EVAL_3211;
  wire  _EVAL_3212;
  reg  _EVAL_3213;
  reg [31:0] _RAND_216;
  wire  _EVAL_3215;
  wire  _EVAL_3217;
  wire [4:0] _EVAL_3219;
  wire  _EVAL_3222;
  reg  _EVAL_3225;
  reg [31:0] _RAND_217;
  wire [31:0] _EVAL_3229;
  wire  _EVAL_3230;
  wire  _EVAL_3233;
  reg  _EVAL_3234;
  reg [31:0] _RAND_218;
  wire  _EVAL_3253;
  wire [25:0] _EVAL_3254;
  wire  _EVAL_3255;
  reg [3:0] _EVAL_3256;
  reg [31:0] _RAND_219;
  wire [25:0] _EVAL_3259;
  wire  _EVAL_3266;
  wire [31:0] _EVAL_3268;
  wire [4:0] _EVAL_3270;
  wire [31:0] _EVAL_3271;
  wire [17:0] _EVAL_3272;
  wire  _EVAL_3273;
  wire [1:0] _EVAL_3274;
  wire [4:0] _EVAL_3275;
  wire [31:0] _EVAL_3277;
  wire  _EVAL_3278;
  reg  _EVAL_3280;
  reg [31:0] _RAND_220;
  wire  _EVAL_3283;
  wire  _EVAL_3285;
  reg  _EVAL_3286;
  reg [31:0] _RAND_221;
  wire [7:0] _EVAL_3289;
  wire  _EVAL_3290;
  wire [31:0] _EVAL_3291;
  wire  _EVAL_3293;
  reg  _EVAL_3294;
  reg [31:0] _RAND_222;
  wire [31:0] _EVAL_3297;
  wire  _EVAL_3298;
  wire [7:0] _EVAL_3299;
  wire  _EVAL_3304;
  wire  _EVAL_3308;
  wire [1:0] _EVAL_3309;
  reg [3:0] _EVAL_3310;
  reg [31:0] _RAND_223;
  wire  _EVAL_3311;
  wire  _EVAL_3317;
  wire  _EVAL_3318;
  wire  _EVAL_3319;
  wire [2:0] _EVAL_3320;
  wire  _EVAL_3324;
  wire  _EVAL_3325;
  reg  _EVAL_3327;
  reg [31:0] _RAND_224;
  wire [7:0] _EVAL_3330;
  wire [31:0] _EVAL_3332;
  wire [15:0] _EVAL_3334;
  wire [2:0] _EVAL_3335;
  wire  _EVAL_3336;
  wire  _EVAL_3339;
  wire  _EVAL_3341;
  wire [7:0] _EVAL_3343;
  wire  _EVAL_3344;
  wire  _EVAL_3345;
  wire  _EVAL_3351;
  wire [4:0] _EVAL_3353;
  wire [7:0] _EVAL_3355;
  wire [31:0] _EVAL_3356;
  wire [25:0] _EVAL_3357;
  wire  _EVAL_3358;
  wire [31:0] _EVAL_3359;
  reg  _EVAL_3363;
  reg [31:0] _RAND_225;
  wire  _EVAL_3365;
  wire [4:0] _EVAL_3368;
  wire  _EVAL_3372;
  reg  _EVAL_3374;
  reg [31:0] _RAND_226;
  wire  _EVAL_3378;
  wire [4:0] _EVAL_3380;
  wire [1:0] _EVAL_3383;
  reg  _EVAL_3384;
  reg [31:0] _RAND_227;
  wire [19:0] _EVAL_3385;
  wire  _EVAL_3389;
  wire  _EVAL_3390;
  wire  _EVAL_3391;
  wire [31:0] _EVAL_3392;
  wire [4:0] _EVAL_3393;
  wire [31:0] _EVAL_3395;
  wire  _EVAL_3397;
  reg  _EVAL_3404;
  reg [31:0] _RAND_228;
  wire  _EVAL_3405;
  wire  _EVAL_3408;
  wire  _EVAL_3410;
  wire [3:0] _EVAL_3411;
  wire [9:0] _EVAL_3415;
  wire [1:0] _EVAL_3416;
  wire  _EVAL_3419;
  wire  _EVAL_3422;
  wire [64:0] _EVAL_3423;
  wire  _EVAL_3426;
  wire [3:0] _EVAL_3427;
  wire [2:0] _EVAL_3428;
  reg [3:0] _EVAL_3429;
  reg [31:0] _RAND_229;
  wire [4:0] _EVAL_3430;
  wire [4:0] _EVAL_3431;
  wire  _EVAL_3434;
  wire  _EVAL_3435;
  wire  _EVAL_3438;
  wire  _EVAL_3439;
  wire  _EVAL_3441;
  wire  _EVAL_3442;
  wire  _EVAL_3443;
  wire [8:0] _EVAL_3444;
  wire  _EVAL_3446;
  reg [3:0] _EVAL_3449;
  reg [31:0] _RAND_230;
  reg  _EVAL_3450;
  reg [31:0] _RAND_231;
  wire [7:0] _EVAL_3452;
  wire [4:0] _EVAL_3454;
  reg  _EVAL_3456;
  reg [31:0] _RAND_232;
  wire [5:0] _EVAL_3460;
  wire [23:0] _EVAL_3463;
  reg [3:0] _EVAL_3464;
  reg [31:0] _RAND_233;
  wire [4:0] _EVAL_3465;
  wire  _EVAL_3466;
  reg [3:0] _EVAL_3467;
  reg [31:0] _RAND_234;
  wire [4:0] _EVAL_3469;
  wire  _EVAL_3472;
  wire  _EVAL_3475;
  wire  _EVAL_3477;
  wire  _EVAL_3479;
  wire [31:0] _EVAL_3482;
  wire [4:0] _EVAL_3483;
  wire  _EVAL_3487;
  wire  _EVAL_3493;
  wire [25:0] _EVAL_3494;
  wire  _EVAL_3496;
  wire  _EVAL_3498;
  wire  _EVAL_3499;
  wire  _EVAL_3501;
  wire  _EVAL_3502;
  wire [7:0] _EVAL_3504;
  wire [31:0] _EVAL_3507;
  wire  _EVAL_3513;
  wire  _EVAL_3516;
  wire  _EVAL_3517;
  wire [4:0] _EVAL_3518;
  wire  _EVAL_3521;
  wire [4:0] _EVAL_3526;
  wire [1:0] _EVAL_3527;
  wire  _EVAL_3530;
  wire [2:0] _EVAL_3532;
  wire  _EVAL_3533;
  wire [3:0] _EVAL_3534;
  wire  _EVAL_3535;
  wire  _EVAL_3537;
  reg [3:0] _EVAL_3538;
  reg [31:0] _RAND_235;
  wire [1:0] _EVAL_3541;
  wire  _EVAL_3542;
  wire  _EVAL_3544;
  wire  _EVAL_3546;
  wire [23:0] _EVAL_3549;
  wire [23:0] _EVAL_3550;
  wire [9:0] _EVAL_3554;
  wire [2:0] _EVAL_3555;
  wire [31:0] _EVAL_3559;
  wire [17:0] _EVAL_3560;
  wire  _EVAL_3561;
  wire  _EVAL_3563;
  wire  _EVAL_3564;
  wire [1:0] _EVAL_3567;
  wire [1:0] _EVAL_3570;
  wire [1:0] _EVAL_3573;
  wire [31:0] _EVAL_3576;
  wire [31:0] _EVAL_3578;
  reg  _EVAL_3580;
  reg [31:0] _RAND_236;
  reg  _EVAL_3584;
  reg [31:0] _RAND_237;
  wire [4:0] _EVAL_3585;
  wire [2:0] _EVAL_3587;
  reg  _EVAL_3589;
  reg [31:0] _RAND_238;
  wire  _EVAL_3590;
  wire  _EVAL_3591;
  reg  _EVAL_3594;
  reg [31:0] _RAND_239;
  wire  _EVAL_3597;
  wire [4:0] _EVAL_3599;
  wire  _EVAL_3603;
  wire [1:0] _EVAL_3604;
  wire  intsink__EVAL;
  wire  intsink__EVAL_0;
  wire  intsink__EVAL_1;
  wire  intsink__EVAL_2;
  wire [31:0] _EVAL_3605;
  wire [31:0] _EVAL_3606;
  reg  _EVAL_3607;
  reg [31:0] _RAND_240;
  reg  _EVAL_3609;
  reg [31:0] _RAND_241;
  wire [1:0] _EVAL_3612;
  wire  _EVAL_3613;
  wire [23:0] _EVAL_3614;
  wire  _EVAL_3615;
  wire  _EVAL_3618;
  wire  _EVAL_3619;
  wire  _EVAL_3620;
  wire  _EVAL_3621;
  wire [31:0] _EVAL_3623;
  wire [1:0] _EVAL_3625;
  wire  _EVAL_3627;
  reg  _EVAL_3629;
  reg [31:0] _RAND_242;
  wire [17:0] _EVAL_3633;
  reg  _EVAL_3634;
  reg [31:0] _RAND_243;
  wire  _EVAL_3635;
  wire  _EVAL_3636;
  wire  _EVAL_3637;
  reg  _EVAL_3639;
  reg [31:0] _RAND_244;
  wire  _EVAL_3641;
  wire  _EVAL_3642;
  wire [31:0] _EVAL_3643;
  wire  _EVAL_3644;
  wire [7:0] _EVAL_3645;
  wire  _EVAL_3646;
  reg  _EVAL_3652;
  reg [31:0] _RAND_245;
  wire [31:0] _EVAL_3653;
  wire [4:0] _EVAL_3654;
  wire [4:0] _EVAL_3656;
  wire [31:0] _EVAL_3661;
  wire  _EVAL_3662;
  wire  _EVAL_3665;
  wire [31:0] _EVAL_3666;
  wire  _EVAL_3667;
  wire  _EVAL_3668;
  wire  _EVAL_3670;
  wire  _EVAL_3671;
  reg [3:0] _EVAL_3673;
  reg [31:0] _RAND_246;
  wire [7:0] _EVAL_3674;
  wire  _EVAL_3675;
  reg [3:0] _EVAL_3676;
  reg [31:0] _RAND_247;
  wire  _EVAL_3681;
  wire [7:0] _EVAL_3682;
  wire  _EVAL_3683;
  wire [4:0] _EVAL_3685;
  wire  _EVAL_3686;
  reg [3:0] _EVAL_3692;
  reg [31:0] _RAND_248;
  reg [3:0] _EVAL_3693;
  reg [31:0] _RAND_249;
  wire [2:0] _EVAL_3696;
  wire [17:0] _EVAL_3697;
  wire [1:0] _EVAL_3703;
  wire  _EVAL_3705;
  wire [3:0] _EVAL_3709;
  wire [7:0] _EVAL_3711;
  wire [31:0] _EVAL_3713;
  wire [9:0] _EVAL_3715;
  wire  _EVAL_3716;
  wire  _EVAL_3717;
  reg [3:0] _EVAL_3722;
  reg [31:0] _RAND_250;
  wire [1:0] _EVAL_3724;
  wire [4:0] _EVAL_3726;
  wire [25:0] _EVAL_3729;
  wire  _EVAL_3731;
  wire [31:0] _EVAL_3732;
  wire [1:0] _EVAL_3733;
  wire  _EVAL_3735;
  wire  _EVAL_3737;
  wire  _EVAL_3739;
  wire [31:0] _EVAL_3741;
  wire [25:0] _EVAL_3742;
  reg [3:0] _EVAL_3743;
  reg [31:0] _RAND_251;
  wire [1:0] _EVAL_3745;
  wire  _EVAL_3748;
  wire [4:0] _EVAL_3750;
  wire [17:0] _EVAL_3751;
  wire  _EVAL_3752;
  wire  _EVAL_3753;
  wire  _EVAL_3756;
  wire  _EVAL_3757;
  wire  _EVAL_3758;
  wire  _EVAL_3762;
  wire  _EVAL_3763;
  wire  _EVAL_3765;
  reg [3:0] _EVAL_3767;
  reg [31:0] _RAND_252;
  reg [3:0] _EVAL_3771;
  reg [31:0] _RAND_253;
  wire  _EVAL_3772;
  wire  _EVAL_3775;
  wire [1:0] _EVAL_3779;
  reg  _EVAL_3783;
  reg [31:0] _RAND_254;
  wire  _EVAL_3786;
  wire [31:0] _EVAL_3788;
  reg  _EVAL_3789;
  reg [31:0] _RAND_255;
  wire [4:0] _EVAL_3790;
  wire [31:0] _EVAL_3791;
  wire [1:0] _EVAL_3793;
  wire  _EVAL_3795;
  wire [4:0] _EVAL_3796;
  wire [31:0] _EVAL_3797;
  wire  _EVAL_3798;
  wire  _EVAL_3799;
  wire [31:0] _EVAL_3800;
  wire  _EVAL_3805;
  wire [17:0] _EVAL_3806;
  wire [3:0] _EVAL_3808;
  wire  _EVAL_3810;
  wire  _EVAL_3814;
  wire [2:0] _EVAL_3819;
  wire [4:0] _EVAL_3823;
  wire [2:0] _EVAL_3824;
  wire  _EVAL_3827;
  wire  _EVAL_3831;
  wire [7:0] _EVAL_3832;
  wire [4:0] _EVAL_3834;
  wire [15:0] _EVAL_3836;
  wire [6:0] _EVAL_3838;
  wire  _EVAL_3839;
  reg  _EVAL_3843;
  reg [31:0] _RAND_256;
  wire [7:0] _EVAL_3846;
  reg  _EVAL_3847;
  reg [31:0] _RAND_257;
  wire  _EVAL_3848;
  wire [4:0] _EVAL_3851;
  wire  _EVAL_3854;
  wire [2:0] _EVAL_3855;
  reg [3:0] _EVAL_3857;
  reg [31:0] _RAND_258;
  wire  _EVAL_3861;
  wire [1:0] _EVAL_3862;
  wire  _EVAL_3864;
  wire  _EVAL_3865;
  reg  _EVAL_3866;
  reg [31:0] _RAND_259;
  wire [4:0] _EVAL_3870;
  wire [25:0] _EVAL_3871;
  wire  _EVAL_3872;
  wire  _EVAL_3876;
  wire [4:0] _EVAL_3877;
  wire  _EVAL_3879;
  wire [25:0] _EVAL_3883;
  wire [17:0] _EVAL_3885;
  reg  _EVAL_3887;
  reg [31:0] _RAND_260;
  wire  _EVAL_3890;
  wire  _EVAL_3891;
  wire  _EVAL_3892;
  wire [4:0] _EVAL_3893;
  wire [3:0] _EVAL_3895;
  wire  _EVAL_3899;
  wire  _EVAL_3900;
  wire [4:0] _EVAL_3903;
  wire  _EVAL_3905;
  wire [4:0] _EVAL_3906;
  wire [17:0] _EVAL_3907;
  wire  _EVAL_3911;
  wire  _EVAL_3912;
  wire [15:0] _EVAL_3913;
  reg  _EVAL_3914;
  reg [31:0] _RAND_261;
  wire [9:0] _EVAL_3915;
  wire  _EVAL_3916;
  wire [15:0] _EVAL_3918;
  wire  _EVAL_3921;
  wire  _EVAL_3922;
  wire  _EVAL_3925;
  wire  _EVAL_3927;
  wire [1:0] _EVAL_3929;
  wire [31:0] _EVAL_3930;
  wire  _EVAL_3934;
  wire [31:0] _EVAL_3936;
  wire [4:0] _EVAL_3937;
  wire [31:0] _EVAL_3938;
  wire  _EVAL_3939;
  reg  _EVAL_3940;
  reg [31:0] _RAND_262;
  wire  _EVAL_3941;
  wire  _EVAL_3944;
  reg [3:0] _EVAL_3945;
  reg [31:0] _RAND_263;
  reg  _EVAL_3946;
  reg [31:0] _RAND_264;
  wire [31:0] _EVAL_3947;
  wire [15:0] _EVAL_3950;
  wire  _EVAL_3958;
  wire [31:0] _EVAL_3960;
  reg  _EVAL_3962;
  reg [31:0] _RAND_265;
  wire [4:0] _EVAL_3963;
  reg  _EVAL_3965;
  reg [31:0] _RAND_266;
  wire  _EVAL_3967;
  wire [31:0] _EVAL_3970;
  wire [25:0] _EVAL_3971;
  wire [1:0] _EVAL_3975;
  wire  _EVAL_3977;
  wire  _EVAL_3979;
  wire  _EVAL_3980;
  reg  _EVAL_3983;
  reg [31:0] _RAND_267;
  wire  _EVAL_3985;
  reg  _EVAL_3986;
  reg [31:0] _RAND_268;
  wire  _EVAL_3987;
  wire  _EVAL_3989;
  wire [4:0] _EVAL_3997;
  wire  _EVAL_3999;
  wire [4:0] _EVAL_4000;
  wire  _EVAL_4003;
  wire [17:0] _EVAL_4004;
  wire  _EVAL_4005;
  reg  _EVAL_4007;
  reg [31:0] _RAND_269;
  wire  _EVAL_4008;
  wire  _EVAL_4009;
  wire  _EVAL_4010;
  wire  _EVAL_4012;
  wire  _EVAL_4013;
  reg  _EVAL_4014;
  reg [31:0] _RAND_270;
  wire  _EVAL_4015;
  reg [3:0] _EVAL_4019;
  reg [31:0] _RAND_271;
  wire [2:0] _EVAL_4021;
  wire  _EVAL_4025;
  wire [4:0] _EVAL_4026;
  wire  _EVAL_4030;
  wire  _EVAL_4032;
  wire [25:0] _EVAL_4036;
  wire [1:0] _EVAL_4037;
  reg [3:0] _EVAL_4040;
  reg [31:0] _RAND_272;
  wire [25:0] _EVAL_4041;
  reg  _EVAL_4045;
  reg [31:0] _RAND_273;
  wire [1:0] _EVAL_4046;
  wire [1:0] _EVAL_4050;
  reg  _EVAL_4051;
  reg [31:0] _RAND_274;
  reg  _EVAL_4053;
  reg [31:0] _RAND_275;
  wire [4:0] _EVAL_4055;
  wire [23:0] _EVAL_4056;
  wire [4:0] _EVAL_4058;
  wire [4:0] _EVAL_4064;
  reg  _EVAL_4065;
  reg [31:0] _RAND_276;
  wire  _EVAL_4067;
  wire  _EVAL_4068;
  wire [6:0] _EVAL_4070;
  wire  _EVAL_4074;
  wire [1:0] _EVAL_4076;
  reg  _EVAL_4080;
  reg [31:0] _RAND_277;
  wire [25:0] _EVAL_4081;
  reg  _EVAL_4085;
  reg [31:0] _RAND_278;
  reg  _EVAL_4087;
  reg [31:0] _RAND_279;
  wire [3:0] _EVAL_4088;
  wire [4:0] _EVAL_4089;
  wire [25:0] _EVAL_4090;
  wire  _EVAL_4096;
  wire [7:0] _EVAL_4098;
  reg  _EVAL_4103;
  reg [31:0] _RAND_280;
  wire [23:0] _EVAL_4105;
  wire [1:0] _EVAL_4107;
  wire  _EVAL_4115;
  wire  _EVAL_4116;
  wire  _EVAL_4117;
  reg  _EVAL_4119;
  reg [31:0] _RAND_281;
  wire [1:0] _EVAL_4122;
  wire [17:0] _EVAL_4123;
  wire  _EVAL_4124;
  wire  _EVAL_4127;
  wire  _EVAL_4128;
  wire  _EVAL_4131;
  wire  _EVAL_4136;
  wire  _EVAL_4142;
  wire [15:0] _EVAL_4143;
  wire [1:0] _EVAL_4147;
  wire [7:0] _EVAL_4148;
  wire  _EVAL_4153;
  wire [25:0] _EVAL_4156;
  wire  _EVAL_4159;
  wire [23:0] _EVAL_4161;
  wire  _EVAL_4162;
  wire  _EVAL_4164;
  wire [4:0] _EVAL_4165;
  wire  _EVAL_4167;
  wire  _EVAL_4168;
  wire [4:0] _EVAL_4169;
  wire [1:0] _EVAL_4170;
  wire [23:0] _EVAL_4172;
  wire [17:0] _EVAL_4173;
  wire  _EVAL_4174;
  wire [4:0] _EVAL_4176;
  wire  _EVAL_4177;
  wire [4:0] _EVAL_4178;
  wire [7:0] _EVAL_4179;
  reg [3:0] _EVAL_4181;
  reg [31:0] _RAND_282;
  wire [4:0] _EVAL_4182;
  reg  _EVAL_4184;
  reg [31:0] _RAND_283;
  wire [17:0] _EVAL_4195;
  wire [31:0] _EVAL_4197;
  wire  _EVAL_4198;
  wire  _EVAL_4199;
  wire  _EVAL_4204;
  wire [3:0] _EVAL_4213;
  wire  _EVAL_4215;
  wire [15:0] _EVAL_4217;
  wire [9:0] _EVAL_4221;
  wire  _EVAL_4226;
  wire [4:0] _EVAL_4229;
  reg  _EVAL_4233;
  reg [31:0] _RAND_284;
  wire [1:0] _EVAL_4234;
  wire  _EVAL_4236;
  wire [1:0] _EVAL_4237;
  wire [25:0] _EVAL_4238;
  wire  _EVAL_4242;
  wire  _EVAL_4244;
  wire  _EVAL_4246;
  wire  _EVAL_4247;
  wire [2:0] _EVAL_4249;
  wire  _EVAL_4250;
  wire [23:0] _EVAL_4251;
  wire  _EVAL_4252;
  wire  _EVAL_4255;
  wire [1:0] _EVAL_4256;
  wire [31:0] _EVAL_4260;
  wire [1:0] _EVAL_4262;
  reg [3:0] _EVAL_4264;
  reg [31:0] _RAND_285;
  wire [4:0] _EVAL_4266;
  wire [31:0] _EVAL_4267;
  wire  _EVAL_4268;
  wire  _EVAL_4271;
  wire  _EVAL_4272;
  wire [4:0] _EVAL_4274;
  wire [9:0] _EVAL_4275;
  wire  _EVAL_4282;
  wire  _EVAL_4284;
  wire [31:0] _EVAL_4285;
  wire [25:0] _EVAL_4286;
  wire [9:0] _EVAL_4290;
  reg  _EVAL_4291;
  reg [31:0] _RAND_286;
  wire [17:0] _EVAL_4292;
  wire [23:0] _EVAL_4296;
  wire  _EVAL_4297;
  wire [31:0] _EVAL_4298;
  wire  _EVAL_4301;
  wire  _EVAL_4303;
  reg [3:0] _EVAL_4304;
  reg [31:0] _RAND_287;
  wire [17:0] _EVAL_4307;
  reg  _EVAL_4308;
  reg [31:0] _RAND_288;
  wire [23:0] _EVAL_4313;
  wire  _EVAL_4318;
  wire [1:0] _EVAL_4321;
  wire [1:0] _EVAL_4328;
  wire  _EVAL_4331;
  reg  _EVAL_4336;
  reg [31:0] _RAND_289;
  wire  _EVAL_4337;
  reg  _EVAL_4338;
  reg [31:0] _RAND_290;
  wire  _EVAL_4339;
  wire  _EVAL_4340;
  wire  _EVAL_4344;
  wire  _EVAL_4345;
  wire [7:0] _EVAL_4347;
  reg  _EVAL_4348;
  reg [31:0] _RAND_291;
  wire  _EVAL_4349;
  wire [4:0] _EVAL_4352;
  wire [4:0] _EVAL_4354;
  wire  _EVAL_4355;
  wire  _EVAL_4356;
  wire [31:0] _EVAL_4358;
  wire [25:0] _EVAL_4360;
  reg  _EVAL_4367;
  reg [31:0] _RAND_292;
  wire [7:0] _EVAL_4368;
  wire  _EVAL_4370;
  reg  _EVAL_4374;
  reg [31:0] _RAND_293;
  wire [4:0] _EVAL_4376;
  wire  _EVAL_4377;
  wire  _EVAL_4382;
  wire  _EVAL_4384;
  wire  _EVAL_4386;
  wire [4:0] _EVAL_4387;
  wire [6:0] _EVAL_4388;
  reg [3:0] _EVAL_4390;
  reg [31:0] _RAND_294;
  wire  _EVAL_4396;
  reg  _EVAL_4397;
  reg [31:0] _RAND_295;
  reg  _EVAL_4398;
  reg [31:0] _RAND_296;
  wire [9:0] _EVAL_4400;
  wire  _EVAL_4401;
  wire  _EVAL_4402;
  wire  _EVAL_4403;
  reg [3:0] _EVAL_4404;
  reg [31:0] _RAND_297;
  wire  _EVAL_4406;
  wire  _EVAL_4410;
  wire  _EVAL_4412;
  wire  _EVAL_4414;
  wire  _EVAL_4415;
  reg [3:0] _EVAL_4416;
  reg [31:0] _RAND_298;
  wire [9:0] _EVAL_4417;
  wire [15:0] _EVAL_4418;
  wire [31:0] _EVAL_4421;
  wire [9:0] _EVAL_4425;
  wire [23:0] _EVAL_4426;
  wire  _EVAL_4437;
  wire [7:0] _EVAL_4438;
  wire  _EVAL_4440;
  wire  _EVAL_4441;
  reg  _EVAL_4443;
  reg [31:0] _RAND_299;
  wire [4:0] _EVAL_4445;
  wire [31:0] _EVAL_4446;
  wire  _EVAL_4448;
  wire  _EVAL_4449;
  wire  _EVAL_4452;
  wire  _EVAL_4456;
  wire [4:0] _EVAL_4458;
  wire  _EVAL_4465;
  wire  _EVAL_4466;
  wire  _EVAL_4467;
  wire  _EVAL_4469;
  wire [4:0] _EVAL_4474;
  wire  _EVAL_4476;
  wire  _EVAL_4477;
  wire  _EVAL_4478;
  reg [3:0] _EVAL_4479;
  reg [31:0] _RAND_300;
  wire  _EVAL_4480;
  wire [4:0] _EVAL_4482;
  wire [4:0] _EVAL_4483;
  wire [3:0] _EVAL_4484;
  wire  _EVAL_4486;
  wire [7:0] _EVAL_4489;
  wire [7:0] _EVAL_4490;
  wire [23:0] _EVAL_4493;
  wire [1:0] _EVAL_4496;
  wire [1:0] _EVAL_4497;
  wire  _EVAL_4500;
  wire [1:0] _EVAL_4505;
  wire [9:0] _EVAL_4508;
  wire [17:0] _EVAL_4509;
  wire  _EVAL_4510;
  wire [4:0] _EVAL_4511;
  wire [15:0] _EVAL_4515;
  wire  _EVAL_4517;
  reg [3:0] _EVAL_4518;
  reg [31:0] _RAND_301;
  wire [31:0] _EVAL_4520;
  wire  _EVAL_4523;
  wire [2:0] _EVAL_4526;
  wire [7:0] _EVAL_4528;
  wire [4:0] _EVAL_4530;
  wire  _EVAL_4532;
  wire [1:0] _EVAL_4534;
  wire [9:0] _EVAL_4538;
  wire  _EVAL_4539;
  wire [4:0] _EVAL_4540;
  wire [1:0] _EVAL_4541;
  wire [31:0] _EVAL_4542;
  wire [31:0] _EVAL_4546;
  wire  _EVAL_4547;
  wire  _EVAL_4548;
  wire  _EVAL_4549;
  wire  _EVAL_4553;
  wire  _EVAL_4554;
  wire  _EVAL_4556;
  wire  _EVAL_4562;
  wire  _EVAL_4566;
  wire [15:0] _EVAL_4569;
  reg [3:0] _EVAL_4571;
  reg [31:0] _RAND_302;
  reg  _EVAL_4572;
  reg [31:0] _RAND_303;
  reg [3:0] _EVAL_4574;
  reg [31:0] _RAND_304;
  wire  _EVAL_4578;
  wire [25:0] _EVAL_4580;
  wire  _EVAL_4582;
  wire  _EVAL_4583;
  reg  _EVAL_4584;
  reg [31:0] _RAND_305;
  reg  _EVAL_4588;
  reg [31:0] _RAND_306;
  wire [7:0] _EVAL_4590;
  wire [3:0] _EVAL_4595;
  wire  _EVAL_4599;
  wire [1:0] _EVAL_4600;
  wire  _EVAL_4602;
  wire [4:0] _EVAL_4603;
  wire  _EVAL_4606;
  wire  _EVAL_4610;
  wire [2:0] _EVAL_4611;
  reg  _EVAL_4612;
  reg [31:0] _RAND_307;
  wire  _EVAL_4614;
  wire [17:0] _EVAL_4615;
  reg  _EVAL_4620;
  reg [31:0] _RAND_308;
  wire  _EVAL_4621;
  wire [23:0] _EVAL_4622;
  reg [3:0] _EVAL_4624;
  reg [31:0] _RAND_309;
  wire  _EVAL_4626;
  reg [3:0] _EVAL_4631;
  reg [31:0] _RAND_310;
  wire [4:0] _EVAL_4632;
  wire [4:0] _EVAL_4633;
  wire  _EVAL_4634;
  wire [4:0] _EVAL_4636;
  wire  _EVAL_4637;
  wire [1:0] _EVAL_4638;
  wire [7:0] _EVAL_4640;
  wire [1:0] _EVAL_4642;
  wire [4:0] _EVAL_4646;
  wire  _EVAL_4650;
  wire  _EVAL_4653;
  wire [4:0] _EVAL_4657;
  wire [2:0] _EVAL_4658;
  wire [31:0] _EVAL_4659;
  wire [25:0] _EVAL_4660;
  wire  _EVAL_4662;
  wire [31:0] _EVAL_4663;
  wire [31:0] _EVAL_4665;
  wire  _EVAL_4672;
  wire  _EVAL_4676;
  wire [1:0] _EVAL_4677;
  wire [15:0] _EVAL_4679;
  wire  _EVAL_4683;
  wire  _EVAL_4684;
  wire [7:0] _EVAL_4685;
  wire [2:0] _EVAL_4687;
  wire  _EVAL_4696;
  wire [4:0] _EVAL_4699;
  reg [3:0] _EVAL_4700;
  reg [31:0] _RAND_311;
  wire  _EVAL_4704;
  wire [7:0] _EVAL_4705;
  wire [15:0] _EVAL_4708;
  wire [3:0] _EVAL_4709;
  reg [3:0] _EVAL_4711;
  reg [31:0] _RAND_312;
  wire [31:0] _EVAL_4716;
  wire [4:0] _EVAL_4717;
  wire [23:0] _EVAL_4718;
  wire [2:0] _EVAL_4719;
  wire  _EVAL_4721;
  wire [63:0] _EVAL_4725;
  wire  _EVAL_4728;
  reg  _EVAL_4732;
  reg [31:0] _RAND_313;
  wire  _EVAL_4734;
  wire  _EVAL_4735;
  reg  _EVAL_4738;
  reg [31:0] _RAND_314;
  wire [4:0] _EVAL_4740;
  wire [7:0] _EVAL_4741;
  reg  _EVAL_4742;
  reg [31:0] _RAND_315;
  wire  _EVAL_4746;
  wire  _EVAL_4747;
  wire  _EVAL_4749;
  wire [4:0] _EVAL_4752;
  wire  _EVAL_4753;
  wire [4:0] _EVAL_4754;
  wire [25:0] _EVAL_4758;
  wire [25:0] _EVAL_4763;
  wire  _EVAL_4769;
  wire [4:0] _EVAL_4770;
  wire [31:0] _EVAL_4771;
  wire  _EVAL_4772;
  wire [25:0] _EVAL_4774;
  wire [4:0] _EVAL_4776;
  wire  _EVAL_4778;
  reg  _EVAL_4779;
  reg [31:0] _RAND_316;
  reg  _EVAL_4785;
  reg [31:0] _RAND_317;
  reg [3:0] _EVAL_4786;
  reg [31:0] _RAND_318;
  wire  _EVAL_4789;
  wire  _EVAL_4791;
  wire  _EVAL_4797;
  wire [31:0] _EVAL_4799;
  wire [31:0] _EVAL_4805;
  reg  _EVAL_4807;
  reg [31:0] _RAND_319;
  reg  _EVAL_4808;
  reg [31:0] _RAND_320;
  wire  _EVAL_4809;
  reg  _EVAL_4810;
  reg [31:0] _RAND_321;
  wire  _EVAL_4815;
  wire [4:0] _EVAL_4816;
  wire [1:0] _EVAL_4818;
  wire  _EVAL_4819;
  wire  _EVAL_4820;
  wire  _EVAL_4822;
  wire [25:0] _EVAL_4823;
  wire [27:0] _EVAL_4824;
  wire [15:0] _EVAL_4826;
  wire [4:0] _EVAL_4827;
  reg  _EVAL_4828;
  reg [31:0] _RAND_322;
  wire [1:0] _EVAL_4829;
  wire  _EVAL_4835;
  wire [25:0] _EVAL_4837;
  wire  _EVAL_4839;
  wire  _EVAL_4840;
  reg  _EVAL_4843;
  reg [31:0] _RAND_323;
  wire [17:0] _EVAL_4846;
  wire [7:0] _EVAL_4848;
  wire  _EVAL_4849;
  wire [15:0] _EVAL_4852;
  wire [31:0] _EVAL_4853;
  wire [4:0] _EVAL_4858;
  wire [25:0] _EVAL_4860;
  wire  _EVAL_4863;
  wire [4:0] _EVAL_4864;
  wire  _EVAL_4865;
  wire [4:0] _EVAL_4869;
  wire [17:0] _EVAL_4875;
  wire  _EVAL_4876;
  wire  _EVAL_4878;
  wire [2:0] _EVAL_4880;
  wire  _EVAL_4882;
  wire [4:0] _EVAL_4883;
  wire [7:0] _EVAL_4884;
  wire [17:0] _EVAL_4885;
  wire [2:0] _EVAL_4889;
  wire [31:0] _EVAL_4893;
  wire  _EVAL_4894;
  wire  _EVAL_4895;
  wire [25:0] _EVAL_4897;
  wire [9:0] _EVAL_4899;
  wire  _EVAL_4901;
  wire  _EVAL_4902;
  wire [1:0] _EVAL_4903;
  wire [7:0] _EVAL_4905;
  wire [31:0] _EVAL_4906;
  reg [3:0] _EVAL_4908;
  reg [31:0] _RAND_324;
  reg [3:0] _EVAL_4911;
  reg [31:0] _RAND_325;
  wire [4:0] _EVAL_4913;
  wire [23:0] _EVAL_4919;
  wire [31:0] _EVAL_4921;
  reg  _EVAL_4922;
  reg [31:0] _RAND_326;
  wire [1:0] _EVAL_4924;
  reg [3:0] _EVAL_4927;
  reg [31:0] _RAND_327;
  wire  _EVAL_4929;
  reg  _EVAL_4932;
  reg [31:0] _RAND_328;
  wire [15:0] _EVAL_4933;
  wire [1:0] _EVAL_4935;
  wire  _EVAL_4937;
  wire  _EVAL_4940;
  wire [25:0] _EVAL_4941;
  wire  _EVAL_4942;
  wire [4:0] _EVAL_4943;
  reg  _EVAL_4944;
  reg [31:0] _RAND_329;
  wire [3:0] _EVAL_4945;
  wire  _EVAL_4948;
  wire [4:0] _EVAL_4953;
  wire [23:0] _EVAL_4954;
  reg  _EVAL_4955;
  reg [31:0] _RAND_330;
  wire  _EVAL_4956;
  wire [5:0] _EVAL_4958;
  wire  _EVAL_4959;
  reg  _EVAL_4965;
  reg [31:0] _RAND_331;
  wire  _EVAL_4968;
  wire [25:0] _EVAL_4969;
  wire  _EVAL_4970;
  wire [9:0] _EVAL_4972;
  wire [4:0] _EVAL_4973;
  wire [9:0] _EVAL_4977;
  wire  _EVAL_4978;
  wire  _EVAL_4980;
  wire [7:0] _EVAL_4982;
  wire [23:0] _EVAL_4986;
  wire [6:0] _EVAL_4990;
  wire  _EVAL_4992;
  wire  _EVAL_4994;
  wire [7:0] _EVAL_4995;
  reg [3:0] _EVAL_4997;
  reg [31:0] _RAND_332;
  wire [1:0] _EVAL_4998;
  wire [7:0] _EVAL_5000;
  wire [25:0] _EVAL_5001;
  reg  _EVAL_5002;
  reg [31:0] _RAND_333;
  wire [31:0] _EVAL_5004;
  wire  _EVAL_5007;
  reg [3:0] _EVAL_5008;
  reg [31:0] _RAND_334;
  reg [3:0] _EVAL_5009;
  reg [31:0] _RAND_335;
  wire  _EVAL_5010;
  wire [4:0] _EVAL_5011;
  wire  _EVAL_5012;
  wire  _EVAL_5013;
  wire  _EVAL_5014;
  wire  _EVAL_5019;
  wire  _EVAL_5022;
  wire  _EVAL_5024;
  wire [31:0] _EVAL_5026;
  wire  _EVAL_5029;
  wire  _EVAL_5030;
  wire [7:0] _EVAL_5031;
  wire  _EVAL_5034;
  wire [31:0] _EVAL_5038;
  reg [3:0] _EVAL_5039;
  reg [31:0] _RAND_336;
  wire  _EVAL_5041;
  wire [4:0] _EVAL_5044;
  wire  _EVAL_5045;
  wire  _EVAL_5046;
  wire [1:0] _EVAL_5047;
  wire  _EVAL_5048;
  wire  _EVAL_5049;
  wire  _EVAL_5052;
  wire [4:0] _EVAL_5058;
  wire [17:0] _EVAL_5061;
  wire  _EVAL_5062;
  wire  _EVAL_5064;
  wire [15:0] _EVAL_5065;
  wire [1023:0] _EVAL_5068;
  wire  _EVAL_5070;
  wire  _EVAL_5073;
  reg [3:0] _EVAL_5080;
  reg [31:0] _RAND_337;
  wire  _EVAL_5086;
  wire  _EVAL_5089;
  wire  _EVAL_5093;
  wire [31:0] _EVAL_5095;
  wire  _EVAL_5096;
  wire [31:0] _EVAL_5097;
  wire [4:0] _EVAL_5098;
  reg  _EVAL_5101;
  reg [31:0] _RAND_338;
  reg  _EVAL_5104;
  reg [31:0] _RAND_339;
  wire [31:0] _EVAL_5106;
  wire [7:0] _EVAL_5107;
  wire  _EVAL_5108;
  wire  _EVAL_5109;
  wire  _EVAL_5111;
  wire [3:0] _EVAL_5112;
  wire  _EVAL_5113;
  wire  _EVAL_5115;
  wire [31:0] _EVAL_5117;
  wire  _EVAL_5120;
  wire  _EVAL_5125;
  wire [1:0] _EVAL_5126;
  wire  _EVAL_5131;
  wire [9:0] _EVAL_5137;
  reg [3:0] _EVAL_5139;
  reg [31:0] _RAND_340;
  wire [31:0] _EVAL_5140;
  reg [3:0] _EVAL_5142;
  reg [31:0] _RAND_341;
  wire  _EVAL_5143;
  wire  _EVAL_5145;
  wire [23:0] _EVAL_5146;
  reg  _EVAL_5147;
  reg [31:0] _RAND_342;
  wire  _EVAL_5150;
  wire  _EVAL_5151;
  wire  _EVAL_5154;
  wire [15:0] _EVAL_5156;
  reg  _EVAL_5163;
  reg [31:0] _RAND_343;
  wire  _EVAL_5164;
  wire [4:0] _EVAL_5165;
  wire [4:0] _EVAL_5166;
  wire  _EVAL_5168;
  wire  _EVAL_5169;
  wire [3:0] _EVAL_5171;
  wire  _EVAL_5172;
  wire  _EVAL_5174;
  wire [23:0] _EVAL_5176;
  wire [3:0] _EVAL_5180;
  wire [25:0] _EVAL_5181;
  wire [4:0] _EVAL_5183;
  wire [4:0] _EVAL_5185;
  wire [17:0] _EVAL_5186;
  wire  _EVAL_5188;
  reg  _EVAL_5190;
  reg [31:0] _RAND_344;
  wire [31:0] _EVAL_5191;
  wire  _EVAL_5195;
  wire [7:0] _EVAL_5197;
  wire [1:0] _EVAL_5198;
  wire [4:0] _EVAL_5202;
  wire  _EVAL_5203;
  wire [2:0] _EVAL_5204;
  wire [4:0] _EVAL_5220;
  wire  _EVAL_5221;
  wire  _EVAL_5222;
  wire [31:0] _EVAL_5224;
  wire  _EVAL_5225;
  wire [4:0] _EVAL_5227;
  wire [4:0] _EVAL_5231;
  reg  _EVAL_5232;
  reg [31:0] _RAND_345;
  wire [15:0] _EVAL_5237;
  wire [1:0] _EVAL_5244;
  wire [63:0] _EVAL_5247;
  wire [31:0] _EVAL_5248;
  reg  _EVAL_5249;
  reg [31:0] _RAND_346;
  wire  _EVAL_5253;
  wire [7:0] _EVAL_5254;
  reg  _EVAL_5255;
  reg [31:0] _RAND_347;
  wire  _EVAL_5256;
  wire [17:0] _EVAL_5257;
  wire  _EVAL_5258;
  wire [31:0] _EVAL_5262;
  wire [4:0] _EVAL_5263;
  wire [23:0] _EVAL_5265;
  wire  _EVAL_5266;
  wire  _EVAL_5267;
  wire  _EVAL_5269;
  wire [1:0] _EVAL_5270;
  wire  _EVAL_5275;
  wire  _EVAL_5278;
  wire [31:0] _EVAL_5279;
  wire [7:0] _EVAL_5287;
  wire  _EVAL_5288;
  wire [4:0] _EVAL_5290;
  reg  _EVAL_5293;
  reg [31:0] _RAND_348;
  wire  _EVAL_5294;
  wire [31:0] _EVAL_5295;
  wire [4:0] _EVAL_5297;
  reg  _EVAL_5300;
  reg [31:0] _RAND_349;
  wire [1:0] _EVAL_5301;
  reg  _EVAL_5307;
  reg [31:0] _RAND_350;
  reg  _EVAL_5309;
  reg [31:0] _RAND_351;
  reg [3:0] _EVAL_5311;
  reg [31:0] _RAND_352;
  wire [1:0] _EVAL_5312;
  wire  _EVAL_5314;
  reg  _EVAL_5315;
  reg [31:0] _RAND_353;
  wire [15:0] _EVAL_5318;
  wire [1:0] _EVAL_5321;
  wire [4:0] _EVAL_5322;
  wire [1:0] _EVAL_5323;
  wire [31:0] _EVAL_5324;
  wire [4:0] _EVAL_5325;
  wire  _EVAL_5326;
  wire  _EVAL_5330;
  wire  _EVAL_5331;
  wire  _EVAL_5332;
  wire [1:0] _EVAL_5333;
  wire [4:0] _EVAL_5334;
  wire  _EVAL_5335;
  wire  _EVAL_5337;
  wire  _EVAL_5339;
  wire  _EVAL_5340;
  reg  _EVAL_5345;
  reg [31:0] _RAND_354;
  wire [17:0] _EVAL_5346;
  wire  _EVAL_5348;
  wire  _EVAL_5350;
  wire [31:0] _EVAL_5358;
  wire [4:0] _EVAL_5359;
  wire  _EVAL_5363;
  wire [4:0] _EVAL_5364;
  wire [1:0] _EVAL_5366;
  reg  _EVAL_5369;
  reg [31:0] _RAND_355;
  wire [4:0] _EVAL_5373;
  wire  _EVAL_5374;
  wire  _EVAL_5375;
  wire [23:0] _EVAL_5377;
  wire [7:0] _EVAL_5378;
  wire  _EVAL_5382;
  wire [31:0] _EVAL_5384;
  reg  _EVAL_5386;
  reg [31:0] _RAND_356;
  wire [1:0] _EVAL_5388;
  reg [3:0] _EVAL_5389;
  reg [31:0] _RAND_357;
  wire  _EVAL_5390;
  wire  _EVAL_5391;
  wire [9:0] _EVAL_5392;
  wire [1:0] _EVAL_5393;
  wire [17:0] _EVAL_5394;
  reg  _EVAL_5396;
  reg [31:0] _RAND_358;
  wire  _EVAL_5397;
  wire  _EVAL_5399;
  wire  _EVAL_5403;
  wire  _EVAL_5405;
  wire [9:0] _EVAL_5406;
  wire [9:0] _EVAL_5407;
  reg  _EVAL_5409;
  reg [31:0] _RAND_359;
  wire [9:0] _EVAL_5410;
  reg  _EVAL_5411;
  reg [31:0] _RAND_360;
  wire [4:0] _EVAL_5413;
  wire [9:0] _EVAL_5415;
  wire  _EVAL_5421;
  wire [1:0] _EVAL_5426;
  wire  _EVAL_5429;
  wire  _EVAL_5432;
  wire  _EVAL_5435;
  wire [31:0] _EVAL_5436;
  wire [4:0] _EVAL_5441;
  wire [31:0] _EVAL_5442;
  wire  _EVAL_5448;
  wire [31:0] _EVAL_5453;
  wire  _EVAL_5459;
  wire [31:0] _EVAL_5460;
  wire  _EVAL_5462;
  wire [4:0] _EVAL_5463;
  wire [7:0] _EVAL_5467;
  wire  _EVAL_5468;
  wire  _EVAL_5469;
  wire  _EVAL_5472;
  wire  _EVAL_5475;
  reg  _EVAL_5479;
  reg [31:0] _RAND_361;
  wire [4:0] _EVAL_5480;
  wire  _EVAL_5481;
  reg  _EVAL_5484;
  reg [31:0] _RAND_362;
  wire  _EVAL_5485;
  wire [1:0] _EVAL_5487;
  wire  _EVAL_5491;
  wire  _EVAL_5494;
  wire [4:0] _EVAL_5495;
  wire [15:0] _EVAL_5499;
  wire [25:0] _EVAL_5501;
  wire [4:0] _EVAL_5503;
  wire [4:0] _EVAL_5504;
  wire  _EVAL_5505;
  wire  _EVAL_5506;
  wire  _EVAL_5511;
  wire [1:0] _EVAL_5513;
  wire [4:0] _EVAL_5515;
  wire  _EVAL_5516;
  reg [3:0] _EVAL_5518;
  reg [31:0] _RAND_363;
  wire  _EVAL_5519;
  wire  _EVAL_5520;
  reg  _EVAL_5521;
  reg [31:0] _RAND_364;
  wire [1:0] _EVAL_5522;
  wire [31:0] _EVAL_5523;
  wire [25:0] _EVAL_5526;
  wire [17:0] _EVAL_5533;
  reg  _EVAL_5535;
  reg [31:0] _RAND_365;
  wire [9:0] _EVAL_5536;
  reg [3:0] _EVAL_5537;
  reg [31:0] _RAND_366;
  wire  _EVAL_5539;
  wire  _EVAL_5540;
  wire [4:0] _EVAL_5545;
  wire  _EVAL_5546;
  wire [4:0] _EVAL_5547;
  wire  _EVAL_5548;
  wire [25:0] _EVAL_5550;
  wire [4:0] _EVAL_5551;
  wire [25:0] _EVAL_5552;
  wire [17:0] _EVAL_5553;
  wire [15:0] _EVAL_5554;
  wire [4:0] _EVAL_5555;
  wire  _EVAL_5556;
  wire  _EVAL_5557;
  reg  _EVAL_5558;
  reg [31:0] _RAND_367;
  wire [4:0] _EVAL_5562;
  wire  _EVAL_5563;
  wire [4:0] _EVAL_5567;
  wire  _EVAL_5571;
  wire  _EVAL_5577;
  wire [4:0] _EVAL_5579;
  wire [2:0] _EVAL_5580;
  wire [1:0] _EVAL_5581;
  wire  _EVAL_5582;
  wire [31:0] _EVAL_5584;
  wire  _EVAL_5585;
  wire  _EVAL_5591;
  wire  _EVAL_5595;
  wire  _EVAL_5597;
  reg  _EVAL_5600;
  reg [31:0] _RAND_368;
  wire  _EVAL_5603;
  wire  _EVAL_5605;
  reg [3:0] _EVAL_5606;
  reg [31:0] _RAND_369;
  reg  _EVAL_5608;
  reg [31:0] _RAND_370;
  reg  _EVAL_5609;
  reg [31:0] _RAND_371;
  wire  _EVAL_5611;
  wire [7:0] _EVAL_5612;
  wire [1:0] _EVAL_5614;
  wire  _EVAL_5615;
  wire  _EVAL_5617;
  wire  _EVAL_5619;
  wire [25:0] _EVAL_5621;
  reg [3:0] _EVAL_5623;
  reg [31:0] _RAND_372;
  reg [3:0] _EVAL_5624;
  reg [31:0] _RAND_373;
  wire [3:0] _EVAL_5626;
  wire  _EVAL_5627;
  wire  _EVAL_5628;
  reg  _EVAL_5629;
  reg [31:0] _RAND_374;
  reg  _EVAL_5635;
  reg [31:0] _RAND_375;
  wire  _EVAL_5636;
  wire  _EVAL_5637;
  wire [1:0] _EVAL_5638;
  wire  _EVAL_5644;
  wire [1:0] _EVAL_5645;
  wire  _EVAL_5646;
  wire [1:0] _EVAL_5653;
  wire [7:0] _EVAL_5655;
  wire  _EVAL_5657;
  wire [9:0] _EVAL_5658;
  wire [31:0] _EVAL_5660;
  wire [4:0] _EVAL_5661;
  reg [3:0] _EVAL_5665;
  reg [31:0] _RAND_376;
  reg [3:0] _EVAL_5667;
  reg [31:0] _RAND_377;
  wire [9:0] _EVAL_5669;
  reg [3:0] _EVAL_5670;
  reg [31:0] _RAND_378;
  wire  _EVAL_5674;
  reg  _EVAL_5675;
  reg [31:0] _RAND_379;
  wire  _EVAL_5677;
  wire [4:0] _EVAL_5681;
  wire  _EVAL_5682;
  wire  _EVAL_5683;
  reg  _EVAL_5684;
  reg [31:0] _RAND_380;
  wire [1:0] _EVAL_5687;
  wire [31:0] _EVAL_5689;
  wire [2:0] _EVAL_5690;
  wire [1:0] _EVAL_5691;
  wire [15:0] _EVAL_5694;
  reg  _EVAL_5696;
  reg [31:0] _RAND_381;
  reg [3:0] _EVAL_5697;
  reg [31:0] _RAND_382;
  wire [15:0] _EVAL_5698;
  wire  _EVAL_5699;
  wire [15:0] _EVAL_5701;
  wire [4:0] _EVAL_5706;
  wire [7:0] _EVAL_5709;
  wire [17:0] _EVAL_5710;
  wire  _EVAL_5711;
  wire [17:0] _EVAL_5712;
  reg [3:0] _EVAL_5713;
  reg [31:0] _RAND_383;
  wire [9:0] _EVAL_5714;
  wire  _EVAL_5715;
  wire  _EVAL_5716;
  wire  _EVAL_5717;
  wire [7:0] _EVAL_5718;
  wire [4:0] _EVAL_5719;
  wire [4:0] _EVAL_5725;
  reg [3:0] _EVAL_5727;
  reg [31:0] _RAND_384;
  wire [4:0] _EVAL_5728;
  wire  _EVAL_5730;
  wire [23:0] _EVAL_5731;
  wire [4:0] _EVAL_5732;
  reg  _EVAL_5735;
  reg [31:0] _RAND_385;
  wire [1:0] _EVAL_5738;
  reg  _EVAL_5741;
  reg [31:0] _RAND_386;
  wire [31:0] _EVAL_5742;
  reg  _EVAL_5743;
  reg [31:0] _RAND_387;
  wire  _EVAL_5745;
  wire [17:0] _EVAL_5746;
  wire  _EVAL_5748;
  wire [31:0] _EVAL_5749;
  wire  _EVAL_5751;
  wire [9:0] _EVAL_5757;
  wire  _EVAL_5758;
  wire  _EVAL_5759;
  wire  _EVAL_5762;
  wire [4:0] _EVAL_5763;
  reg [3:0] _EVAL_5765;
  reg [31:0] _RAND_388;
  wire [7:0] _EVAL_5767;
  wire [15:0] _EVAL_5768;
  wire  _EVAL_5769;
  wire [31:0] _EVAL_5770;
  wire  _EVAL_5771;
  wire  _EVAL_5777;
  wire  _EVAL_5780;
  reg  _EVAL_5781;
  reg [31:0] _RAND_389;
  wire  _EVAL_5782;
  wire [9:0] _EVAL_5783;
  wire [31:0] _EVAL_5785;
  wire  _EVAL_5787;
  wire  _EVAL_5791;
  wire  _EVAL_5792;
  wire [4:0] _EVAL_5793;
  wire [4:0] _EVAL_5794;
  wire  _EVAL_5799;
  wire  _EVAL_5800;
  wire  _EVAL_5801;
  wire  _EVAL_5802;
  wire [4:0] _EVAL_5803;
  wire [7:0] _EVAL_5804;
  wire [31:0] _EVAL_5805;
  wire  _EVAL_5806;
  wire [4:0] _EVAL_5807;
  wire [9:0] _EVAL_5808;
  wire  _EVAL_5813;
  wire  _EVAL_5815;
  wire [31:0] _EVAL_5817;
  wire  _EVAL_5818;
  wire [17:0] _EVAL_5820;
  wire  _EVAL_5821;
  wire [4:0] _EVAL_5824;
  wire [31:0] _EVAL_5828;
  wire  _EVAL_5829;
  wire [1:0] _EVAL_5830;
  wire  _EVAL_5833;
  wire  _EVAL_5835;
  wire  _EVAL_5836;
  wire  _EVAL_5841;
  wire [31:0] _EVAL_5844;
  reg  _EVAL_5846;
  reg [31:0] _RAND_390;
  wire [9:0] _EVAL_5847;
  wire [17:0] _EVAL_5849;
  wire  _EVAL_5851;
  wire [31:0] _EVAL_5852;
  wire [1:0] _EVAL_5859;
  wire  _EVAL_5860;
  wire [15:0] _EVAL_5861;
  wire  _EVAL_5862;
  wire [31:0] _EVAL_5863;
  wire [7:0] _EVAL_5864;
  wire [15:0] _EVAL_5865;
  wire [31:0] _EVAL_5870;
  wire  _EVAL_5871;
  wire  _EVAL_5872;
  wire  _EVAL_5873;
  wire [25:0] _EVAL_5875;
  wire [13:0] _EVAL_5876;
  reg  _EVAL_5878;
  reg [31:0] _RAND_391;
  wire  _EVAL_5881;
  wire  _EVAL_5883;
  wire [2:0] _EVAL_5884;
  wire  _EVAL_5885;
  reg  _EVAL_5890;
  reg [31:0] _RAND_392;
  wire [23:0] _EVAL_5891;
  wire  _EVAL_5894;
  wire  _EVAL_5898;
  wire [4:0] _EVAL_5899;
  wire [31:0] _EVAL_5901;
  wire  _EVAL_5903;
  wire [3:0] _EVAL_5905;
  wire  _EVAL_5906;
  wire  _EVAL_5907;
  wire [15:0] _EVAL_5908;
  wire  _EVAL_5909;
  wire [15:0] _EVAL_5910;
  wire [3:0] _EVAL_5913;
  wire [7:0] _EVAL_5915;
  reg  _EVAL_5916;
  reg [31:0] _RAND_393;
  wire [3:0] _EVAL_5918;
  wire [4:0] _EVAL_5923;
  reg  _EVAL_5924;
  reg [31:0] _RAND_394;
  wire [4:0] _EVAL_5925;
  wire [7:0] _EVAL_5926;
  wire  _EVAL_5928;
  wire  _EVAL_5929;
  wire  _EVAL_5931;
  wire  _EVAL_5933;
  wire [15:0] _EVAL_5934;
  wire  _EVAL_5935;
  wire  _EVAL_5939;
  reg  _EVAL_5940;
  reg [31:0] _RAND_395;
  wire  _EVAL_5942;
  wire [31:0] _EVAL_5944;
  wire [7:0] _EVAL_5949;
  wire  _EVAL_5951;
  wire [4:0] _EVAL_5952;
  wire  _EVAL_5957;
  wire [31:0] _EVAL_5958;
  wire  _EVAL_5960;
  wire [23:0] _EVAL_5961;
  reg [3:0] _EVAL_5962;
  reg [31:0] _RAND_396;
  wire [23:0] _EVAL_5963;
  wire  _EVAL_5965;
  wire  _EVAL_5966;
  wire  _EVAL_5967;
  wire [7:0] _EVAL_5969;
  wire [4:0] _EVAL_5972;
  reg [3:0] _EVAL_5981;
  reg [31:0] _RAND_397;
  wire  _EVAL_5983;
  wire  _EVAL_5984;
  reg  _EVAL_5985;
  reg [31:0] _RAND_398;
  wire [15:0] _EVAL_5989;
  wire  _EVAL_5993;
  wire  _EVAL_5995;
  wire [4:0] _EVAL_5996;
  wire  _EVAL_5997;
  wire  _EVAL_6000;
  wire  _EVAL_6004;
  wire [31:0] _EVAL_6006;
  wire  _EVAL_6009;
  wire  _EVAL_6012;
  wire [31:0] _EVAL_6013;
  wire  _EVAL_6014;
  wire [17:0] _EVAL_6016;
  wire [2:0] _EVAL_6018;
  wire [17:0] _EVAL_6019;
  wire [25:0] _EVAL_6020;
  reg  _EVAL_6021;
  reg [31:0] _RAND_399;
  wire  _EVAL_6023;
  wire  _EVAL_6025;
  wire [15:0] _EVAL_6027;
  reg  _EVAL_6030;
  reg [31:0] _RAND_400;
  wire [4:0] _EVAL_6031;
  wire [17:0] _EVAL_6034;
  wire  _EVAL_6035;
  reg [3:0] _EVAL_6040;
  reg [31:0] _RAND_401;
  wire [23:0] _EVAL_6041;
  wire  _EVAL_6042;
  wire  _EVAL_6043;
  wire [15:0] _EVAL_6044;
  wire  _EVAL_6046;
  wire  _EVAL_6049;
  wire  _EVAL_6052;
  wire  _EVAL_6053;
  wire  _EVAL_6056;
  wire [31:0] _EVAL_6058;
  wire  _EVAL_6060;
  wire  _EVAL_6061;
  wire [4:0] _EVAL_6063;
  wire  _EVAL_6064;
  wire [4:0] _EVAL_6066;
  wire [7:0] _EVAL_6067;
  wire  _EVAL_6071;
  wire [23:0] _EVAL_6072;
  wire  _EVAL_6073;
  wire  _EVAL_6074;
  wire  _EVAL_6078;
  wire [31:0] _EVAL_6079;
  wire  _EVAL_6081;
  wire [31:0] _EVAL_6082;
  wire [5:0] _EVAL_6091;
  wire  _EVAL_6092;
  reg  _EVAL_6098;
  reg [31:0] _RAND_402;
  wire [4:0] _EVAL_6100;
  wire  _EVAL_6101;
  _EVAL_115 Queue (
    ._EVAL(Queue__EVAL),
    ._EVAL_0(Queue__EVAL_0),
    ._EVAL_1(Queue__EVAL_1),
    ._EVAL_2(Queue__EVAL_2),
    ._EVAL_3(Queue__EVAL_3),
    ._EVAL_4(Queue__EVAL_4),
    ._EVAL_5(Queue__EVAL_5),
    ._EVAL_6(Queue__EVAL_6),
    ._EVAL_7(Queue__EVAL_7),
    ._EVAL_8(Queue__EVAL_8),
    ._EVAL_9(Queue__EVAL_9),
    ._EVAL_10(Queue__EVAL_10),
    ._EVAL_11(Queue__EVAL_11),
    ._EVAL_12(Queue__EVAL_12),
    ._EVAL_13(Queue__EVAL_13),
    ._EVAL_14(Queue__EVAL_14),
    ._EVAL_15(Queue__EVAL_15),
    ._EVAL_16(Queue__EVAL_16)
  );
  _EVAL_113 intsink (
    ._EVAL(intsink__EVAL),
    ._EVAL_0(intsink__EVAL_0),
    ._EVAL_1(intsink__EVAL_1),
    ._EVAL_2(intsink__EVAL_2)
  );
  assign _EVAL_505 = {{6'd0}, _EVAL_499};
  assign _EVAL_2811 = {{6'd0}, _EVAL_4837};
  assign _EVAL_3345 = _EVAL_1730 & _EVAL_1506;
  assign _EVAL_749 = {1'h0,_EVAL_5629};
  assign _EVAL_1872 = {{1'd0}, _EVAL_448};
  assign _EVAL_5262 = _EVAL_6025 ? _EVAL_190 : _EVAL_1435;
  assign _EVAL_5480 = {_EVAL_3053,_EVAL_5623};
  assign _EVAL_4852 = {{6'd0}, _EVAL_2623};
  assign _EVAL_2693 = _EVAL_5068[668];
  assign _EVAL_6034 = {1'h0,_EVAL_3171,_EVAL_6044};
  assign _EVAL_5297 = {_EVAL_229,_EVAL_1289};
  assign _EVAL_2042 = 10'h292 == _EVAL_5757;
  assign _EVAL_3365 = _EVAL_5068[589];
  assign _EVAL_556 = _EVAL_4556 & _EVAL_2350;
  assign _EVAL_2389 = {{6'd0}, _EVAL_5653};
  assign _EVAL_968 = _EVAL_5836 & _EVAL_2350;
  assign _EVAL_1950 = {_EVAL_5862,_EVAL_4997};
  assign _EVAL_5415 = {1'h0,_EVAL_4398,_EVAL_4368};
  assign _EVAL_3534 = {{1'd0}, _EVAL_2820};
  assign _EVAL_866 = _EVAL_4772 ? _EVAL_3653 : _EVAL_5852;
  assign _EVAL_3987 = _EVAL_5732 > 5'h0;
  assign _EVAL_2392 = _EVAL_3866 & _EVAL_3196;
  assign _EVAL_5001 = {1'h0,_EVAL_4087,_EVAL_838};
  assign _EVAL_403 = _EVAL_1770 ? _EVAL_715 : _EVAL_3268;
  assign _EVAL_1261 = _EVAL_4865 & _EVAL_3154;
  assign _EVAL_1705 = Queue__EVAL_8[12];
  assign _EVAL_945 = 10'h219 == _EVAL_5757;
  assign _EVAL_6031 = {_EVAL_5818,_EVAL_1318};
  assign _EVAL_4347 = {{6'd0}, _EVAL_5126};
  assign _EVAL_1890 = _EVAL_1686[4];
  assign _EVAL_3023 = {_EVAL_5506,_EVAL_2557};
  assign _EVAL_5258 = 10'h20f == _EVAL_5757;
  assign _EVAL_5782 = _EVAL_5068[586];
  assign _EVAL_4406 = _EVAL_5113 & _EVAL_417;
  assign _EVAL_2240 = {1'h0,_EVAL_3286,_EVAL_4251};
  assign _EVAL_5690 = 3'h4 | _EVAL_420;
  assign _EVAL_5169 = _EVAL_5068[672];
  assign _EVAL_5997 = _EVAL_5068[583];
  assign _EVAL_5337 = 10'h2a3 == _EVAL_5757;
  assign _EVAL_338 = Queue__EVAL[0];
  assign _EVAL_240 = {{6'd0}, _EVAL_4899};
  assign _EVAL_1265 = 2'h2 | _EVAL_167;
  assign _EVAL_5711 = _EVAL_5068[666];
  assign _EVAL_1899 = {{6'd0}, _EVAL_1923};
  assign _EVAL_3098 = {1'h0,_EVAL_2086,_EVAL_2600};
  assign _EVAL_3742 = {1'h0,_EVAL_4932,_EVAL_6072};
  assign _EVAL_301 = _EVAL_1323 | _EVAL_2091;
  assign _EVAL_1849 = _EVAL_2968 ? _EVAL_2543 : _EVAL_4260;
  assign _EVAL_2216 = _EVAL_5068[590];
  assign _EVAL_4418 = {{6'd0}, _EVAL_1693};
  assign _EVAL_4425 = {1'h0,_EVAL_507,_EVAL_1345};
  assign _EVAL_3681 = _EVAL_5951 & _EVAL_2216;
  assign _EVAL_806 = {{6'd0}, _EVAL_1823};
  assign _EVAL_4237 = {1'h0,_EVAL_3589};
  assign _EVAL_4884 = _EVAL_2218[63:56];
  assign _EVAL_5725 = {_EVAL_4271,_EVAL_5606};
  assign _EVAL_5653 = {1'h0,_EVAL_4374};
  assign _EVAL_4030 = _EVAL_1746 == 4'h8;
  assign _EVAL_203 = _EVAL_3814 & _EVAL_417;
  assign _EVAL_1089 = _EVAL_5068[654];
  assign _EVAL_4880 = _EVAL_4728 ? {{1'd0}, _EVAL_2090} : _EVAL_1174;
  assign _EVAL_2691 = _EVAL_3979 ? _EVAL_673 : _EVAL_2173;
  assign _EVAL_4331 = _EVAL_3834 > _EVAL_2055;
  assign _EVAL_2446 = _EVAL_4415 ? 1'h0 : 1'h1;
  assign _EVAL_3733 = {1'h0,_EVAL_5600};
  assign _EVAL_3215 = _EVAL_423 & _EVAL_673;
  assign _EVAL_4548 = _EVAL_2638 ? 1'h0 : 1'h1;
  assign _EVAL_3493 = _EVAL_796 & _EVAL_4477;
  assign _EVAL_5442 = {_EVAL_2984,4'hf,_EVAL_5008,4'hf,_EVAL_5670,4'hf,_EVAL_653,4'hf};
  assign _EVAL_1414 = _EVAL_2166 ? _EVAL_5413 : _EVAL_1688;
  assign _EVAL_4474 = _EVAL_2470 ? _EVAL_459 : _EVAL_2348;
  assign _EVAL_5421 = _EVAL_5432 & _EVAL_847;
  assign _EVAL_3550 = {{6'd0}, _EVAL_4885};
  assign _EVAL_4426 = {{6'd0}, _EVAL_180};
  assign _EVAL_3293 = _EVAL_1968 > 5'h0;
  assign _EVAL_4753 = _EVAL_5151 & _EVAL_2350;
  assign _EVAL_3644 = _EVAL_2583 & _EVAL_3946;
  assign _EVAL_2989 = {{6'd0}, _EVAL_3554};
  assign _EVAL_3434 = _EVAL_2778 & _EVAL_5781;
  assign _EVAL_1111 = _EVAL_1751 & _EVAL_417;
  assign _EVAL_978 = _EVAL_6073 & _EVAL_847;
  assign _EVAL_1400 = {{6'd0}, _EVAL_991};
  assign _EVAL_5550 = {1'h0,_EVAL_3404,24'h0};
  assign _EVAL_5966 = _EVAL_5629 & _EVAL_4732;
  assign _EVAL_3119 = {_EVAL_2666,_EVAL_5039};
  assign _EVAL_4937 = _EVAL_2155 & _EVAL_2756;
  assign _EVAL_1306 = {{1'd0}, _EVAL_2527};
  assign _EVAL_2901 = {1'h0,_EVAL_3652,_EVAL_3918};
  assign _EVAL_4948 = _EVAL_4089 > _EVAL_5263;
  assign _EVAL_5346 = {1'h0,_EVAL_2233,_EVAL_4418};
  assign _EVAL_2315 = {_EVAL_3410,_EVAL_1273};
  assign _EVAL_5331 = _EVAL_5064 & _EVAL_1937;
  assign _EVAL_3938 = _EVAL_3083 ? _EVAL_2654 : _EVAL_1279;
  assign _EVAL_4826 = {{6'd0}, _EVAL_1205};
  assign _EVAL_3913 = {{6'd0}, _EVAL_5406};
  assign _EVAL_2413 = _EVAL_3499 & _EVAL_3487;
  assign _EVAL_1217 = 10'h295 == _EVAL_5757;
  assign _EVAL_4448 = 10'h21e == _EVAL_5757;
  assign _EVAL_4906 = _EVAL_3671 ? _EVAL_4197 : _EVAL_2727;
  assign _EVAL_5626 = {{1'd0}, _EVAL_4021};
  assign _EVAL_6009 = _EVAL_2857 & _EVAL_847;
  assign _EVAL_3259 = {1'h0,_EVAL_3225,_EVAL_2152};
  assign _EVAL_2463 = {1'h0,_EVAL_891};
  assign _EVAL_6063 = {_EVAL_4599,_EVAL_4181};
  assign _EVAL_4182 = _EVAL_3477 ? _EVAL_2227 : _EVAL_4973;
  assign _EVAL_4396 = 10'h29c == _EVAL_5757;
  assign _EVAL_2264 = {1'h0,_EVAL_5293,_EVAL_2257};
  assign _EVAL_3339 = _EVAL_4994 & _EVAL_673;
  assign _EVAL_4360 = {1'h0,_EVAL_5190,_EVAL_3123};
  assign _EVAL_5926 = {{6'd0}, _EVAL_452};
  assign _EVAL_4465 = _EVAL_5108 | _EVAL_879;
  assign _EVAL_3285 = _EVAL_2380 & _EVAL_4477;
  assign _EVAL_835 = 10'h254 == _EVAL_5757;
  assign _EVAL_5646 = _EVAL_597 & _EVAL_847;
  assign _EVAL_658 = _EVAL_3225 & _EVAL_2301;
  assign _EVAL_693 = {1'h0,_EVAL_5479,_EVAL_1899};
  assign _EVAL_5000 = _EVAL_1159[15:8];
  assign _EVAL_2053 = {{1'd0}, _EVAL_1498};
  assign _EVAL_3144 = {_EVAL_3958,_EVAL_1610};
  assign _EVAL_5605 = 10'h20b == _EVAL_5757;
  assign _EVAL_3378 = _EVAL_3671 ? _EVAL_673 : _EVAL_5278;
  assign _EVAL_1583 = {{1'd0}, _EVAL_3793};
  assign _EVAL_1260 = 4'h8 | _EVAL_5180;
  assign _EVAL_3392 = {{6'd0}, _EVAL_2264};
  assign _EVAL_4356 = _EVAL_198 > _EVAL_1474;
  assign _EVAL_3537 = _EVAL_3499 & _EVAL_4477;
  assign _EVAL_5125 = _EVAL_3319 & _EVAL_673;
  assign _EVAL_1507 = _EVAL_4869 > _EVAL_872;
  assign _EVAL_4935 = {{1'd0}, _EVAL_3189};
  assign _EVAL_3059 = _EVAL_4749 ? _EVAL_1540 : _EVAL_5870;
  assign _EVAL_5522 = {1'h0,_EVAL_3450};
  assign _EVAL_1267 = {{6'd0}, _EVAL_2434};
  assign _EVAL_2776 = {1'h0,_EVAL_1670,_EVAL_3645};
  assign _EVAL_1367 = _EVAL_5010 & _EVAL_1937;
  assign _EVAL_5151 = _EVAL_1732 & _EVAL_673;
  assign _EVAL_4382 = _EVAL_2905 & _EVAL_1544;
  assign _EVAL_3939 = _EVAL_5096 & _EVAL_3154;
  assign _EVAL_3832 = {{6'd0}, _EVAL_5321};
  assign _EVAL_5758 = _EVAL_3681 & _EVAL_673;
  assign _EVAL_2880 = _EVAL_3591 ? _EVAL_673 : _EVAL_195;
  assign _EVAL_5270 = 2'h2 | _EVAL_1416;
  assign _EVAL_5526 = {1'h0,_EVAL_5735,_EVAL_2211};
  assign _EVAL_2439 = {{6'd0}, _EVAL_450};
  assign _EVAL_1537 = _EVAL_5615 & _EVAL_3043;
  assign _EVAL_6067 = Queue__EVAL[7:0];
  assign _EVAL_671 = _EVAL_5068[644];
  assign _EVAL_4178 = {_EVAL_4403,_EVAL_3172};
  assign _EVAL_3797 = {{6'd0}, _EVAL_3011};
  assign _EVAL_3790 = _EVAL_3088 ? _EVAL_2788 : _EVAL_5495;
  assign _EVAL_3343 = {{6'd0}, _EVAL_3120};
  assign _EVAL_1617 = {{6'd0}, _EVAL_2226};
  assign _EVAL_4860 = {1'h0,_EVAL_236,_EVAL_505};
  assign _EVAL_234 = _EVAL_5068[580];
  assign _EVAL_5746 = {1'h0,_EVAL_2339,_EVAL_2487};
  assign _EVAL_5191 = _EVAL_519 ? _EVAL_4285 : _EVAL_5097;
  assign _EVAL_3114 = 2'h2 | _EVAL_4638;
  assign _EVAL_1531 = _EVAL_427 ? 1'h0 : 1'h1;
  assign _EVAL_2618 = {{6'd0}, _EVAL_3494};
  assign _EVAL_6016 = {1'h0,_EVAL_5609,_EVAL_2094};
  assign _EVAL_3620 = _EVAL_1825 & _EVAL_417;
  assign _EVAL_2832 = {1'h0,_EVAL_4810,_EVAL_379};
  assign _EVAL_2521 = _EVAL_1753 & _EVAL_4477;
  assign _EVAL_229 = _EVAL_4828 & _EVAL_3384;
  assign _EVAL_2857 = _EVAL_1713 & _EVAL_673;
  assign _EVAL_5097 = _EVAL_4523 ? _EVAL_3392 : _EVAL_5140;
  assign _EVAL_3148 = {{6'd0}, _EVAL_2866};
  assign _EVAL_500 = _EVAL_5951 & _EVAL_676;
  assign _EVAL_4818 = {1'h0,_EVAL_4732};
  assign _EVAL_273 = {1'h0,_EVAL_5386,_EVAL_2681};
  assign _EVAL_4164 = _EVAL_1408 & _EVAL_3194;
  assign _EVAL_6027 = {{6'd0}, _EVAL_4508};
  assign _EVAL_1855 = {{6'd0}, _EVAL_4615};
  assign _EVAL_2610 = _EVAL_912 ? _EVAL_1785 : _EVAL_2752;
  assign _EVAL_683 = {1'h0,_EVAL_1293,_EVAL_4493};
  assign _EVAL_5501 = {1'h0,_EVAL_3152,_EVAL_6041};
  assign _EVAL_2343 = _EVAL_1235 & _EVAL_5696;
  assign _EVAL_5096 = _EVAL_384 & _EVAL_673;
  assign _EVAL_618 = _EVAL_2058 & _EVAL_1937;
  assign _EVAL_1556 = {1'h0,_EVAL_4738,_EVAL_2797};
  assign _EVAL_3027 = {{1'd0}, _EVAL_3703};
  assign _EVAL_5254 = _EVAL_1775[63:56];
  assign _EVAL_1969 = {{6'd0}, _EVAL_273};
  assign _EVAL_5806 = 10'h25b == _EVAL_5757;
  assign _EVAL_459 = {_EVAL_3980,_EVAL_5667};
  assign _EVAL_2884 = _EVAL_5068[669];
  assign _EVAL_898 = _EVAL_6066 > _EVAL_1998;
  assign _EVAL_226 = _EVAL_3093 ? 1'h0 : 1'h1;
  assign Queue__EVAL_3 = _EVAL_34;
  assign _EVAL_2596 = 10'h288 == _EVAL_5757;
  assign _EVAL_2566 = 10'h25a == _EVAL_5757;
  assign _EVAL_1091 = {{6'd0}, _EVAL_4818};
  assign _EVAL_466 = _EVAL_3731 ? _EVAL_4646 : _EVAL_2761;
  assign _EVAL_796 = _EVAL_4215 & _EVAL_673;
  assign _EVAL_3636 = _EVAL_762 & _EVAL_417;
  assign _EVAL_5817 = _EVAL_4448 ? _EVAL_1160 : _EVAL_5958;
  assign _EVAL_2303 = {1'h0,_EVAL_3203,_EVAL_1091};
  assign _EVAL_2141 = _EVAL_4308 & _EVAL_1131;
  assign _EVAL_5933 = _EVAL_3083 ? _EVAL_673 : _EVAL_2199;
  assign _EVAL_632 = _EVAL_2352 ? _EVAL_3275 : _EVAL_5824;
  assign _EVAL_4582 = _EVAL_2470 ? 1'h0 : 1'h1;
  assign _EVAL_5533 = {1'h0,_EVAL_5345,_EVAL_5861};
  assign _EVAL_4858 = _EVAL_4412 ? _EVAL_2751 : _EVAL_1023;
  assign _EVAL_5378 = {{6'd0}, _EVAL_2692};
  assign _EVAL_4153 = _EVAL_945 ? _EVAL_673 : _EVAL_3563;
  assign _EVAL_3477 = _EVAL_2227 > _EVAL_4973;
  assign _EVAL_3713 = {{6'd0}, _EVAL_1060};
  assign _EVAL_4848 = {{6'd0}, _EVAL_1496};
  assign _EVAL_6058 = _EVAL_1217 ? _EVAL_1249 : _EVAL_5844;
  assign _EVAL_3452 = _EVAL_2218[47:40];
  assign _EVAL_5617 = _EVAL_5545 > _EVAL_5373;
  assign _EVAL_5399 = 10'h21d == _EVAL_5757;
  assign _EVAL_2501 = {{6'd0}, _EVAL_5621};
  assign _EVAL_2996 = {{6'd0}, _EVAL_3715};
  assign _EVAL_1160 = {{6'd0}, _EVAL_2563};
  assign _EVAL_729 = _EVAL_1626 ? _EVAL_5220 : _EVAL_4229;
  assign _EVAL_2683 = _EVAL_3927 & _EVAL_673;
  assign _EVAL_3271 = {{6'd0}, _EVAL_5001};
  assign _EVAL_4699 = {_EVAL_3207,_EVAL_272};
  assign _EVAL_519 = 10'h221 == _EVAL_5757;
  assign _EVAL_1682 = _EVAL_1403 & _EVAL_2350;
  assign _EVAL_6064 = _EVAL_5951 & _EVAL_2515;
  assign _EVAL_1436 = _EVAL_3273 & _EVAL_673;
  assign _EVAL_5852 = _EVAL_3670 ? _EVAL_5660 : _EVAL_439;
  assign _EVAL_3320 = 3'h4 | _EVAL_5580;
  assign _EVAL_4252 = _EVAL_5951 & _EVAL_5637;
  assign _EVAL_2739 = {{1'd0}, _EVAL_1842};
  assign _EVAL_5070 = _EVAL_5951 & _EVAL_3365;
  assign _EVAL_304 = {1'h0,_EVAL_4843,_EVAL_3550};
  assign _EVAL_1608 = _EVAL_1002 & _EVAL_673;
  assign _EVAL_4117 = _EVAL_5052 & _EVAL_847;
  assign _EVAL_3298 = _EVAL_5068[587];
  assign _EVAL_3308 = _EVAL_5972 > _EVAL_4770;
  assign _EVAL_6013 = {_EVAL_5254,_EVAL_3504,_EVAL_545,_EVAL_851};
  assign _EVAL_293 = {1'h0,_EVAL_5315};
  assign _EVAL_2281 = _EVAL_5068[512];
  assign _EVAL_5802 = _EVAL_5758 & _EVAL_3487;
  assign _EVAL_185 = _EVAL_2197 ? _EVAL_673 : _EVAL_6012;
  assign _EVAL_2559 = {{1'd0}, _EVAL_4634};
  assign _EVAL_6071 = _EVAL_4014 & _EVAL_4932;
  assign _EVAL_881 = _EVAL_5951 & _EVAL_3502;
  assign _EVAL_4684 = _EVAL_2857 & _EVAL_3154;
  assign _EVAL_366 = {{6'd0}, _EVAL_5847};
  assign _EVAL_3643 = _EVAL_5995 ? _EVAL_5785 : _EVAL_5262;
  assign _EVAL_2741 = _EVAL_2621 & _EVAL_3487;
  assign _EVAL_1759 = {{6'd0}, _EVAL_3751};
  assign _EVAL_992 = _EVAL_3308 ? 1'h0 : 1'h1;
  assign _EVAL_3618 = _EVAL_1560 > _EVAL_903;
  assign _EVAL_2492 = Queue__EVAL[31:24];
  assign _EVAL_1002 = _EVAL_5951 & _EVAL_1464;
  assign _EVAL_1415 = _EVAL_3318 & _EVAL_3154;
  assign _EVAL_786 = _EVAL_5068[584];
  assign _EVAL_3483 = _EVAL_1507 ? {{1'd0}, _EVAL_305} : _EVAL_1114;
  assign _EVAL_2630 = _EVAL_3197 & _EVAL_1388;
  assign _EVAL_4846 = {1'h0,_EVAL_1311,_EVAL_1522};
  assign _EVAL_2914 = _EVAL_3887 & _EVAL_1331;
  assign _EVAL_4538 = {1'h0,_EVAL_3789,_EVAL_1760};
  assign _EVAL_4940 = _EVAL_1787 > _EVAL_4883;
  assign _EVAL_3900 = _EVAL_2190 ? _EVAL_673 : _EVAL_5965;
  assign _EVAL_6041 = {{6'd0}, _EVAL_3697};
  assign _EVAL_3087 = _EVAL_5432 & _EVAL_3154;
  assign _EVAL_4486 = _EVAL_3635 & _EVAL_673;
  assign _EVAL_2743 = _EVAL_4176 > _EVAL_632;
  assign _EVAL_1987 = {1'h0,_EVAL_4808,_EVAL_1473};
  assign _EVAL_2113 = {1'h0,_EVAL_666,_EVAL_593};
  assign _EVAL_3088 = _EVAL_2788 > _EVAL_5495;
  assign _EVAL_2764 = _EVAL_5792 ? _EVAL_673 : _EVAL_4136;
  assign _EVAL_450 = {1'h0,_EVAL_5309,_EVAL_2508};
  assign _EVAL_1575 = _EVAL_246 & _EVAL_2350;
  assign _EVAL_2332 = {_EVAL_1922,_EVAL_5727};
  assign _EVAL_1460 = {1'h0,_EVAL_3594};
  assign _EVAL_3925 = _EVAL_4740 > _EVAL_4776;
  assign _EVAL_5689 = {{6'd0}, _EVAL_250};
  assign _EVAL_4370 = _EVAL_5780 | _EVAL_3899;
  assign _EVAL_1860 = _EVAL_267 & _EVAL_673;
  assign _EVAL_1871 = _EVAL_5113 & _EVAL_1937;
  assign _EVAL_445 = _EVAL_4614 ? _EVAL_4603 : _EVAL_3380;
  assign _EVAL_1462 = _EVAL_3092 & _EVAL_2756;
  assign _EVAL_2964 = _EVAL_5363 ? _EVAL_2492 : _EVAL_5254;
  assign _EVAL_4496 = {1'h0,_EVAL_4828};
  assign _EVAL_6061 = _EVAL_4058 > _EVAL_2819;
  assign _EVAL_785 = 10'h28b == _EVAL_5757;
  assign _EVAL_276 = _EVAL_1668 ? _EVAL_5463 : _EVAL_4953;
  assign _EVAL_3892 = _EVAL_762 & _EVAL_1937;
  assign _EVAL_553 = _EVAL_4865 & _EVAL_4477;
  assign _EVAL_2661 = _EVAL_5068[611];
  assign _EVAL_569 = _EVAL_4978 ? _EVAL_1577 : _EVAL_3790;
  assign _EVAL_3502 = _EVAL_5068[649];
  assign _EVAL_3083 = 10'h0 == _EVAL_5757;
  assign _EVAL_1964 = {1'h0,_EVAL_4944,_EVAL_399};
  assign _EVAL_810 = _EVAL_511 & _EVAL_3487;
  assign _EVAL_4169 = {_EVAL_3434,_EVAL_1442};
  assign _EVAL_874 = _EVAL_5758 & _EVAL_3154;
  assign _EVAL_4242 = _EVAL_4865 & _EVAL_3487;
  assign _EVAL_4621 = _EVAL_2883 > _EVAL_405;
  assign _EVAL_4497 = _EVAL_5815 ? {{1'd0}, _EVAL_5375} : _EVAL_1222;
  assign _EVAL_2396 = {1'h0,_EVAL_5635,24'h0};
  assign _EVAL_68 = Queue__EVAL_0;
  assign _EVAL_4510 = _EVAL_1286 == 8'h0;
  assign _EVAL_2600 = {{6'd0}, _EVAL_5410};
  assign _EVAL_4897 = {1'h0,_EVAL_616,_EVAL_2641};
  assign _EVAL_3158 = _EVAL_4556 & _EVAL_1937;
  assign _EVAL_3115 = {{6'd0}, _EVAL_3357};
  assign _EVAL_4517 = _EVAL_4356 ? 1'h0 : 1'h1;
  assign _EVAL_5691 = {1'h0,_EVAL_2988};
  assign _EVAL_432 = _EVAL_519 ? _EVAL_673 : _EVAL_1683;
  assign _EVAL_2820 = _EVAL_4746 ? {{1'd0}, _EVAL_1829} : _EVAL_2004;
  assign _EVAL_4440 = _EVAL_3152 & _EVAL_4087;
  assign _EVAL_5865 = {{6'd0}, _EVAL_3022};
  assign _EVAL_1998 = _EVAL_3765 ? _EVAL_720 : _EVAL_2869;
  assign _EVAL_5540 = _EVAL_2372 & _EVAL_673;
  assign _EVAL_325 = Queue__EVAL_8 & 22'h1fecc0;
  assign _EVAL_863 = {_EVAL_624,_EVAL_1351};
  assign _EVAL_4199 = 10'h293 == _EVAL_5757;
  assign _EVAL_2660 = _EVAL_3339 & _EVAL_4477;
  assign _EVAL_5520 = Queue__EVAL_8[9];
  assign _EVAL_5335 = _EVAL_3851 > _EVAL_5480;
  assign _EVAL_1788 = _EVAL_3454 > _EVAL_5227;
  assign _EVAL_495 = _EVAL_3344 ? _EVAL_5579 : _EVAL_4864;
  assign _EVAL_5330 = _EVAL_1609 > _EVAL_664;
  assign _EVAL_1247 = _EVAL_5147 & _EVAL_2837;
  assign _EVAL_4865 = _EVAL_1377 & _EVAL_673;
  assign _EVAL_2936 = _EVAL_1119 > _EVAL_5925;
  assign _EVAL_4296 = {{6'd0}, _EVAL_2832};
  assign _EVAL_762 = _EVAL_1704 & _EVAL_673;
  assign _EVAL_1454 = _EVAL_2474 & _EVAL_417;
  assign _EVAL_1379 = {1'h0,_EVAL_3847,_EVAL_2415};
  assign _EVAL_1417 = 4'h8 | _EVAL_1872;
  assign _EVAL_2541 = _EVAL_1770 ? _EVAL_673 : _EVAL_1410;
  assign _EVAL_4774 = {1'h0,_EVAL_4051,_EVAL_833};
  assign _EVAL_4716 = _EVAL_5636 ? _EVAL_3713 : _EVAL_5901;
  assign _EVAL_4388 = 7'h40 | _EVAL_4070;
  assign _EVAL_3030 = _EVAL_2701 & _EVAL_417;
  assign _EVAL_1825 = _EVAL_5382 & _EVAL_673;
  assign _EVAL_2935 = _EVAL_2474 & _EVAL_2350;
  assign _EVAL_4067 = _EVAL_988 ? _EVAL_673 : _EVAL_4704;
  assign _EVAL_3017 = {1'h0,_EVAL_3384,24'h0};
  assign _EVAL_2138 = 2'h2 | _EVAL_2276;
  assign _EVAL_1766 = _EVAL_3670 ? _EVAL_673 : _EVAL_4032;
  assign _EVAL_5295 = {{6'd0}, _EVAL_4660};
  assign _EVAL_2473 = 10'h245 == _EVAL_5757;
  assign _EVAL_3937 = {_EVAL_1117,_EVAL_2781};
  assign _EVAL_3022 = {1'h0,_EVAL_3843,_EVAL_3024};
  assign _EVAL_2147 = _EVAL_163 ? _EVAL_1930 : _EVAL_4659;
  assign _EVAL_991 = {1'h0,_EVAL_1645,_EVAL_1855};
  assign _EVAL_5935 = _EVAL_2261 > _EVAL_1457;
  assign _EVAL_166 = _EVAL_1775[23:16];
  assign _EVAL_4469 = 10'h291 == _EVAL_5757;
  assign _EVAL_3665 = 10'h296 == _EVAL_5757;
  assign _EVAL_844 = _EVAL_1378 & _EVAL_417;
  assign _EVAL_2261 = {_EVAL_4500,_EVAL_5713};
  assign _EVAL_575 = {{6'd0}, _EVAL_3567};
  assign _EVAL_5394 = {1'h0,_EVAL_1929,_EVAL_2547};
  assign _EVAL_2800 = _EVAL_4199 ? _EVAL_673 : _EVAL_4009;
  assign _EVAL_215 = _EVAL_3498 ? _EVAL_673 : _EVAL_4849;
  assign _EVAL_5007 = _EVAL_5681 > _EVAL_4717;
  assign _EVAL_5364 = _EVAL_1507 ? _EVAL_4869 : _EVAL_872;
  assign _EVAL_3590 = _EVAL_5511 & _EVAL_3154;
  assign _EVAL_427 = _EVAL_5165 > _EVAL_2228;
  assign _EVAL_1263 = {1'h0,_EVAL_487,_EVAL_4852};
  assign _EVAL_3024 = {{6'd0}, _EVAL_2463};
  assign _EVAL_1908 = _EVAL_4331 ? 1'h0 : 1'h1;
  assign _EVAL_3980 = _EVAL_1593 & _EVAL_4808;
  assign _EVAL_3521 = _EVAL_1112 | _EVAL_2406;
  assign _EVAL_4970 = _EVAL_5951 & _EVAL_671;
  assign _EVAL_3053 = _EVAL_4612 & _EVAL_1166;
  assign _EVAL_5993 = _EVAL_5540 & _EVAL_2350;
  assign _EVAL_3533 = _EVAL_333 ? _EVAL_673 : _EVAL_2398;
  assign _EVAL_4953 = _EVAL_4244 ? _EVAL_4274 : _EVAL_5555;
  assign _EVAL_5257 = {1'h0,_EVAL_2312,_EVAL_6027};
  assign _EVAL_1481 = {1'h0,_EVAL_880,_EVAL_1597};
  assign _EVAL_743 = _EVAL_930 ? _EVAL_1517 : _EVAL_3823;
  assign _EVAL_1934 = _EVAL_5010 & _EVAL_417;
  assign _EVAL_2248 = _EVAL_3662 ? _EVAL_2780 : _EVAL_3666;
  assign _EVAL_977 = {{6'd0}, _EVAL_436};
  assign _EVAL_3290 = _EVAL_1040 & _EVAL_2381;
  assign _EVAL_1927 = {{6'd0}, _EVAL_1181};
  assign _EVAL_5883 = 10'h257 == _EVAL_5757;
  assign _EVAL_4534 = _EVAL_3786 ? {{1'd0}, _EVAL_3762} : _EVAL_2591;
  assign _EVAL_5183 = _EVAL_5683 ? _EVAL_995 : _EVAL_4354;
  assign _EVAL_1805 = _EVAL_3477 ? 1'h0 : 1'h1;
  assign _EVAL_3499 = _EVAL_3668 & _EVAL_673;
  assign _EVAL_514 = _EVAL_3391 ? _EVAL_6067 : _EVAL_1282;
  assign _EVAL_2633 = _EVAL_3278 & _EVAL_673;
  assign _EVAL_3696 = {{1'd0}, _EVAL_4600};
  assign _EVAL_5204 = _EVAL_2342 ? {{1'd0}, _EVAL_4170} : _EVAL_1304;
  assign _EVAL_5830 = _EVAL_3372 ? {{1'd0}, _EVAL_1492} : _EVAL_1265;
  assign _EVAL_4539 = _EVAL_5995 ? _EVAL_673 : _EVAL_3442;
  assign _EVAL_4809 = _EVAL_2824 > _EVAL_3353;
  assign _EVAL_3819 = _EVAL_3905 ? 3'h3 : _EVAL_4658;
  assign _EVAL_368 = {_EVAL_893,_EVAL_4711};
  assign _EVAL_2815 = _EVAL_3609 & _EVAL_5479;
  assign _EVAL_628 = _EVAL_3339 & _EVAL_3154;
  assign _EVAL_4990 = _EVAL_4318 ? {{1'd0}, _EVAL_4958} : _EVAL_4388;
  assign _EVAL_423 = _EVAL_5951 & _EVAL_2898;
  assign _EVAL_1129 = _EVAL_1502 ? {{1'd0}, _EVAL_3573} : _EVAL_3320;
  assign _EVAL_2794 = {{6'd0}, _EVAL_1883};
  assign _EVAL_1249 = {_EVAL_542,4'hf,_EVAL_994,4'hf,_EVAL_5623,4'hf,_EVAL_2493,4'hf};
  assign _EVAL_5481 = _EVAL_3989 & _EVAL_847;
  assign _EVAL_5064 = _EVAL_500 & _EVAL_673;
  assign _EVAL_2353 = {1'h0,_EVAL_3866,_EVAL_1690};
  assign _EVAL_4633 = _EVAL_5873 ? _EVAL_5807 : _EVAL_5166;
  assign _EVAL_924 = {1'h0,1'h0,_EVAL_291};
  assign _EVAL_4876 = _EVAL_5609 & _EVAL_896;
  assign _EVAL_1674 = _EVAL_5989 | _EVAL_4515;
  assign _EVAL_2756 = _EVAL_4213 == 4'hf;
  assign _EVAL_2185 = 3'h4 | _EVAL_1898;
  assign _EVAL_353 = _EVAL_6035 ? _EVAL_673 : _EVAL_5062;
  assign _EVAL_2146 = _EVAL_1621 ? _EVAL_1337 : _EVAL_3654;
  assign _EVAL_4508 = {1'h0,_EVAL_5743,_EVAL_5718};
  assign _EVAL_3283 = _EVAL_1956 & _EVAL_673;
  assign _EVAL_3507 = _EVAL_785 ? _EVAL_5436 : _EVAL_2944;
  assign _EVAL_2092 = 10'h252 == _EVAL_5757;
  assign _EVAL_2883 = {_EVAL_5391,_EVAL_3538};
  assign _EVAL_912 = _EVAL_1785 > _EVAL_2752;
  assign _EVAL_3397 = _EVAL_3750 > _EVAL_495;
  assign _EVAL_5391 = _EVAL_891 & _EVAL_5232;
  assign _EVAL_5718 = {{6'd0}, _EVAL_293};
  assign _EVAL_1345 = {{6'd0}, _EVAL_2017};
  assign _EVAL_4606 = _EVAL_2787 > _EVAL_5325;
  assign _EVAL_3911 = _EVAL_516 & _EVAL_3154;
  assign _EVAL_5041 = _EVAL_6052 & _EVAL_3154;
  assign _EVAL_5799 = _EVAL_2050 ? _EVAL_673 : _EVAL_1219;
  assign _EVAL_5580 = {{1'd0}, _EVAL_1128};
  assign _EVAL_1140 = 10'h255 == _EVAL_5757;
  assign _EVAL_3253 = _EVAL_2092 ? _EVAL_673 : _EVAL_4894;
  assign _EVAL_5582 = _EVAL_5068[607];
  assign _EVAL_2774 = {_EVAL_6101,_EVAL_2984};
  assign _EVAL_3019 = {1'h0,_EVAL_4779,_EVAL_2989};
  assign _EVAL_2711 = _EVAL_3171 & _EVAL_3129;
  assign _EVAL_5714 = {1'h0,_EVAL_2669,_EVAL_5197};
  assign _EVAL_4229 = _EVAL_5007 ? _EVAL_5681 : _EVAL_4717;
  assign _EVAL_6043 = _EVAL_5758 & _EVAL_4477;
  assign _EVAL_2385 = _EVAL_4948 ? _EVAL_4089 : _EVAL_5263;
  assign _EVAL_4307 = {1'h0,_EVAL_1342,_EVAL_1204};
  assign _EVAL_5154 = _EVAL_3283 & _EVAL_1937;
  assign _EVAL_2265 = _EVAL_3339 & _EVAL_3487;
  assign _EVAL_1504 = {_EVAL_1247,_EVAL_1052};
  assign _EVAL_2623 = {1'h0,_EVAL_1166,_EVAL_1190};
  assign _EVAL_3877 = {_EVAL_5881,_EVAL_412};
  assign _EVAL_142 = Queue__EVAL_14;
  assign _EVAL_4709 = Queue__EVAL[23:20];
  assign _EVAL_812 = _EVAL_1504 > _EVAL_5996;
  assign _EVAL_3831 = _EVAL_5314 & _EVAL_3487;
  assign _EVAL_2182 = _EVAL_1626 ? {{1'd0}, _EVAL_5585} : _EVAL_5312;
  assign _EVAL_999 = {1'h0,_EVAL_1664,_EVAL_178};
  assign _EVAL_2351 = 10'h218 == _EVAL_5757;
  assign _EVAL_489 = _EVAL_1860 & _EVAL_4477;
  assign _EVAL_5475 = Queue__EVAL_8[21];
  assign _EVAL_3685 = _EVAL_1502 ? _EVAL_3270 : _EVAL_5231;
  assign _EVAL_3805 = _EVAL_5068[257];
  assign _EVAL_1771 = {{6'd0}, _EVAL_4538};
  assign _EVAL_2928 = _EVAL_2979 ? {{1'd0}, _EVAL_3309} : _EVAL_3335;
  assign _EVAL_1592 = _EVAL_5821 & _EVAL_4477;
  assign _EVAL_4238 = {1'h0,_EVAL_4348,_EVAL_3463};
  assign _EVAL_4553 = 10'h217 == _EVAL_5757;
  assign _EVAL_198 = {_EVAL_3169,_EVAL_3767};
  assign _EVAL_2547 = {{6'd0}, _EVAL_5137};
  assign _EVAL_5506 = _EVAL_1917 & _EVAL_2669;
  assign _EVAL_2722 = {1'h0,_EVAL_2162,_EVAL_5377};
  assign _EVAL_3753 = _EVAL_2009 & _EVAL_5101;
  assign _EVAL_4933 = {{6'd0}, _EVAL_4400};
  assign _EVAL_2036 = 10'h206 == _EVAL_5757;
  assign _EVAL_1866 = _EVAL_1074 > _EVAL_6100;
  assign _EVAL_1059 = _EVAL_2444 & _EVAL_4119;
  assign _EVAL_2523 = _EVAL_6053 & _EVAL_2756;
  assign _EVAL_4595 = {{1'd0}, _EVAL_4880};
  assign _EVAL_4882 = _EVAL_1314 & _EVAL_507;
  assign _EVAL_5436 = {_EVAL_4997,4'hf,_EVAL_4040,4'hf,_EVAL_2561,4'hf,_EVAL_2806,4'hf};
  assign _EVAL_438 = {_EVAL_899,4'hf,_EVAL_1629,4'hf,_EVAL_1882,4'hf,_EVAL_2293,4'hf};
  assign _EVAL_2503 = _EVAL_5684 & _EVAL_1510;
  assign _EVAL_189 = _EVAL_343 ? _EVAL_2636 : _EVAL_5334;
  assign _EVAL_1138 = _EVAL_5951 & _EVAL_2864;
  assign _EVAL_4128 = _EVAL_2128 ? 1'h0 : 1'h1;
  assign _EVAL_5332 = _EVAL_2703 ? _EVAL_673 : _EVAL_2691;
  assign _EVAL_2119 = _EVAL_1075 & _EVAL_417;
  assign _EVAL_2862 = _EVAL_4511 > _EVAL_3430;
  assign _EVAL_3666 = _EVAL_3597 ? _EVAL_5004 : _EVAL_567;
  assign _EVAL_2101 = 10'h240 == _EVAL_5757;
  assign _EVAL_3675 = _EVAL_2034 ? _EVAL_673 : _EVAL_2933;
  assign _EVAL_295 = _EVAL_5045 ? _EVAL_5803 : _EVAL_1284;
  assign _EVAL_437 = {1'h0,_EVAL_2065,_EVAL_3682};
  assign _EVAL_3475 = _EVAL_2247 & _EVAL_3286;
  assign _EVAL_4354 = _EVAL_270 ? _EVAL_1812 : _EVAL_1983;
  assign _EVAL_3044 = _EVAL_3986 & _EVAL_355;
  assign _EVAL_4797 = _EVAL_4653 & _EVAL_3154;
  assign _EVAL_3146 = 10'h204 == _EVAL_5757;
  assign _EVAL_4665 = _EVAL_4337 ? _EVAL_2501 : _EVAL_5095;
  assign _EVAL_3709 = Queue__EVAL[31:28];
  assign _EVAL_5384 = _EVAL_5605 ? _EVAL_3947 : _EVAL_3643;
  assign _EVAL_4820 = _EVAL_2467 > _EVAL_1354;
  assign _EVAL_420 = {{1'd0}, _EVAL_4050};
  assign _EVAL_3674 = _EVAL_1775[15:8];
  assign _EVAL_1497 = {{6'd0}, _EVAL_5487};
  assign _EVAL_211 = {{6'd0}, _EVAL_5710};
  assign _EVAL_5709 = {{6'd0}, _EVAL_3975};
  assign _EVAL_6035 = 10'h24c == _EVAL_5757;
  assign _EVAL_5392 = {1'h0,_EVAL_4785,_EVAL_2158};
  assign _EVAL_4213 = _EVAL_1159[31:28];
  assign _EVAL_5657 = _EVAL_2229 & _EVAL_1777;
  assign _EVAL_3086 = _EVAL_2351 ? _EVAL_673 : _EVAL_4153;
  assign _EVAL_2486 = _EVAL_636 & _EVAL_673;
  assign _EVAL_3385 = {4'h0,_EVAL_4679};
  assign _EVAL_5770 = _EVAL_5960 ? _EVAL_1572 : _EVAL_1335;
  assign _EVAL_3266 = _EVAL_2595 & _EVAL_2350;
  assign _EVAL_264 = {1'h0,_EVAL_5675,24'h0};
  assign _EVAL_488 = _EVAL_3215 & _EVAL_2350;
  assign _EVAL_5499 = {{6'd0}, _EVAL_1963};
  assign _EVAL_5287 = _EVAL_879 ? _EVAL_3102 : _EVAL_681;
  assign _EVAL_3653 = {{6'd0}, _EVAL_5181};
  assign _EVAL_2168 = _EVAL_516 & _EVAL_4477;
  assign _EVAL_5539 = _EVAL_2621 & _EVAL_847;
  assign _EVAL_3960 = _EVAL_1018 ? _EVAL_980 : {{8'd0}, _EVAL_2579};
  assign _EVAL_5312 = 2'h2 | _EVAL_655;
  assign _EVAL_1128 = _EVAL_5145 ? {{1'd0}, _EVAL_3839} : _EVAL_840;
  assign _EVAL_647 = {_EVAL_3753,_EVAL_5765};
  assign _EVAL_526 = {{6'd0}, _EVAL_4425};
  assign _EVAL_1930 = {{6'd0}, _EVAL_4081};
  assign _EVAL_5851 = _EVAL_6049 & _EVAL_4477;
  assign _EVAL_3958 = _EVAL_5890 & _EVAL_2847;
  assign _EVAL_3929 = _EVAL_823 ? {{1'd0}, _EVAL_5571} : _EVAL_3114;
  assign _EVAL_3846 = {{6'd0}, _EVAL_3570};
  assign _EVAL_270 = _EVAL_1812 > _EVAL_1983;
  assign _EVAL_2282 = {{6'd0}, _EVAL_5849};
  assign Queue__EVAL_15 = _EVAL_140;
  assign _EVAL_763 = {_EVAL_6014,_EVAL_994};
  assign _EVAL_2801 = {{6'd0}, _EVAL_5550};
  assign _EVAL_2639 = {{1'd0}, _EVAL_5830};
  assign _EVAL_1823 = {1'h0,_EVAL_1331,_EVAL_5731};
  assign _EVAL_611 = _EVAL_5951 & _EVAL_1093;
  assign _EVAL_305 = _EVAL_2104 ? {{1'd0}, _EVAL_274} : _EVAL_1260;
  assign _EVAL_5563 = _EVAL_2286 ? _EVAL_673 : _EVAL_5799;
  assign _EVAL_1519 = {{6'd0}, _EVAL_3915};
  assign _EVAL_3836 = {{4'd0}, _EVAL_1280};
  assign _EVAL_5621 = {1'h0,_EVAL_1245,_EVAL_2010};
  assign _EVAL_1898 = {{1'd0}, _EVAL_502};
  assign _EVAL_1753 = _EVAL_485 & _EVAL_673;
  assign _EVAL_3359 = {{6'd0}, _EVAL_683};
  assign _EVAL_2922 = _EVAL_1806 & _EVAL_4477;
  assign _EVAL_4321 = 2'h2 | _EVAL_2429;
  assign _EVAL_1323 = _EVAL_2225 | _EVAL_2714;
  assign _EVAL_4602 = ~Queue__EVAL_2;
  assign _EVAL_1597 = {{6'd0}, _EVAL_5407};
  assign _EVAL_4402 = 10'h207 == _EVAL_5757;
  assign _EVAL_86 = _EVAL_1286;
  assign _EVAL_2520 = _EVAL_5068[656];
  assign _EVAL_4599 = _EVAL_4080 & _EVAL_5535;
  assign _EVAL_1469 = {_EVAL_3345,_EVAL_2490};
  assign _EVAL_411 = _EVAL_2406 ? _EVAL_1035 : _EVAL_3504;
  assign _EVAL_401 = {{6'd0}, _EVAL_3971};
  assign _EVAL_527 = _EVAL_6049 & _EVAL_3154;
  assign _EVAL_657 = {1'h0,_EVAL_3609,_EVAL_1232};
  assign _EVAL_5983 = _EVAL_1423 ? 1'h0 : 1'h1;
  assign _EVAL_2971 = {1'h0,_EVAL_1544};
  assign _EVAL_2022 = _EVAL_4486 & _EVAL_2350;
  assign _EVAL_246 = _EVAL_1659 & _EVAL_673;
  assign _EVAL_1264 = _EVAL_2862 ? {{1'd0}, _EVAL_2838} : _EVAL_522;
  assign _EVAL_15 = _EVAL_4510 ? 8'h0 : _EVAL_3190;
  assign _EVAL_3358 = _EVAL_2701 & _EVAL_2350;
  assign _EVAL_5791 = _EVAL_3067 > _EVAL_1120;
  assign _EVAL_1255 = _EVAL_3363 & _EVAL_3962;
  assign _EVAL_384 = _EVAL_5951 & _EVAL_5997;
  assign _EVAL_6081 = _EVAL_5928 & _EVAL_417;
  assign _EVAL_4540 = _EVAL_1788 ? _EVAL_3454 : _EVAL_5227;
  assign _EVAL_3518 = _EVAL_5049 ? _EVAL_919 : _EVAL_4816;
  assign _EVAL_5117 = _EVAL_4778 ? _EVAL_5689 : _EVAL_2535;
  assign _EVAL_851 = _EVAL_1775[39:32];
  assign _EVAL_4687 = _EVAL_4672 ? {{1'd0}, _EVAL_2182} : _EVAL_2185;
  assign _EVAL_1937 = _EVAL_3427 == 4'hf;
  assign _EVAL_4954 = {{6'd0}, _EVAL_3098};
  assign _EVAL_5403 = _EVAL_1656 ? 1'h0 : 1'h1;
  assign _EVAL_1018 = 10'h2a2 == _EVAL_5757;
  assign _EVAL_4483 = {_EVAL_3739,_EVAL_702};
  assign _EVAL_425 = {{1'd0}, _EVAL_4262};
  assign _EVAL_1437 = _EVAL_368 > _EVAL_5098;
  assign _EVAL_2530 = _EVAL_1753 & _EVAL_3487;
  assign _EVAL_815 = {{6'd0}, _EVAL_4195};
  assign _EVAL_5195 = _EVAL_5511 & _EVAL_4477;
  assign _EVAL_2178 = {{6'd0}, _EVAL_3871};
  assign _EVAL_502 = _EVAL_1903 ? {{1'd0}, _EVAL_1218} : _EVAL_4677;
  assign _EVAL_3309 = _EVAL_5120 ? {{1'd0}, _EVAL_1748} : _EVAL_3096;
  assign _EVAL_2091 = _EVAL_2728 & _EVAL_4247;
  assign _EVAL_1851 = _EVAL_5540 & _EVAL_1937;
  assign _EVAL_1740 = {{6'd0}, _EVAL_5687};
  assign _EVAL_5052 = _EVAL_742 & _EVAL_673;
  assign _EVAL_2869 = _EVAL_2862 ? _EVAL_4511 : _EVAL_3430;
  assign _EVAL_934 = _EVAL_5468 & _EVAL_2350;
  assign _EVAL_5547 = _EVAL_5935 ? _EVAL_2261 : _EVAL_1457;
  assign _EVAL_3380 = {_EVAL_760,_EVAL_5624};
  assign _EVAL_913 = _EVAL_4785 & _EVAL_1880;
  assign _EVAL_4313 = {{6'd0}, _EVAL_5061};
  assign _EVAL_5763 = _EVAL_4142 ? _EVAL_2146 : _EVAL_5322;
  assign _EVAL_2276 = {{1'd0}, _EVAL_4747};
  assign _EVAL_5669 = {1'h0,1'h0,_EVAL_4982};
  assign _EVAL_2681 = {{6'd0}, _EVAL_979};
  assign _EVAL_2595 = _EVAL_2322 & _EVAL_673;
  assign _EVAL_1357 = 2'h2 | _EVAL_3625;
  assign _EVAL_2024 = {_EVAL_3464,4'hf,_EVAL_1610,4'hf,_EVAL_5981,4'hf,_EVAL_2827,4'hf};
  assign _EVAL_2760 = _EVAL_727 & _EVAL_3133;
  assign _EVAL_2143 = _EVAL_2703 ? _EVAL_3359 : _EVAL_1632;
  assign _EVAL_1959 = _EVAL_5519 ? 8'hff : 8'h0;
  assign _EVAL_414 = _EVAL_945 ? _EVAL_401 : _EVAL_5453;
  assign _EVAL_2410 = {1'h0,_EVAL_3280,_EVAL_5908};
  assign _EVAL_5227 = {_EVAL_3999,_EVAL_1882};
  assign _EVAL_923 = _EVAL_5068[578];
  assign _EVAL_2108 = _EVAL_2954 & _EVAL_847;
  assign _EVAL_4520 = _EVAL_1030 ? _EVAL_294 : _EVAL_3578;
  assign _EVAL_3999 = _EVAL_4085 & _EVAL_3634;
  assign _EVAL_5694 = {{6'd0}, _EVAL_5808};
  assign _EVAL_5202 = 4'h8 - _EVAL_1746;
  assign _EVAL_3800 = _EVAL_4553 ? _EVAL_2491 : _EVAL_5863;
  assign _EVAL_5661 = _EVAL_1903 ? _EVAL_1472 : _EVAL_3997;
  assign _EVAL_3513 = _EVAL_5007 ? 1'h0 : 1'h1;
  assign _EVAL_2755 = _EVAL_2481 & _EVAL_847;
  assign _EVAL_5326 = _EVAL_2380 & _EVAL_3154;
  assign _EVAL_3654 = _EVAL_4940 ? _EVAL_1787 : _EVAL_4883;
  assign _EVAL_2855 = _EVAL_733 > _EVAL_647;
  assign _EVAL_1666 = _EVAL_3339 & _EVAL_847;
  assign _EVAL_747 = _EVAL_5068[641];
  assign _EVAL_2461 = _EVAL_1153 ? _EVAL_673 : _EVAL_3872;
  assign _EVAL_6073 = _EVAL_5787 & _EVAL_673;
  assign _EVAL_4449 = _EVAL_1403 & _EVAL_417;
  assign _EVAL_336 = _EVAL_5951 & _EVAL_1665;
  assign _EVAL_4721 = _EVAL_3521 | _EVAL_5363;
  assign _EVAL_1336 = _EVAL_5674 ? _EVAL_901 : _EVAL_1534;
  assign _EVAL_4969 = {1'h0,_EVAL_1121,_EVAL_741};
  assign _EVAL_3526 = {_EVAL_406,_EVAL_542};
  assign _EVAL_3390 = _EVAL_5615 & _EVAL_1292;
  assign _EVAL_5318 = {{6'd0}, _EVAL_5714};
  assign _EVAL_678 = _EVAL_597 & _EVAL_4477;
  assign _EVAL_3667 = _EVAL_1140 ? _EVAL_673 : _EVAL_2943;
  assign _EVAL_3930 = _EVAL_5883 ? _EVAL_2874 : _EVAL_6006;
  assign _EVAL_2692 = {1'h0,_EVAL_5307};
  assign _EVAL_3211 = _EVAL_5068[605];
  assign _EVAL_5698 = {{6'd0}, _EVAL_2303};
  assign _EVAL_636 = _EVAL_5951 & _EVAL_5711;
  assign _EVAL_3219 = _EVAL_3372 ? _EVAL_642 : _EVAL_466;
  assign _EVAL_4274 = _EVAL_898 ? _EVAL_6066 : _EVAL_1998;
  assign _EVAL_5731 = {{6'd0}, _EVAL_598};
  assign _EVAL_5925 = _EVAL_5791 ? _EVAL_3067 : _EVAL_1120;
  assign _EVAL_2489 = _EVAL_3499 & _EVAL_3154;
  assign _EVAL_3605 = _EVAL_5275 ? _EVAL_3576 : _EVAL_4799;
  assign _EVAL_2967 = {_EVAL_2392,_EVAL_4304};
  assign _EVAL_4569 = {{6'd0}, _EVAL_2767};
  assign _EVAL_3100 = _EVAL_5951 & _EVAL_2176;
  assign _EVAL_3612 = {1'h0,_EVAL_3327};
  assign _EVAL_3573 = _EVAL_3798 ? {{1'd0}, _EVAL_3627} : _EVAL_1390;
  assign _EVAL_6020 = {1'h0,_EVAL_4367,_EVAL_497};
  assign _EVAL_4772 = 10'h261 == _EVAL_5757;
  assign _EVAL_18 = Queue__EVAL_9;
  assign _EVAL_4615 = {1'h0,_EVAL_1618,_EVAL_3950};
  assign _EVAL_980 = {_EVAL_3743,4'hf,_EVAL_5667,4'hf,_EVAL_1440,4'hf,_EVAL_3467,4'hf};
  assign _EVAL_285 = {_EVAL_4068,_EVAL_1676};
  assign _EVAL_1298 = 4'h8 | _EVAL_4484;
  assign _EVAL_1476 = _EVAL_4562 ? _EVAL_673 : _EVAL_4284;
  assign _EVAL_5176 = {{6'd0}, _EVAL_1263};
  assign _EVAL_399 = {{6'd0}, _EVAL_4972};
  assign _EVAL_3737 = _EVAL_3989 & _EVAL_3487;
  assign _EVAL_5046 = _EVAL_2616 & _EVAL_1670;
  assign _EVAL_981 = {{4'd0}, _EVAL_4824};
  assign _EVAL_691 = _EVAL_5644 & _EVAL_3487;
  assign _EVAL_4683 = _EVAL_846 ? 1'h0 : 1'h1;
  assign _EVAL_1477 = _EVAL_3544 & _EVAL_673;
  assign _EVAL_597 = _EVAL_1438 & _EVAL_673;
  assign _EVAL_2622 = _EVAL_5222 & _EVAL_1937;
  assign _EVAL_1550 = {{6'd0}, _EVAL_4941};
  assign _EVAL_571 = _EVAL_597 & _EVAL_3487;
  assign _EVAL_1422 = {{6'd0}, _EVAL_447};
  assign _EVAL_182 = {{6'd0}, _EVAL_2854};
  assign _EVAL_2017 = {1'h0,_EVAL_1942};
  assign _EVAL_3036 = _EVAL_3391 | _EVAL_2063;
  assign _EVAL_3104 = _EVAL_4865 & _EVAL_847;
  assign _EVAL_4662 = _EVAL_2486 & _EVAL_417;
  assign _EVAL_3989 = _EVAL_3140 & _EVAL_673;
  assign _EVAL_1024 = _EVAL_2484 & _EVAL_4233;
  assign _EVAL_2283 = {1'h0,_EVAL_4922,_EVAL_2940};
  assign _EVAL_2980 = Queue__EVAL_4[2];
  assign _EVAL_5894 = _EVAL_6049 & _EVAL_3487;
  assign _EVAL_3705 = _EVAL_1753 & _EVAL_847;
  assign _EVAL_1282 = _EVAL_1775[7:0];
  assign _EVAL_2638 = _EVAL_3144 > _EVAL_4026;
  assign _EVAL_4541 = {1'h0,_EVAL_3363};
  assign _EVAL_5908 = {{6'd0}, _EVAL_667};
  assign _EVAL_676 = _EVAL_5068[673];
  assign _EVAL_261 = _EVAL_3099 ? _EVAL_5442 : _EVAL_2802;
  assign _EVAL_5829 = _EVAL_5068[652];
  assign _EVAL_893 = _EVAL_2154 & _EVAL_3374;
  assign _EVAL_2887 = 2'h2 | _EVAL_1306;
  assign _EVAL_4368 = {{6'd0}, _EVAL_766};
  assign _EVAL_5467 = {{6'd0}, _EVAL_5691};
  assign _EVAL_5107 = _EVAL_2063 ? _EVAL_3102 : _EVAL_3674;
  assign _EVAL_2605 = _EVAL_3092 & _EVAL_417;
  assign _EVAL_5366 = 2'h2 | _EVAL_2109;
  assign _EVAL_3748 = _EVAL_2784 & _EVAL_1937;
  assign _EVAL_1431 = _EVAL_5951 & _EVAL_5203;
  assign _EVAL_1075 = _EVAL_5898 & _EVAL_673;
  assign _EVAL_2164 = {_EVAL_5765,4'hf,_EVAL_2537,4'hf,_EVAL_3771,4'hf,_EVAL_834,4'hf};
  assign _EVAL_1177 = {1'h0,_EVAL_2148,_EVAL_5865};
  assign _EVAL_4349 = _EVAL_4250 ? _EVAL_673 : _EVAL_5611;
  assign _EVAL_382 = {{6'd0}, _EVAL_2777};
  assign _EVAL_3217 = _EVAL_5951 & _EVAL_5266;
  assign _EVAL_439 = _EVAL_2316 ? {{8'd0}, _EVAL_5963} : _EVAL_958;
  assign _EVAL_4659 = _EVAL_5048 ? _EVAL_173 : _EVAL_1698;
  assign _EVAL_2048 = _EVAL_3921 ? _EVAL_673 : _EVAL_6056;
  assign _EVAL_5156 = {{6'd0}, _EVAL_1172};
  assign _EVAL_6000 = _EVAL_3665 ? _EVAL_673 : _EVAL_3080;
  assign _EVAL_1445 = {1'h0,_EVAL_1040,_EVAL_716};
  assign _EVAL_4636 = _EVAL_1032 ? _EVAL_3191 : _EVAL_2115;
  assign _EVAL_1433 = {{1'd0}, _EVAL_3555};
  assign _EVAL_1704 = _EVAL_5951 & _EVAL_5829;
  assign _EVAL_1225 = _EVAL_5432 & _EVAL_3487;
  assign _EVAL_4869 = _EVAL_2104 ? _EVAL_5763 : _EVAL_4913;
  assign _EVAL_289 = _EVAL_5068[588];
  assign _EVAL_2694 = {1'h0,_EVAL_3374,_EVAL_240};
  assign _EVAL_5004 = {{6'd0}, _EVAL_5501};
  assign _EVAL_2319 = _EVAL_3591 ? _EVAL_5828 : _EVAL_3605;
  assign _EVAL_1787 = {_EVAL_340,_EVAL_1288};
  assign _EVAL_5168 = _EVAL_1763 <= 4'h8;
  assign _EVAL_5485 = _EVAL_1430 ? 1'h0 : 1'h1;
  assign _EVAL_3703 = _EVAL_343 ? {{1'd0}, _EVAL_2867} : _EVAL_4998;
  assign _EVAL_4355 = _EVAL_5951 & _EVAL_3200;
  assign _EVAL_145 = _EVAL_3404;
  assign _EVAL_2777 = {1'h0,_EVAL_3965,_EVAL_1026};
  assign _EVAL_2532 = {{1'd0}, _EVAL_2813};
  assign _EVAL_706 = {1'h0,_EVAL_5484};
  assign _EVAL_5019 = _EVAL_4553 ? _EVAL_673 : _EVAL_3086;
  assign _EVAL_4822 = _EVAL_2912 & _EVAL_417;
  assign _EVAL_3127 = {{6'd0}, _EVAL_4505};
  assign _EVAL_4924 = 2'h2 | _EVAL_1918;
  assign _EVAL_3885 = {1'h0,_EVAL_1229,_EVAL_4217};
  assign _EVAL_2535 = _EVAL_2473 ? _EVAL_1943 : _EVAL_5460;
  assign _EVAL_642 = _EVAL_308 ? _EVAL_2003 : _EVAL_1469;
  assign _EVAL_730 = {_EVAL_5024,_EVAL_2629};
  assign _EVAL_5405 = _EVAL_5068[582];
  assign _EVAL_5804 = _EVAL_4583 ? 8'hff : 8'h0;
  assign _EVAL_3912 = _EVAL_3047 == 4'hf;
  assign _EVAL_5745 = _EVAL_1477 & _EVAL_847;
  assign _EVAL_5762 = 10'h260 == _EVAL_5757;
  assign _EVAL_598 = {1'h0,_EVAL_3584,_EVAL_5065};
  assign _EVAL_841 = _EVAL_930 ? 1'h0 : 1'h1;
  assign _EVAL_557 = _EVAL_1608 & _EVAL_4477;
  assign _EVAL_2352 = _EVAL_3275 > _EVAL_5824;
  assign _EVAL_3353 = {_EVAL_3876,_EVAL_1720};
  assign _EVAL_5820 = {1'h0,_EVAL_5535,_EVAL_366};
  assign _EVAL_545 = _EVAL_1775[47:40];
  assign _EVAL_732 = _EVAL_2092 ? _EVAL_1400 : _EVAL_494;
  assign _EVAL_78 = _EVAL_1581;
  assign _EVAL_4943 = {{1'd0}, _EVAL_3411};
  assign _EVAL_669 = _EVAL_5125 & _EVAL_1937;
  assign _EVAL_3922 = _EVAL_6021 & _EVAL_906;
  assign _EVAL_2752 = {_EVAL_3516,_EVAL_3449};
  assign _EVAL_2499 = _EVAL_5174 & _EVAL_4247;
  assign _EVAL_3012 = {1'h0,_EVAL_355};
  assign _EVAL_2098 = _EVAL_4402 ? _EVAL_673 : _EVAL_5253;
  assign _EVAL_5944 = _EVAL_3941 ? _EVAL_5279 : _EVAL_665;
  assign _EVAL_2575 = _EVAL_5314 & _EVAL_3154;
  assign _EVAL_4127 = 10'h21a == _EVAL_5757;
  assign _EVAL_5928 = _EVAL_4478 & _EVAL_673;
  assign _EVAL_4328 = {1'h0,_EVAL_1765};
  assign _EVAL_3735 = _EVAL_1378 & _EVAL_1937;
  assign _EVAL_2010 = {{6'd0}, _EVAL_2694};
  assign _EVAL_2434 = {1'h0,_EVAL_2847,_EVAL_5701};
  assign _EVAL_1508 = 6'h20 | _EVAL_2114;
  assign _EVAL_5628 = _EVAL_1030 ? _EVAL_673 : _EVAL_3090;
  assign _EVAL_2882 = _EVAL_4637 ? _EVAL_371 : _EVAL_2391;
  assign _EVAL_4505 = {1'h0,_EVAL_2291};
  assign _EVAL_2391 = _EVAL_2190 ? _EVAL_4893 : _EVAL_3936;
  assign _EVAL_5126 = {1'h0,_EVAL_2484};
  assign _EVAL_5495 = {_EVAL_4344,_EVAL_1484};
  assign _EVAL_3559 = {_EVAL_5389,4'hf,_EVAL_4404,4'hf,_EVAL_1273,4'hf,_EVAL_272,4'hf};
  assign _EVAL_2707 = 10'h283 == _EVAL_5757;
  assign _EVAL_3469 = {_EVAL_6074,_EVAL_3857};
  assign _EVAL_4556 = _EVAL_5835 & _EVAL_673;
  assign _EVAL_1257 = _EVAL_5089 ? _EVAL_673 : _EVAL_3016;
  assign _EVAL_4746 = _EVAL_3465 > _EVAL_5183;
  assign _EVAL_4142 = _EVAL_2146 > _EVAL_5322;
  assign _EVAL_1572 = {_EVAL_4884,_EVAL_3289,_EVAL_3452,_EVAL_2865};
  assign _EVAL_5903 = _EVAL_301 | _EVAL_5221;
  assign _EVAL_1333 = _EVAL_325 == 22'h2cc0;
  assign _EVAL_3268 = _EVAL_393 ? _EVAL_3277 : _EVAL_3960;
  assign _EVAL_4285 = {{6'd0}, _EVAL_3729};
  assign _EVAL_1238 = _EVAL_5557 ? _EVAL_6067 : _EVAL_2865;
  assign _EVAL_2912 = _EVAL_1431 & _EVAL_673;
  assign _EVAL_2709 = {{1'd0}, _EVAL_4128};
  assign _EVAL_765 = _EVAL_2380 & _EVAL_847;
  assign _EVAL_4895 = 10'h215 == _EVAL_5757;
  assign _EVAL_1844 = _EVAL_5511 & _EVAL_847;
  assign _EVAL_5963 = {{6'd0}, _EVAL_677};
  assign _EVAL_1683 = _EVAL_4523 ? _EVAL_673 : _EVAL_3865;
  assign _EVAL_1251 = _EVAL_3843 & _EVAL_1831;
  assign _EVAL_5567 = _EVAL_4244 ? {{1'd0}, _EVAL_2642} : _EVAL_604;
  assign _EVAL_3099 = 10'h29b == _EVAL_5757;
  assign _EVAL_5862 = _EVAL_5002 & _EVAL_1041;
  assign _EVAL_4771 = {{6'd0}, _EVAL_4758};
  assign _EVAL_4980 = _EVAL_5951 & _EVAL_5267;
  assign _EVAL_4046 = {1'h0,_EVAL_1235};
  assign _EVAL_2249 = _EVAL_5846 & _EVAL_1407;
  assign _EVAL_2070 = _EVAL_1229 & _EVAL_1602;
  assign _EVAL_5504 = {_EVAL_4901,_EVAL_3692};
  assign _EVAL_4298 = {_EVAL_4574,4'hf,_EVAL_1288,4'hf,_EVAL_3692,4'hf,_EVAL_1672,4'hf};
  assign _EVAL_2160 = _EVAL_212 & _EVAL_3280;
  assign _EVAL_2853 = {{6'd0}, _EVAL_2330};
  assign _EVAL_1976 = _EVAL_1564[7:0];
  assign _EVAL_1119 = _EVAL_4621 ? _EVAL_2883 : _EVAL_405;
  assign _EVAL_2949 = {_EVAL_5537,4'hf,_EVAL_2030,4'hf,_EVAL_5962,4'hf,_EVAL_5606,4'hf};
  assign _EVAL_2267 = {1'h0,_EVAL_1057};
  assign _EVAL_2958 = _EVAL_5728 > _EVAL_2159;
  assign _EVAL_3795 = _EVAL_2058 & _EVAL_417;
  assign _EVAL_3656 = {_EVAL_3443,_EVAL_2546};
  assign _EVAL_1258 = {1'h0,_EVAL_4443,_EVAL_1527};
  assign _EVAL_738 = {1'h0,_EVAL_1826,_EVAL_2439};
  assign _EVAL_5885 = _EVAL_4226 ? _EVAL_673 : _EVAL_5942;
  assign _EVAL_3517 = _EVAL_3814 & _EVAL_1937;
  assign _EVAL_1595 = _EVAL_3783 & _EVAL_1383;
  assign _EVAL_5472 = _EVAL_5951 & _EVAL_2281;
  assign intsink__EVAL_2 = _EVAL_60;
  assign _EVAL_1949 = _EVAL_6049 & _EVAL_847;
  assign _EVAL_1662 = 3'h4 | _EVAL_3696;
  assign _EVAL_4247 = _EVAL_350 == 8'hff;
  assign Queue__EVAL_16 = _EVAL_4986[21:0];
  assign _EVAL_161 = {1'h0,_EVAL_1396,_EVAL_3020};
  assign _EVAL_4509 = {1'h0,_EVAL_1211,_EVAL_1868};
  assign _EVAL_2598 = _EVAL_762 & _EVAL_2756;
  assign _EVAL_838 = {{6'd0}, _EVAL_1556};
  assign _EVAL_5909 = _EVAL_3212 & _EVAL_2756;
  assign _EVAL_1253 = _EVAL_942 ? {{1'd0}, _EVAL_1168} : _EVAL_3862;
  assign _EVAL_5951 = _EVAL_970 & _EVAL_4602;
  assign _EVAL_3140 = _EVAL_5951 & _EVAL_5556;
  assign _EVAL_5957 = _EVAL_5511 & _EVAL_3487;
  assign _EVAL_2512 = _EVAL_6035 ? _EVAL_518 : _EVAL_4716;
  assign _EVAL_4875 = {1'h0,_EVAL_5300,_EVAL_5694};
  assign _EVAL_5010 = _EVAL_1843 & _EVAL_673;
  assign _EVAL_4477 = _EVAL_1159[16];
  assign _EVAL_2534 = {1'h0,1'h0,_EVAL_5265};
  assign _EVAL_948 = _EVAL_5052 & _EVAL_3487;
  assign _EVAL_1218 = _EVAL_3864 ? 1'h0 : 1'h1;
  assign _EVAL_160 = 10'h243 == _EVAL_5757;
  assign _EVAL_1614 = 10'h209 == _EVAL_5757;
  assign _EVAL_3808 = 4'h8 | _EVAL_3534;
  assign _EVAL_4282 = _EVAL_1751 & _EVAL_1937;
  assign _EVAL_2137 = {1'h0,_EVAL_3194,_EVAL_2549};
  assign _EVAL_2674 = _EVAL_1790 & _EVAL_847;
  assign _EVAL_1522 = {{6'd0}, _EVAL_286};
  assign _EVAL_2350 = _EVAL_5905 == 4'hf;
  assign _EVAL_2867 = _EVAL_4809 ? 1'h0 : 1'h1;
  assign _EVAL_1990 = _EVAL_381 & _EVAL_4922;
  assign _EVAL_5712 = {1'h0,_EVAL_5255,_EVAL_526};
  assign _EVAL_4905 = {{6'd0}, _EVAL_5301};
  assign _EVAL_1093 = _EVAL_5068[604];
  assign _EVAL_2861 = _EVAL_1608 & _EVAL_3154;
  assign _EVAL_4076 = {1'h0,_EVAL_2215};
  assign _EVAL_2114 = {{1'd0}, _EVAL_5567};
  assign _EVAL_4249 = {{1'd0}, _EVAL_5198};
  assign _EVAL_1589 = _EVAL_5151 & _EVAL_1937;
  assign _EVAL_4741 = _EVAL_2218[23:16];
  assign _EVAL_5682 = _EVAL_4291 & _EVAL_1287;
  assign _EVAL_1106 = _EVAL_2218[31:24];
  assign _EVAL_394 = {{6'd0}, _EVAL_2267};
  assign _EVAL_3827 = _EVAL_559 ? _EVAL_673 : _EVAL_3637;
  assign _EVAL_397 = _EVAL_5096 & _EVAL_847;
  assign _EVAL_559 = 10'h211 == _EVAL_5757;
  assign _EVAL_2938 = _EVAL_3597 ? _EVAL_673 : _EVAL_4303;
  assign _EVAL_2186 = {{6'd0}, _EVAL_6020};
  assign _EVAL_2111 = Queue__EVAL_8[5];
  assign _EVAL_3154 = _EVAL_1159[8];
  assign _EVAL_2237 = _EVAL_3423[63:0];
  assign _EVAL_5701 = {{6'd0}, _EVAL_639};
  assign _EVAL_5413 = _EVAL_2936 ? _EVAL_1119 : _EVAL_5925;
  assign _EVAL_5429 = _EVAL_5951 & _EVAL_3757;
  assign _EVAL_5562 = {{1'd0}, _EVAL_3895};
  assign _EVAL_609 = {{6'd0}, _EVAL_2336};
  assign _EVAL_3890 = _EVAL_1598 ? _EVAL_673 : _EVAL_5109;
  assign _EVAL_4268 = _EVAL_5951 & _EVAL_2394;
  assign _EVAL_1250 = _EVAL_5836 & _EVAL_1937;
  assign _EVAL_5513 = {{1'd0}, _EVAL_1531};
  assign _EVAL_2716 = {{6'd0}, _EVAL_750};
  assign _EVAL_2120 = _EVAL_4978 ? {{1'd0}, _EVAL_5677} : _EVAL_170;
  assign _EVAL_5611 = _EVAL_2596 ? _EVAL_673 : _EVAL_3621;
  assign _EVAL_2054 = {_EVAL_4301,_EVAL_5665};
  assign _EVAL_4412 = _EVAL_2751 > _EVAL_1023;
  assign _EVAL_1219 = _EVAL_5093 ? _EVAL_673 : _EVAL_5459;
  assign _EVAL_1174 = 3'h4 | _EVAL_2856;
  assign _EVAL_4116 = 10'h286 == _EVAL_5757;
  assign _EVAL_1335 = _EVAL_1598 ? _EVAL_2812 : _EVAL_5805;
  assign _EVAL_267 = _EVAL_5951 & _EVAL_4162;
  assign _EVAL_416 = _EVAL_2197 ? _EVAL_1422 : _EVAL_5384;
  assign _EVAL_1918 = {{1'd0}, _EVAL_1979};
  assign _EVAL_3985 = _EVAL_5068[658];
  assign _EVAL_1005 = _EVAL_4734 & _EVAL_417;
  assign _EVAL_494 = _EVAL_2369 ? _EVAL_1550 : _EVAL_959;
  assign _EVAL_3916 = _EVAL_3987 ? 1'h0 : 1'h1;
  assign _EVAL_2932 = {{6'd0}, _EVAL_4823};
  assign _EVAL_2804 = _EVAL_5010 & _EVAL_2350;
  assign _EVAL_3411 = _EVAL_2112 ? {{1'd0}, _EVAL_548} : _EVAL_969;
  assign _EVAL_3018 = {1'h0,_EVAL_1641};
  assign _EVAL_2077 = _EVAL_5068[645];
  assign _EVAL_6072 = {{6'd0}, _EVAL_4875};
  assign _EVAL_1785 = {_EVAL_3922,_EVAL_5080};
  assign _EVAL_5595 = _EVAL_1309 ? _EVAL_673 : _EVAL_5019;
  assign _EVAL_760 = _EVAL_4053 & _EVAL_1645;
  assign _EVAL_4345 = _EVAL_430 > _EVAL_4165;
  assign _EVAL_3111 = 2'h2 | _EVAL_5645;
  assign _EVAL_4484 = {{1'd0}, _EVAL_2136};
  assign _EVAL_3031 = _EVAL_4749 ? _EVAL_673 : _EVAL_4067;
  assign _EVAL_3970 = _EVAL_520 ? _EVAL_2186 : _EVAL_4921;
  assign _EVAL_5655 = {{6'd0}, _EVAL_2843};
  assign _EVAL_5863 = _EVAL_2351 ? _EVAL_5523 : _EVAL_414;
  assign _EVAL_5742 = {_EVAL_5624,4'hf,_EVAL_4927,4'hf,_EVAL_5139,4'hf,_EVAL_607,4'hf};
  assign _EVAL_4610 = _EVAL_2595 & _EVAL_417;
  assign _EVAL_3621 = _EVAL_3941 ? _EVAL_673 : _EVAL_1476;
  assign _EVAL_5783 = {1'h0,_EVAL_2229,_EVAL_2389};
  assign _EVAL_2257 = {{6'd0}, _EVAL_3272};
  assign _EVAL_220 = _EVAL_2603 ? _EVAL_5044 : _EVAL_3219;
  assign _EVAL_939 = 10'h29f == _EVAL_5757;
  assign _EVAL_3899 = _EVAL_5174 & _EVAL_5871;
  assign _EVAL_4626 = 10'h220 == _EVAL_5757;
  assign _EVAL_2052 = _EVAL_5068[599];
  assign _EVAL_5913 = _EVAL_1159[15:12];
  assign _EVAL_3786 = _EVAL_4636 > _EVAL_5441;
  assign _EVAL_3758 = _EVAL_1347 & _EVAL_847;
  assign _EVAL_2666 = _EVAL_2308 & _EVAL_3580;
  assign _EVAL_3530 = _EVAL_246 & _EVAL_1937;
  assign _EVAL_4068 = _EVAL_644 & _EVAL_5484;
  assign _EVAL_3791 = _EVAL_1309 ? _EVAL_3229 : _EVAL_3800;
  assign _EVAL_4256 = {1'h0,_EVAL_1493};
  assign _EVAL_3757 = _EVAL_5068[0];
  assign _EVAL_1806 = _EVAL_5073 & _EVAL_673;
  assign _EVAL_3979 = 10'h248 == _EVAL_5757;
  assign _EVAL_2522 = _EVAL_1228 ? _EVAL_4064 : _EVAL_1904;
  assign _EVAL_813 = _EVAL_3456 & _EVAL_5409;
  assign _EVAL_483 = {_EVAL_4815,_EVAL_2626};
  assign _EVAL_3613 = _EVAL_5068[610];
  assign _EVAL_1848 = _EVAL_4772 ? _EVAL_673 : _EVAL_1766;
  assign _EVAL_3045 = {_EVAL_1863,4'hf,_EVAL_3040,4'hf,_EVAL_2307,4'hf,_EVAL_3256,4'hf};
  assign _EVAL_5093 = 10'h250 == _EVAL_5757;
  assign _EVAL_3563 = _EVAL_4127 ? _EVAL_673 : _EVAL_3426;
  assign _EVAL_1403 = _EVAL_6064 & _EVAL_673;
  assign _EVAL_1474 = {_EVAL_6071,_EVAL_4700};
  assign Queue__EVAL_1 = _EVAL_77;
  assign _EVAL_2621 = _EVAL_4340 & _EVAL_673;
  assign _EVAL_3793 = _EVAL_3717 ? {{1'd0}, _EVAL_1098} : _EVAL_1912;
  assign _EVAL_1072 = _EVAL_5068[674];
  assign _EVAL_2491 = {{6'd0}, _EVAL_4897};
  assign _EVAL_953 = {_EVAL_1515,4'hf,_EVAL_4390,4'hf,_EVAL_4624,4'hf,_EVAL_5009,4'hf};
  assign _EVAL_4386 = _EVAL_5068[592];
  assign _EVAL_5150 = _EVAL_6073 & _EVAL_4477;
  assign _EVAL_4234 = _EVAL_4820 ? {{1'd0}, _EVAL_5715} : _EVAL_2887;
  assign _EVAL_2337 = {{6'd0}, _EVAL_5394};
  assign _EVAL_4725 = {_EVAL_2964,_EVAL_411,_EVAL_4438,_EVAL_3299,_EVAL_4489,_EVAL_4528,_EVAL_5107,_EVAL_514};
  assign _EVAL_1444 = _EVAL_2215 & _EVAL_3294;
  assign _EVAL_3426 = _EVAL_1935 ? _EVAL_673 : _EVAL_5885;
  assign _EVAL_662 = {{6'd0}, _EVAL_4107};
  assign _EVAL_4603 = {_EVAL_4467,_EVAL_4927};
  assign _EVAL_986 = {_EVAL_2781,4'hf,_EVAL_2626,4'hf,_EVAL_3857,4'hf,_EVAL_1186,4'hf};
  assign _EVAL_2970 = {{6'd0}, _EVAL_4046};
  assign _EVAL_324 = {{6'd0}, _EVAL_3724};
  assign _EVAL_5972 = {_EVAL_2070,_EVAL_4518};
  assign _EVAL_2226 = {1'h0,_EVAL_5411,_EVAL_4161};
  assign _EVAL_5881 = _EVAL_3404 & _EVAL_5635;
  assign _EVAL_2952 = _EVAL_5068[600];
  assign _EVAL_3494 = {1'h0,_EVAL_2381,_EVAL_1267};
  assign _EVAL_5923 = {_EVAL_5390,_EVAL_5981};
  assign _EVAL_5614 = _EVAL_4272 ? {{1'd0}, _EVAL_3446} : _EVAL_3745;
  assign _EVAL_5098 = {_EVAL_1200,_EVAL_4019};
  assign _EVAL_4968 = _EVAL_1057 & _EVAL_5307;
  assign _EVAL_784 = _EVAL_2961 ? _EVAL_4771 : _EVAL_2512;
  assign _EVAL_4244 = _EVAL_4274 > _EVAL_5555;
  assign _EVAL_317 = _EVAL_2341 & _EVAL_2203;
  assign _EVAL_3564 = _EVAL_5068[648];
  assign _EVAL_4410 = 10'h297 == _EVAL_5757;
  assign _EVAL_5494 = _EVAL_2719 ? 1'h0 : 1'h1;
  assign _EVAL_5847 = {1'h0,_EVAL_3940,_EVAL_4179};
  assign _EVAL_6046 = _EVAL_5468 & _EVAL_2756;
  assign _EVAL_3368 = {_EVAL_2160,_EVAL_5008};
  assign _EVAL_5591 = _EVAL_5836 & _EVAL_417;
  assign _EVAL_4339 = _EVAL_2058 & _EVAL_2350;
  assign _EVAL_1877 = _EVAL_1860 & _EVAL_847;
  assign _EVAL_405 = {_EVAL_1251,_EVAL_1797};
  assign _EVAL_3724 = {1'h0,_EVAL_3986};
  assign _EVAL_5224 = {{6'd0}, _EVAL_1445};
  assign _EVAL_879 = _EVAL_5174 & _EVAL_3043;
  assign _EVAL_716 = {{6'd0}, _EVAL_962};
  assign _EVAL_3110 = _EVAL_5337 ? _EVAL_673 : _EVAL_4466;
  assign _EVAL_497 = {{6'd0}, _EVAL_3019};
  assign _EVAL_306 = _EVAL_2784 & _EVAL_2756;
  assign _EVAL_5835 = _EVAL_5951 & _EVAL_2520;
  assign _EVAL_5115 = _EVAL_5068[609];
  assign _EVAL_742 = _EVAL_5951 & _EVAL_3613;
  assign _EVAL_3325 = _EVAL_2967 > _EVAL_1799;
  assign _EVAL_6074 = _EVAL_5940 & _EVAL_4398;
  assign _EVAL_648 = {1'h0,_EVAL_6030};
  assign _EVAL_2823 = _EVAL_3662 ? _EVAL_673 : _EVAL_2938;
  assign _EVAL_1275 = {{1'd0}, _EVAL_400};
  assign _EVAL_2654 = {{30'd0}, _EVAL_4496};
  assign _EVAL_959 = _EVAL_835 ? _EVAL_3271 : _EVAL_1368;
  assign _EVAL_3277 = {_EVAL_5518,4'hf,_EVAL_2920,4'hf,_EVAL_3676,4'hf,_EVAL_5713,4'hf};
  assign _EVAL_547 = _EVAL_3499 & _EVAL_847;
  assign _EVAL_5585 = _EVAL_1737 ? 1'h0 : 1'h1;
  assign _EVAL_889 = _EVAL_796 & _EVAL_3487;
  assign _EVAL_3751 = {1'h0,_EVAL_2993,_EVAL_2488};
  assign _EVAL_3542 = _EVAL_5222 & _EVAL_2350;
  assign _EVAL_1907 = _EVAL_1875 & _EVAL_5558;
  assign _EVAL_3997 = _EVAL_4356 ? _EVAL_198 : _EVAL_1474;
  assign _EVAL_5571 = _EVAL_320 ? 1'h0 : 1'h1;
  assign _EVAL_180 = {1'h0,_EVAL_1131,_EVAL_1519};
  assign _EVAL_3042 = 2'h2 | _EVAL_2053;
  assign _EVAL_4583 = Queue__EVAL_4[3];
  assign _EVAL_3391 = _EVAL_2683 & _EVAL_1292;
  assign _EVAL_4511 = _EVAL_6061 ? _EVAL_4058 : _EVAL_2819;
  assign _EVAL_2671 = {1'h0,_EVAL_2667};
  assign _EVAL_5222 = _EVAL_5801 & _EVAL_673;
  assign _EVAL_3927 = _EVAL_5951 & _EVAL_2706;
  assign _EVAL_1159 = {_EVAL_5804,_EVAL_1080,_EVAL_1959,_EVAL_5969};
  assign _EVAL_3048 = _EVAL_1159[31:24];
  assign _EVAL_67 = _EVAL_5933 ? _EVAL_3938 : 32'h0;
  assign _EVAL_4056 = {{6'd0}, _EVAL_2156};
  assign _EVAL_1968 = _EVAL_3987 ? _EVAL_5732 : 5'h0;
  assign _EVAL_1117 = _EVAL_2782 & _EVAL_666;
  assign _EVAL_501 = _EVAL_285 > _EVAL_3023;
  assign _EVAL_696 = _EVAL_1403 & _EVAL_2756;
  assign _EVAL_3729 = {1'h0,_EVAL_5684,_EVAL_2408};
  assign _EVAL_1042 = _EVAL_1654 ? 1'h0 : 1'h1;
  assign _EVAL_3716 = _EVAL_3318 & _EVAL_4477;
  assign _EVAL_344 = {{4'd0}, _EVAL_3385};
  assign _EVAL_393 = 10'h2a1 == _EVAL_5757;
  assign _EVAL_2158 = {{6'd0}, _EVAL_1330};
  assign _EVAL_1252 = _EVAL_4458 > _EVAL_1571;
  assign _EVAL_1699 = _EVAL_5068[675];
  assign _EVAL_4611 = 3'h4 | _EVAL_4719;
  assign _EVAL_379 = {{6'd0}, _EVAL_2448};
  assign _EVAL_1248 = 10'h212 == _EVAL_5757;
  assign _EVAL_2898 = _EVAL_5068[671];
  assign _EVAL_3304 = _EVAL_5883 ? _EVAL_673 : _EVAL_1257;
  assign _EVAL_601 = _EVAL_4556 & _EVAL_2756;
  assign _EVAL_1565 = _EVAL_4010 & _EVAL_3154;
  assign _EVAL_4452 = 10'h284 == _EVAL_5757;
  assign _EVAL_6019 = {1'h0,_EVAL_896,_EVAL_188};
  assign _EVAL_5137 = {1'h0,_EVAL_1880,_EVAL_5915};
  assign _EVAL_4204 = 10'h24a == _EVAL_5757;
  assign _EVAL_3796 = _EVAL_812 ? _EVAL_1504 : _EVAL_5996;
  assign _EVAL_1549 = {{6'd0}, _EVAL_4509};
  assign _EVAL_1903 = _EVAL_1472 > _EVAL_3997;
  assign _EVAL_2359 = _EVAL_3925 ? _EVAL_4740 : _EVAL_4776;
  assign _EVAL_3745 = 2'h2 | _EVAL_5393;
  assign _EVAL_5815 = _EVAL_3431 > _EVAL_685;
  assign _EVAL_2311 = _EVAL_5521 & _EVAL_2918;
  assign _EVAL_1466 = {{6'd0}, _EVAL_4292};
  assign _EVAL_3876 = _EVAL_4965 & _EVAL_1820;
  assign _EVAL_1092 = _EVAL_5768[15:1];
  assign _EVAL_3597 = 10'h214 == _EVAL_5757;
  assign _EVAL_4526 = _EVAL_4948 ? {{1'd0}, _EVAL_1429} : _EVAL_1817;
  assign _EVAL_5803 = {_EVAL_4942,_EVAL_4404};
  assign _EVAL_2189 = _EVAL_5951 & _EVAL_3805;
  assign _EVAL_4376 = _EVAL_4124 ? _EVAL_4699 : _EVAL_2315;
  assign _EVAL_3123 = {{6'd0}, _EVAL_2845};
  assign _EVAL_5710 = {1'h0,_EVAL_3607,_EVAL_3334};
  assign _EVAL_2408 = {{6'd0}, _EVAL_2901};
  assign _EVAL_1074 = {_EVAL_1066,_EVAL_1629};
  assign _EVAL_5555 = _EVAL_1252 ? _EVAL_4458 : _EVAL_1571;
  assign _EVAL_705 = _EVAL_2428 ? _EVAL_4298 : _EVAL_1857;
  assign _EVAL_2018 = _EVAL_4621 ? 1'h0 : 1'h1;
  assign _EVAL_308 = _EVAL_2003 > _EVAL_1469;
  assign _EVAL_1222 = 2'h2 | _EVAL_2532;
  assign _EVAL_2563 = {1'h0,_EVAL_2782,_EVAL_1969};
  assign _EVAL_2013 = _EVAL_3847 & _EVAL_5878;
  assign _EVAL_3003 = {{6'd0}, _EVAL_3604};
  assign _EVAL_4358 = _EVAL_2050 ? _EVAL_4267 : _EVAL_5324;
  assign _EVAL_2377 = _EVAL_5068[598];
  assign _EVAL_371 = {_EVAL_780,4'hf,_EVAL_4518,4'hf,_EVAL_493,4'hf,_EVAL_1052,4'hf};
  assign _EVAL_4105 = {{6'd0}, _EVAL_2410};
  assign _EVAL_2519 = _EVAL_516 & _EVAL_3487;
  assign _EVAL_4246 = _EVAL_5068[663];
  assign _EVAL_6004 = _EVAL_5068[255];
  assign _EVAL_4036 = {1'h0,_EVAL_2247,_EVAL_5891};
  assign _EVAL_350 = _EVAL_1159[23:16];
  assign _EVAL_3839 = _EVAL_2180 ? 1'h0 : 1'h1;
  assign _EVAL_5730 = _EVAL_6053 & _EVAL_1937;
  assign _EVAL_1748 = _EVAL_1758 ? 1'h0 : 1'h1;
  assign _EVAL_2866 = {1'h0,_EVAL_1188,_EVAL_3141};
  assign _EVAL_516 = _EVAL_5769 & _EVAL_673;
  assign intsink__EVAL = _EVAL_106;
  assign _EVAL_5314 = _EVAL_3763 & _EVAL_673;
  assign _EVAL_2156 = {1'h0,_EVAL_4588,_EVAL_3913};
  assign _EVAL_5143 = _EVAL_2968 ? _EVAL_673 : _EVAL_3351;
  assign _EVAL_3482 = {{6'd0}, _EVAL_2137};
  assign _EVAL_1809 = _EVAL_1806 & _EVAL_847;
  assign _EVAL_312 = {1'h0,_EVAL_2690,_EVAL_165};
  assign _EVAL_5603 = _EVAL_5821 & _EVAL_847;
  assign _EVAL_4899 = {1'h0,_EVAL_2357,_EVAL_5709};
  assign _EVAL_5785 = {{6'd0}, _EVAL_4090};
  assign _EVAL_1221 = {_EVAL_913,_EVAL_2307};
  assign _EVAL_1303 = {{1'd0}, _EVAL_1554};
  assign _EVAL_1429 = _EVAL_3618 ? {{1'd0}, _EVAL_855} : _EVAL_2138;
  assign _EVAL_5048 = 10'h201 == _EVAL_5757;
  assign _EVAL_4791 = Queue__EVAL_2;
  assign _EVAL_3560 = {1'h0,_EVAL_4080,_EVAL_4143};
  assign _EVAL_297 = _EVAL_3796 > _EVAL_700;
  assign _EVAL_3879 = _EVAL_5951 & _EVAL_5516;
  assign _EVAL_901 = _EVAL_5330 ? _EVAL_1609 : _EVAL_664;
  assign _EVAL_4271 = _EVAL_2516 & _EVAL_2580;
  assign _EVAL_3299 = _EVAL_3390 ? _EVAL_6067 : _EVAL_851;
  assign _EVAL_1456 = {{4'd0}, _EVAL_902};
  assign _EVAL_2372 = _EVAL_5951 & _EVAL_1706;
  assign _EVAL_5836 = _EVAL_881 & _EVAL_673;
  assign _EVAL_2874 = {{6'd0}, _EVAL_738};
  assign _EVAL_1621 = _EVAL_1337 > _EVAL_3654;
  assign _EVAL_1315 = _EVAL_2046 ? _EVAL_3732 : _EVAL_1849;
  assign _EVAL_4972 = {1'h0,_EVAL_1917,_EVAL_4848};
  assign _EVAL_685 = _EVAL_3325 ? _EVAL_2967 : _EVAL_1799;
  assign _EVAL_3357 = {1'h0,_EVAL_4620,_EVAL_1466};
  assign _EVAL_2061 = {{6'd0}, _EVAL_918};
  assign _EVAL_5172 = _EVAL_1477 & _EVAL_4477;
  assign _EVAL_1372 = {_EVAL_1106,_EVAL_4741,_EVAL_681,_EVAL_1011};
  assign _EVAL_4272 = _EVAL_4540 > _EVAL_1359;
  assign _EVAL_5323 = _EVAL_5435 ? 2'h0 : 2'h3;
  assign _EVAL_1815 = _EVAL_4266 > _EVAL_863;
  assign _EVAL_5146 = {{6'd0}, _EVAL_5346};
  assign _EVAL_5821 = _EVAL_4355 & _EVAL_673;
  assign _EVAL_4749 = 10'h29d == _EVAL_5757;
  assign _EVAL_5256 = 10'h294 == _EVAL_5757;
  assign _EVAL_5120 = _EVAL_5952 > _EVAL_5503;
  assign _EVAL_3043 = _EVAL_5000 == 8'hff;
  assign _EVAL_4058 = {_EVAL_2895,_EVAL_2806};
  assign _EVAL_1021 = _EVAL_1900 ? {{1'd0}, _EVAL_4497} : _EVAL_1230;
  assign _EVAL_4236 = _EVAL_5432 & _EVAL_4477;
  assign _EVAL_3799 = _EVAL_2912 & _EVAL_1937;
  assign _EVAL_2728 = _EVAL_1569 & _EVAL_1333;
  assign _EVAL_2196 = {1'h0,_EVAL_5916,_EVAL_5176};
  assign _EVAL_2865 = _EVAL_2218[39:32];
  assign _EVAL_5551 = _EVAL_846 ? _EVAL_1441 : _EVAL_3035;
  assign _EVAL_3662 = 10'h213 == _EVAL_5757;
  assign _EVAL_2155 = _EVAL_4268 & _EVAL_673;
  assign _EVAL_2824 = {_EVAL_2851,_EVAL_6040};
  assign _EVAL_4156 = {1'h0,_EVAL_5846,_EVAL_4622};
  assign _EVAL_3907 = {1'h0,_EVAL_4308,_EVAL_2716};
  assign _EVAL_4009 = _EVAL_5256 ? _EVAL_673 : _EVAL_3105;
  assign _EVAL_2136 = _EVAL_3925 ? {{1'd0}, _EVAL_2590} : _EVAL_5884;
  assign _EVAL_2428 = 10'h298 == _EVAL_5757;
  assign _EVAL_1843 = _EVAL_5951 & _EVAL_3466;
  assign _EVAL_6066 = _EVAL_4672 ? _EVAL_729 : _EVAL_5661;
  assign _EVAL_4161 = {{6'd0}, _EVAL_1964};
  assign _EVAL_5491 = _EVAL_5068[660];
  assign _EVAL_2961 = 10'h24b == _EVAL_5757;
  assign _EVAL_463 = _EVAL_5468 & _EVAL_417;
  assign _EVAL_2342 = _EVAL_4387 > _EVAL_3893;
  assign _EVAL_3870 = _EVAL_1184 - 4'h1;
  assign _EVAL_3731 = _EVAL_4646 > _EVAL_2761;
  assign _EVAL_4685 = 8'h80 | _EVAL_1456;
  assign _EVAL_1362 = {1'h0,_EVAL_727,_EVAL_4590};
  assign _EVAL_2719 = _EVAL_2188 > _EVAL_2332;
  assign _EVAL_5931 = Queue__EVAL_8[0];
  assign _EVAL_2279 = {{6'd0}, _EVAL_2309};
  assign _EVAL_3212 = _EVAL_907 & _EVAL_673;
  assign _EVAL_5339 = _EVAL_4456 & _EVAL_673;
  assign _EVAL_4050 = _EVAL_4769 ? {{1'd0}, _EVAL_230} : _EVAL_5047;
  assign _EVAL_5278 = _EVAL_5939 ? _EVAL_673 : _EVAL_5462;
  assign _EVAL_3479 = _EVAL_5293 & _EVAL_4348;
  assign _EVAL_970 = Queue__EVAL_14 & _EVAL_34;
  assign _EVAL_5967 = _EVAL_270 ? 1'h0 : 1'h1;
  assign _EVAL_1979 = _EVAL_5791 ? 1'h0 : 1'h1;
  assign _EVAL_2380 = _EVAL_5577 & _EVAL_673;
  assign _EVAL_5390 = _EVAL_3181 & _EVAL_887;
  assign _EVAL_5996 = {_EVAL_1178,_EVAL_493};
  assign _EVAL_5876 = _EVAL_5989[15:2];
  assign _EVAL_2322 = _EVAL_5951 & _EVAL_1089;
  assign _EVAL_3274 = 2'h2 | _EVAL_4122;
  assign _EVAL_3332 = _EVAL_5397 ? _EVAL_806 : _EVAL_2896;
  assign _EVAL_520 = 10'h208 == _EVAL_5757;
  assign _EVAL_1368 = _EVAL_1140 ? _EVAL_5358 : _EVAL_3741;
  assign _EVAL_3020 = {{6'd0}, _EVAL_1961};
  assign _EVAL_2161 = 10'h205 == _EVAL_5757;
  assign _EVAL_1124 = {{1'd0}, _EVAL_2287};
  assign _EVAL_2843 = {1'h0,_EVAL_4233};
  assign _EVAL_1726 = _EVAL_5548 & _EVAL_673;
  assign _EVAL_3408 = _EVAL_2848 > _EVAL_672;
  assign _EVAL_5388 = {1'h0,_EVAL_2837};
  assign _EVAL_5813 = _EVAL_2065 & _EVAL_2766;
  assign _EVAL_1066 = _EVAL_2876 & _EVAL_4738;
  assign _EVAL_2090 = _EVAL_3891 ? {{1'd0}, _EVAL_4683} : _EVAL_3274;
  assign _EVAL_4704 = _EVAL_939 ? _EVAL_673 : _EVAL_2541;
  assign _EVAL_4292 = {1'h0,_EVAL_212,_EVAL_1859};
  assign _EVAL_1200 = _EVAL_1206 & _EVAL_1245;
  assign _EVAL_5374 = _EVAL_4159 ? _EVAL_673 : _EVAL_3827;
  assign _EVAL_1486 = 10'h256 == _EVAL_5757;
  assign _EVAL_1154 = _EVAL_163 ? _EVAL_673 : _EVAL_595;
  assign _EVAL_5768 = 16'h1 << _EVAL_5112;
  assign _EVAL_3823 = {_EVAL_1990,_EVAL_5139};
  assign _EVAL_197 = _EVAL_5821 & _EVAL_3154;
  assign _EVAL_2805 = {_EVAL_1595,_EVAL_3693};
  assign _EVAL_3854 = _EVAL_1806 & _EVAL_3487;
  assign _EVAL_700 = _EVAL_3308 ? _EVAL_5972 : _EVAL_4770;
  assign _EVAL_190 = {{6'd0}, _EVAL_4156};
  assign _EVAL_811 = {1'h0,_EVAL_1777,_EVAL_5767};
  assign _EVAL_1912 = 2'h2 | _EVAL_3416;
  assign _EVAL_4986 = _EVAL_131[25:2];
  assign _EVAL_3893 = _EVAL_1381 ? _EVAL_329 : _EVAL_4530;
  assign _EVAL_2025 = _EVAL_2954 & _EVAL_4477;
  assign _EVAL_720 = _EVAL_3615 ? _EVAL_687 : _EVAL_4632;
  assign _EVAL_3427 = _EVAL_1159[7:4];
  assign _EVAL_4829 = _EVAL_2936 ? {{1'd0}, _EVAL_2018} : _EVAL_4924;
  assign _EVAL_2577 = _EVAL_1825 & _EVAL_1937;
  assign _EVAL_665 = _EVAL_4562 ? _EVAL_2435 : _EVAL_3507;
  assign _EVAL_5942 = _EVAL_5399 ? _EVAL_673 : _EVAL_1749;
  assign _EVAL_650 = _EVAL_5010 & _EVAL_2756;
  assign _EVAL_320 = _EVAL_674 > _EVAL_2080;
  assign _EVAL_2394 = _EVAL_5068[667];
  assign _EVAL_3131 = _EVAL_2180 ? _EVAL_5725 : _EVAL_5793;
  assign _EVAL_1560 = _EVAL_3752 ? _EVAL_4827 : _EVAL_3469;
  assign _EVAL_3603 = _EVAL_2366 & _EVAL_4051;
  assign _EVAL_1232 = {{6'd0}, _EVAL_2749};
  assign _EVAL_850 = _EVAL_5951 & _EVAL_2077;
  assign _EVAL_4377 = Queue__EVAL_8[3];
  assign _EVAL_2784 = _EVAL_4970 & _EVAL_673;
  assign _EVAL_1868 = {{6'd0}, _EVAL_1362};
  assign _EVAL_5807 = {_EVAL_5111,_EVAL_3005};
  assign _EVAL_1963 = {1'h0,_EVAL_2277,_EVAL_1497};
  assign _EVAL_1321 = 10'h249 == _EVAL_5757;
  assign _EVAL_1576 = _EVAL_427 ? _EVAL_5165 : _EVAL_2228;
  assign _EVAL_4978 = _EVAL_1577 > _EVAL_3790;
  assign _EVAL_2080 = {_EVAL_3056,_EVAL_1427};
  assign _EVAL_4679 = {{4'd0}, _EVAL_1587};
  assign _EVAL_1215 = _EVAL_1664 & _EVAL_3940;
  assign _EVAL_3496 = _EVAL_5951 & _EVAL_1072;
  assign _EVAL_2063 = _EVAL_2683 & _EVAL_3043;
  assign _EVAL_1352 = _EVAL_5068[577];
  assign _EVAL_4387 = _EVAL_5929 ? _EVAL_3585 : _EVAL_5058;
  assign _EVAL_3270 = _EVAL_3798 ? _EVAL_1520 : _EVAL_3126;
  assign _EVAL_3058 = _EVAL_1159[7:0];
  assign _EVAL_2854 = {1'h0,_EVAL_4584,_EVAL_3003};
  assign _EVAL_4493 = {{6'd0}, _EVAL_5186};
  assign _EVAL_846 = _EVAL_1441 > _EVAL_3035;
  assign _EVAL_3864 = _EVAL_3903 > _EVAL_3656;
  assign _EVAL_2239 = _EVAL_2701 & _EVAL_1937;
  assign _EVAL_4547 = _EVAL_5928 & _EVAL_1937;
  assign _EVAL_3535 = _EVAL_5068[655];
  assign _EVAL_5515 = _EVAL_320 ? _EVAL_674 : _EVAL_2080;
  assign _EVAL_1517 = {_EVAL_2343,_EVAL_607};
  assign _EVAL_4286 = {1'h0,_EVAL_582,_EVAL_1398};
  assign _EVAL_2787 = {_EVAL_2630,_EVAL_4479};
  assign _EVAL_5934 = {{6'd0}, _EVAL_4275};
  assign _EVAL_6079 = {{6'd0}, _EVAL_4041};
  assign _EVAL_1681 = Queue__EVAL_8[4];
  assign _EVAL_1141 = {{1'd0}, _EVAL_4517};
  assign _EVAL_2510 = _EVAL_4010 & _EVAL_3487;
  assign _EVAL_5844 = _EVAL_3665 ? _EVAL_2164 : _EVAL_1710;
  assign _EVAL_2199 = _EVAL_4863 ? _EVAL_1333 : _EVAL_1768;
  assign _EVAL_2603 = _EVAL_5044 > _EVAL_3219;
  assign _EVAL_606 = _EVAL_2757 & _EVAL_673;
  assign _EVAL_1925 = {1'h0,_EVAL_643};
  assign _EVAL_3317 = _EVAL_349 > _EVAL_3393;
  assign _EVAL_5958 = _EVAL_1153 ? _EVAL_1503 : _EVAL_3661;
  assign _EVAL_1534 = _EVAL_2958 ? _EVAL_5728 : _EVAL_2159;
  assign _EVAL_1564 = _EVAL_1674 | _EVAL_3836;
  assign _EVAL_5237 = {{6'd0}, _EVAL_2102};
  assign _EVAL_2212 = _EVAL_812 ? 1'h0 : 1'h1;
  assign _EVAL_5873 = _EVAL_5807 > _EVAL_5166;
  assign _EVAL_2034 = 10'h28c == _EVAL_5757;
  assign _EVAL_4663 = {{6'd0}, _EVAL_3742};
  assign _EVAL_4653 = _EVAL_5070 & _EVAL_673;
  assign _EVAL_4945 = _EVAL_5330 ? {{1'd0}, _EVAL_1021} : _EVAL_3808;
  assign _EVAL_1307 = _EVAL_3814 & _EVAL_2350;
  assign _EVAL_340 = _EVAL_2339 & _EVAL_4184;
  assign _EVAL_3606 = _EVAL_2161 ? _EVAL_3204 : _EVAL_5038;
  assign _EVAL_4994 = _EVAL_5951 & _EVAL_4386;
  assign _EVAL_1347 = _EVAL_3546 & _EVAL_673;
  assign _EVAL_1237 = _EVAL_2961 ? _EVAL_673 : _EVAL_353;
  assign _EVAL_255 = _EVAL_939 ? _EVAL_3559 : _EVAL_403;
  assign _EVAL_1654 = _EVAL_1997 > _EVAL_1221;
  assign _EVAL_294 = {_EVAL_1028,4'hf,_EVAL_4304,4'hf,_EVAL_3673,4'hf,_EVAL_563,4'hf};
  assign _EVAL_4176 = _EVAL_4272 ? _EVAL_4540 : _EVAL_1359;
  assign _EVAL_4173 = {1'h0,_EVAL_3629,_EVAL_182};
  assign _EVAL_5397 = 10'h259 == _EVAL_5757;
  assign _EVAL_5732 = {_EVAL_576,_EVAL_5311};
  assign _EVAL_3454 = {_EVAL_2457,_EVAL_2293};
  assign _EVAL_1495 = 6'h20 | _EVAL_6091;
  assign _EVAL_4143 = {{6'd0}, _EVAL_999};
  assign _EVAL_3204 = {{6'd0}, _EVAL_4580};
  assign _EVAL_4528 = _EVAL_4956 ? _EVAL_1035 : _EVAL_166;
  assign _EVAL_3549 = {{6'd0}, _EVAL_1791};
  assign _EVAL_4827 = {_EVAL_5225,_EVAL_1186};
  assign _EVAL_4255 = _EVAL_3965 & _EVAL_661;
  assign _EVAL_3335 = 3'h4 | _EVAL_3587;
  assign _EVAL_4717 = {_EVAL_1999,_EVAL_1515};
  assign _EVAL_4642 = {{1'd0}, _EVAL_226};
  assign _EVAL_2758 = _EVAL_5052 & _EVAL_3154;
  assign _EVAL_1353 = {1'h0,_EVAL_2308};
  assign _EVAL_5767 = {{6'd0}, _EVAL_1460};
  assign _EVAL_4823 = {1'h0,_EVAL_2301,_EVAL_4296};
  assign _EVAL_533 = _EVAL_3344 ? 1'h0 : 1'h1;
  assign _EVAL_966 = {{6'd0}, _EVAL_5392};
  assign _EVAL_4956 = _EVAL_2683 & _EVAL_4247;
  assign _EVAL_833 = {{6'd0}, _EVAL_1648};
  assign _EVAL_4090 = {1'h0,_EVAL_356,_EVAL_288};
  assign _EVAL_3093 = _EVAL_730 > _EVAL_431;
  assign _EVAL_47 = _EVAL_4572 & _EVAL_1890;
  assign _EVAL_238 = {_EVAL_5813,_EVAL_5697};
  assign _EVAL_5022 = _EVAL_4486 & _EVAL_2756;
  assign _EVAL_3963 = {_EVAL_1779,_EVAL_164};
  assign _EVAL_5321 = {1'h0,_EVAL_2583};
  assign _EVAL_5805 = _EVAL_1054 ? _EVAL_6013 : _EVAL_2147;
  assign _EVAL_1737 = _EVAL_5899 > _EVAL_858;
  assign _EVAL_673 = _EVAL_325 == 22'h0;
  assign _EVAL_1623 = _EVAL_278 ? _EVAL_2664 : _EVAL_3788;
  assign _EVAL_343 = _EVAL_2636 > _EVAL_5334;
  assign _EVAL_1330 = {1'h0,_EVAL_2422};
  assign _EVAL_5961 = {{6'd0}, _EVAL_5820};
  assign _EVAL_2234 = {_EVAL_1289,28'hf000000};
  assign _EVAL_1148 = 10'h29a == _EVAL_5757;
  assign _EVAL_1821 = _EVAL_4452 ? _EVAL_2263 : _EVAL_4853;
  assign _EVAL_1123 = 4'h8 | _EVAL_4595;
  assign _EVAL_5793 = {_EVAL_2760,_EVAL_5962};
  assign _EVAL_1874 = 2'h2 | _EVAL_2739;
  assign _EVAL_5627 = _EVAL_6052 & _EVAL_3487;
  assign _EVAL_1632 = _EVAL_3979 ? _EVAL_3148 : _EVAL_2747;
  assign _EVAL_4107 = {1'h0,_EVAL_4007};
  assign _EVAL_3711 = {{6'd0}, _EVAL_3527};
  assign _EVAL_2447 = _EVAL_4226 ? _EVAL_5295 : _EVAL_1425;
  assign _EVAL_5253 = _EVAL_520 ? _EVAL_673 : _EVAL_524;
  assign _EVAL_930 = _EVAL_1517 > _EVAL_3823;
  assign _EVAL_1191 = _EVAL_4754 > _EVAL_5719;
  assign _EVAL_2309 = {1'h0,1'h0,_EVAL_1573};
  assign _EVAL_5658 = {1'h0,_EVAL_3634,_EVAL_5949};
  assign _EVAL_3035 = {_EVAL_5046,_EVAL_1440};
  assign _EVAL_3278 = _EVAL_5951 & _EVAL_747;
  assign _EVAL_5841 = _EVAL_1075 & _EVAL_2756;
  assign _EVAL_5290 = {_EVAL_3641,_EVAL_3310};
  assign _EVAL_5221 = _EVAL_2728 & _EVAL_5871;
  assign _EVAL_3422 = _EVAL_1403 & _EVAL_1937;
  assign _EVAL_5861 = {{6'd0}, _EVAL_2995};
  assign _EVAL_1339 = {_EVAL_4968,_EVAL_653};
  assign _EVAL_2840 = {{6'd0}, _EVAL_5552};
  assign _EVAL_1598 = 10'h100 == _EVAL_5757;
  assign _EVAL_3516 = _EVAL_1396 & _EVAL_1293;
  assign _EVAL_4530 = _EVAL_1423 ? _EVAL_3368 : _EVAL_2774;
  assign _EVAL_1566 = _EVAL_1656 ? _EVAL_6031 : _EVAL_5290;
  assign _EVAL_2448 = {1'h0,_EVAL_1831,_EVAL_3846};
  assign _EVAL_3591 = 10'h25e == _EVAL_5757;
  assign _EVAL_1540 = {_EVAL_5142,4'hf,_EVAL_3722,4'hf,_EVAL_2490,4'hf,_EVAL_4416,4'hf};
  assign _EVAL_4417 = {1'h0,_EVAL_1875,_EVAL_394};
  assign _EVAL_5552 = {1'h0,_EVAL_2910,_EVAL_717};
  assign _EVAL_5407 = {1'h0,_EVAL_1147,_EVAL_1101};
  assign _EVAL_4344 = _EVAL_5411 & _EVAL_2162;
  assign _EVAL_3336 = _EVAL_2954 & _EVAL_3154;
  assign _EVAL_5706 = 5'h10 | _EVAL_5562;
  assign _EVAL_2786 = _EVAL_1621 ? {{1'd0}, _EVAL_5485} : _EVAL_3042;
  assign _EVAL_444 = _EVAL_3989 & _EVAL_3154;
  assign _EVAL_2369 = 10'h253 == _EVAL_5757;
  assign _EVAL_1114 = 5'h10 | _EVAL_4943;
  assign _EVAL_3614 = {{6'd0}, _EVAL_3560};
  assign _EVAL_1626 = _EVAL_5220 > _EVAL_4229;
  assign _EVAL_4000 = {{1'd0}, _EVAL_805};
  assign _EVAL_750 = {1'h0,_EVAL_5741,_EVAL_662};
  assign _EVAL_2259 = _EVAL_1347 & _EVAL_3154;
  assign _EVAL_186 = {1'h0,_EVAL_6098,_EVAL_4148};
  assign _EVAL_2316 = 10'h263 == _EVAL_5757;
  assign _EVAL_1953 = {{6'd0}, _EVAL_2722};
  assign _EVAL_639 = {1'h0,_EVAL_887,_EVAL_5655};
  assign _EVAL_5459 = _EVAL_675 ? _EVAL_673 : _EVAL_3253;
  assign _EVAL_1609 = _EVAL_1900 ? _EVAL_5011 : _EVAL_3037;
  assign _EVAL_3289 = _EVAL_2218[55:48];
  assign _EVAL_915 = _EVAL_2596 ? _EVAL_953 : _EVAL_5944;
  assign _EVAL_3585 = _EVAL_4331 ? _EVAL_3834 : _EVAL_2055;
  assign _EVAL_2128 = _EVAL_6063 > _EVAL_3963;
  assign _EVAL_367 = _EVAL_6052 & _EVAL_4477;
  assign _EVAL_4672 = _EVAL_729 > _EVAL_5661;
  assign Queue__EVAL_12 = _EVAL_26;
  assign _EVAL_2112 = _EVAL_220 > _EVAL_2385;
  assign _EVAL_4226 = 10'h21c == _EVAL_5757;
  assign _EVAL_5516 = _EVAL_5068[651];
  assign _EVAL_120 = Queue__EVAL_11;
  assign _EVAL_1751 = _EVAL_1156 & _EVAL_673;
  assign _EVAL_4147 = {1'h0,_EVAL_2096};
  assign _EVAL_1205 = {1'h0,_EVAL_3181,_EVAL_4347};
  assign _EVAL_3604 = {1'h0,_EVAL_5608};
  assign _EVAL_548 = _EVAL_2603 ? {{1'd0}, _EVAL_4234} : _EVAL_3125;
  assign _EVAL_4096 = _EVAL_1608 & _EVAL_3487;
  assign _EVAL_525 = {{6'd0}, _EVAL_657};
  assign _EVAL_4863 = 10'hfe == _EVAL_5757;
  assign _EVAL_3646 = _EVAL_5151 & _EVAL_2756;
  assign _EVAL_6060 = _EVAL_2380 & _EVAL_3487;
  assign _EVAL_3824 = 3'h4 | _EVAL_3027;
  assign _EVAL_1571 = _EVAL_5906 ? _EVAL_569 : _EVAL_189;
  assign _EVAL_5382 = _EVAL_5951 & _EVAL_3977;
  assign _EVAL_1423 = _EVAL_3368 > _EVAL_2774;
  assign _EVAL_1648 = {1'h0,_EVAL_603,_EVAL_5554};
  assign _EVAL_2767 = {1'h0,_EVAL_661,_EVAL_848};
  assign _EVAL_1943 = {{6'd0}, _EVAL_4774};
  assign _EVAL_5687 = {1'h0,_EVAL_3197};
  assign _EVAL_3389 = _EVAL_1075 & _EVAL_1937;
  assign _EVAL_2740 = _EVAL_4734 & _EVAL_2350;
  assign _EVAL_5553 = {1'h0,_EVAL_3983,_EVAL_966};
  assign _EVAL_3967 = _EVAL_2155 & _EVAL_417;
  assign _EVAL_4013 = _EVAL_246 & _EVAL_2756;
  assign _EVAL_3443 = _EVAL_5743 & _EVAL_454;
  assign _EVAL_3415 = {1'h0,_EVAL_5924,_EVAL_3711};
  assign _EVAL_672 = _EVAL_823 ? _EVAL_5515 : _EVAL_1566;
  assign _EVAL_4889 = {{1'd0}, _EVAL_1253};
  assign _EVAL_5031 = {{6'd0}, _EVAL_1925};
  assign _EVAL_2418 = {1'h0,_EVAL_1383,_EVAL_2981};
  assign _EVAL_3633 = {1'h0,1'h0,_EVAL_2157};
  assign _EVAL_3741 = _EVAL_1486 ? _EVAL_609 : _EVAL_3930;
  assign _EVAL_4168 = _EVAL_1477 & _EVAL_3487;
  assign _EVAL_3671 = 10'h241 == _EVAL_5757;
  assign _EVAL_4165 = {_EVAL_4929,_EVAL_2393};
  assign _EVAL_4098 = {{6'd0}, _EVAL_3018};
  assign _EVAL_614 = {{6'd0}, _EVAL_749};
  assign _EVAL_1031 = _EVAL_2910 & _EVAL_582;
  assign _EVAL_1208 = {{6'd0}, _EVAL_2765};
  assign _EVAL_3772 = _EVAL_5547 > _EVAL_4182;
  assign _EVAL_5738 = _EVAL_3293 ? {{1'd0}, _EVAL_3916} : 2'h3;
  assign _EVAL_4032 = _EVAL_2316 ? _EVAL_673 : _EVAL_215;
  assign _EVAL_1172 = {1'h0,_EVAL_4085,_EVAL_1192};
  assign _EVAL_3544 = _EVAL_5951 & _EVAL_4992;
  assign _EVAL_1502 = _EVAL_3270 > _EVAL_5231;
  assign _EVAL_5275 = 10'h25f == _EVAL_5757;
  assign _EVAL_5106 = {{6'd0}, _EVAL_4286};
  assign _EVAL_5581 = 2'h2 | _EVAL_5426;
  assign _EVAL_1390 = 2'h2 | _EVAL_2709;
  assign _EVAL_2841 = _EVAL_4843 & _EVAL_5190;
  assign _EVAL_3851 = {_EVAL_3044,_EVAL_2493};
  assign _EVAL_2159 = _EVAL_3408 ? _EVAL_2848 : _EVAL_672;
  assign _EVAL_5503 = _EVAL_3093 ? _EVAL_730 : _EVAL_431;
  assign _EVAL_1309 = 10'h216 == _EVAL_5757;
  assign _EVAL_2761 = {_EVAL_4164,_EVAL_5142};
  assign _EVAL_4172 = {{6'd0}, _EVAL_5257};
  assign _EVAL_4853 = _EVAL_5792 ? _EVAL_2949 : _EVAL_4805;
  assign _EVAL_5185 = {_EVAL_1444,_EVAL_703};
  assign _EVAL_5660 = {{6'd0}, _EVAL_4238};
  assign _EVAL_3670 = 10'h262 == _EVAL_5757;
  assign _EVAL_433 = _EVAL_5951 & _EVAL_5984;
  assign _EVAL_4894 = _EVAL_2369 ? _EVAL_673 : _EVAL_3619;
  assign _EVAL_4352 = {_EVAL_1278,_EVAL_563};
  assign _EVAL_4074 = _EVAL_5762 ? _EVAL_673 : _EVAL_1848;
  assign _EVAL_5045 = _EVAL_5803 > _EVAL_1284;
  assign _EVAL_4740 = _EVAL_1191 ? _EVAL_4754 : _EVAL_5719;
  assign _EVAL_3645 = {{6'd0}, _EVAL_2971};
  assign _EVAL_4037 = {1'h0,_EVAL_5104};
  assign _EVAL_605 = {{6'd0}, _EVAL_4004};
  assign _EVAL_5073 = _EVAL_5951 & _EVAL_5582;
  assign _EVAL_2527 = _EVAL_1437 ? 1'h0 : 1'h1;
  assign _EVAL_634 = {_EVAL_1024,_EVAL_2827};
  assign _EVAL_1914 = _EVAL_3293 ? _EVAL_1968 : 5'h0;
  assign _EVAL_5780 = _EVAL_4465 | _EVAL_2499;
  assign _EVAL_447 = {1'h0,_EVAL_4338,_EVAL_1013};
  assign _EVAL_1643 = {_EVAL_4019,4'hf,_EVAL_4711,4'hf,_EVAL_1891,4'hf,_EVAL_4479,4'hf};
  assign _EVAL_3037 = _EVAL_3397 ? _EVAL_3750 : _EVAL_495;
  assign _EVAL_5393 = {{1'd0}, _EVAL_4003};
  assign _EVAL_595 = _EVAL_5048 ? _EVAL_673 : _EVAL_3533;
  assign _EVAL_5901 = _EVAL_2286 ? _EVAL_1953 : _EVAL_4358;
  assign _EVAL_4421 = {_EVAL_3062,4'hf,_EVAL_3108,4'hf,_EVAL_5697,4'hf,_EVAL_703,4'hf};
  assign _EVAL_1230 = 3'h4 | _EVAL_425;
  assign _EVAL_2286 = 10'h24e == _EVAL_5757;
  assign _EVAL_3641 = _EVAL_616 & _EVAL_1826;
  assign _EVAL_2648 = _EVAL_2042 ? _EVAL_673 : _EVAL_2800;
  assign _EVAL_1060 = {1'h0,_EVAL_1407,_EVAL_2282};
  assign _EVAL_4415 = _EVAL_1339 > _EVAL_3599;
  assign _EVAL_1457 = {_EVAL_5682,_EVAL_3676};
  assign _EVAL_2838 = _EVAL_6061 ? 1'h0 : 1'h1;
  assign _EVAL_4250 = 10'h287 == _EVAL_5757;
  assign _EVAL_1812 = {_EVAL_791,_EVAL_3040};
  assign _EVAL_4901 = _EVAL_2717 & _EVAL_3203;
  assign Queue__EVAL_10 = _EVAL_88 == 3'h4;
  assign _EVAL_3810 = Queue__EVAL_8[1];
  assign _EVAL_2995 = {1'h0,_EVAL_1506,_EVAL_1892};
  assign _EVAL_723 = _EVAL_5335 ? 1'h0 : 1'h1;
  assign _EVAL_3324 = _EVAL_2855 ? 1'h0 : 1'h1;
  assign _EVAL_3255 = _EVAL_5951 & _EVAL_5115;
  assign _EVAL_6056 = _EVAL_1148 ? _EVAL_673 : _EVAL_5717;
  assign _EVAL_3546 = _EVAL_5951 & _EVAL_3298;
  assign _EVAL_4162 = _EVAL_5068[595];
  assign _EVAL_4864 = {_EVAL_3475,_EVAL_3062};
  assign Queue__EVAL_6 = _EVAL_112;
  assign _EVAL_858 = {_EVAL_4882,_EVAL_4624};
  assign _EVAL_1613 = _EVAL_5951 & _EVAL_2377;
  assign _EVAL_2406 = _EVAL_5615 & _EVAL_4247;
  assign _EVAL_1714 = _EVAL_5068[647];
  assign _EVAL_4769 = _EVAL_3726 > _EVAL_4858;
  assign _EVAL_188 = {{6'd0}, _EVAL_312};
  assign _EVAL_3207 = _EVAL_4955 & _EVAL_643;
  assign _EVAL_550 = _EVAL_5068[640];
  assign _EVAL_1527 = {{6'd0}, _EVAL_5415};
  assign _EVAL_2055 = {_EVAL_5657,_EVAL_4264};
  assign _EVAL_3233 = _EVAL_2036 ? _EVAL_673 : _EVAL_2098;
  assign _EVAL_5808 = {1'h0,_EVAL_454,_EVAL_3127};
  assign _EVAL_4124 = _EVAL_4699 > _EVAL_2315;
  assign _EVAL_2896 = _EVAL_2566 ? _EVAL_929 : _EVAL_5584;
  assign _EVAL_1779 = _EVAL_277 & _EVAL_3914;
  assign _EVAL_719 = {{6'd0}, _EVAL_1353};
  assign _EVAL_4942 = _EVAL_4045 & _EVAL_506;
  assign _EVAL_2664 = {{6'd0}, _EVAL_2534};
  assign _EVAL_2544 = {_EVAL_3172,4'hf,_EVAL_296,4'hf,_EVAL_4264,4'hf,_EVAL_1356,4'hf};
  assign _EVAL_5548 = _EVAL_5951 & _EVAL_2661;
  assign _EVAL_2981 = {{6'd0}, _EVAL_4307};
  assign _EVAL_4177 = _EVAL_3685 > _EVAL_2359;
  assign _EVAL_4903 = 2'h2 | _EVAL_890;
  assign _EVAL_4778 = 10'h244 == _EVAL_5757;
  assign _EVAL_3200 = _EVAL_5068[602];
  assign _EVAL_3395 = _EVAL_1148 ? _EVAL_2544 : _EVAL_261;
  assign _EVAL_3527 = {1'h0,_EVAL_5147};
  assign _EVAL_6091 = {{1'd0}, _EVAL_3483};
  assign _EVAL_1130 = {{1'd0}, _EVAL_689};
  assign _EVAL_195 = _EVAL_5275 ? _EVAL_673 : _EVAL_4074;
  assign _EVAL_4284 = _EVAL_785 ? _EVAL_673 : _EVAL_3675;
  assign _EVAL_5545 = {_EVAL_1255,_EVAL_2889};
  assign _EVAL_5012 = _EVAL_1726 & _EVAL_4477;
  assign _EVAL_5511 = _EVAL_3100 & _EVAL_673;
  assign _EVAL_5265 = {{6'd0}, _EVAL_3633};
  assign _EVAL_400 = _EVAL_2352 ? {{1'd0}, _EVAL_723} : _EVAL_3383;
  assign _EVAL_1799 = {_EVAL_1031,_EVAL_1028};
  assign _EVAL_5038 = _EVAL_2036 ? _EVAL_5224 : _EVAL_313;
  assign _EVAL_1425 = _EVAL_5399 ? _EVAL_2811 : _EVAL_5817;
  assign _EVAL_3090 = _EVAL_4469 ? _EVAL_673 : _EVAL_2648;
  assign _EVAL_4437 = _EVAL_4653 & _EVAL_4477;
  assign _EVAL_855 = _EVAL_3752 ? 1'h0 : 1'h1;
  assign _EVAL_1110 = {1'h0,_EVAL_277,_EVAL_3614};
  assign _EVAL_4590 = {{6'd0}, _EVAL_1803};
  assign _EVAL_4554 = _EVAL_4653 & _EVAL_3487;
  assign _EVAL_2115 = {_EVAL_2815,_EVAL_3771};
  assign _EVAL_5536 = {1'h0,_EVAL_4742,_EVAL_719};
  assign _EVAL_4480 = _EVAL_5163 & _EVAL_2357;
  assign _EVAL_2450 = {{6'd0}, _EVAL_443};
  assign _EVAL_4438 = _EVAL_1537 ? _EVAL_3102 : _EVAL_545;
  assign _EVAL_3446 = _EVAL_1788 ? 1'h0 : 1'h1;
  assign _EVAL_1153 = 10'h21f == _EVAL_5757;
  assign _EVAL_736 = {{1'd0}, _EVAL_5738};
  assign _EVAL_5267 = _EVAL_5068[579];
  assign Queue__EVAL_7 = _EVAL_106;
  assign _EVAL_4660 = {1'h0,_EVAL_1206,_EVAL_815};
  assign _EVAL_5358 = {{6'd0}, _EVAL_2196};
  assign _EVAL_1761 = _EVAL_1320 & _EVAL_673;
  assign _EVAL_3739 = _EVAL_5249 & _EVAL_2690;
  assign _EVAL_3205 = _EVAL_5935 ? 1'h0 : 1'h1;
  assign _EVAL_883 = _EVAL_4345 ? _EVAL_430 : _EVAL_4165;
  assign _EVAL_1320 = _EVAL_5951 & _EVAL_3211;
  assign _EVAL_2637 = {{6'd0}, _EVAL_5536};
  assign _EVAL_4754 = _EVAL_219 ? _EVAL_634 : _EVAL_5923;
  assign _EVAL_4542 = {{6'd0}, _EVAL_161};
  assign _EVAL_1552 = {1'h0,_EVAL_4807,_EVAL_2637};
  assign _EVAL_522 = 2'h2 | _EVAL_1303;
  assign _EVAL_1922 = _EVAL_3639 & _EVAL_2828;
  assign _EVAL_3936 = _EVAL_3039 ? _EVAL_5248 : _EVAL_4520;
  assign _EVAL_4977 = {1'h0,_EVAL_1820,_EVAL_1295};
  assign _EVAL_3463 = {{6'd0}, _EVAL_1987};
  assign _EVAL_4467 = _EVAL_2086 & _EVAL_1618;
  assign _EVAL_2029 = _EVAL_5683 ? {{1'd0}, _EVAL_1042} : _EVAL_5270;
  assign _EVAL_5014 = _EVAL_4010 & _EVAL_4477;
  assign _EVAL_2636 = _EVAL_4809 ? _EVAL_2824 : _EVAL_3353;
  assign _EVAL_219 = _EVAL_634 > _EVAL_5923;
  assign _EVAL_5198 = _EVAL_1381 ? {{1'd0}, _EVAL_2446} : _EVAL_4903;
  assign _EVAL_4446 = _EVAL_5258 ? _EVAL_2450 : _EVAL_2099;
  assign _EVAL_1770 = 10'h2a0 == _EVAL_5757;
  assign _EVAL_1239 = {1'h0,_EVAL_4184,_EVAL_5698};
  assign _EVAL_604 = 5'h10 | _EVAL_2994;
  assign _EVAL_1284 = {_EVAL_2841,_EVAL_5389};
  assign _EVAL_5363 = _EVAL_5615 & _EVAL_5871;
  assign _EVAL_5186 = {1'h0,_EVAL_906,_EVAL_4569};
  assign _EVAL_3487 = _EVAL_1159[0];
  assign _EVAL_3341 = _EVAL_5951 & _EVAL_543;
  assign _EVAL_4217 = {{6'd0}, _EVAL_3415};
  assign _EVAL_4297 = _EVAL_880 & _EVAL_3584;
  assign _EVAL_1181 = {1'h0,_EVAL_2905};
  assign _EVAL_728 = {{1'd0}, _EVAL_615};
  assign _EVAL_4123 = {1'h0,_EVAL_5409,_EVAL_3149};
  assign _EVAL_1710 = _EVAL_4410 ? _EVAL_1712 : _EVAL_705;
  assign _EVAL_1278 = _EVAL_2988 & _EVAL_3001;
  assign _EVAL_3501 = _EVAL_246 & _EVAL_417;
  assign _EVAL_1669 = _EVAL_3092 & _EVAL_1937;
  assign _EVAL_1472 = _EVAL_3864 ? _EVAL_3903 : _EVAL_3656;
  assign _EVAL_5969 = _EVAL_359 ? 8'hff : 8'h0;
  assign _EVAL_3862 = 2'h2 | _EVAL_1130;
  assign _EVAL_6018 = _EVAL_2743 ? {{1'd0}, _EVAL_5614} : _EVAL_3855;
  assign _EVAL_1803 = {1'h0,_EVAL_2516};
  assign _EVAL_311 = _EVAL_640 ? 1'h0 : 1'h1;
  assign _EVAL_3555 = _EVAL_3765 ? {{1'd0}, _EVAL_592} : _EVAL_852;
  assign _EVAL_2435 = {_EVAL_1351,4'hf,_EVAL_1822,4'hf,_EVAL_702,4'hf,_EVAL_558,4'hf};
  assign _EVAL_5131 = _EVAL_6053 & _EVAL_417;
  assign _EVAL_2474 = _EVAL_433 & _EVAL_673;
  assign _EVAL_2780 = {{6'd0}, _EVAL_3168};
  assign _EVAL_1115 = _EVAL_4396 ? _EVAL_673 : _EVAL_3031;
  assign _EVAL_1337 = _EVAL_1430 ? _EVAL_1216 : _EVAL_5504;
  assign _EVAL_4982 = {{6'd0}, _EVAL_4037};
  assign _EVAL_499 = {1'h0,_EVAL_2203,_EVAL_5910};
  assign _EVAL_3190 = _EVAL_1686 | _EVAL_404;
  assign _EVAL_1656 = _EVAL_6031 > _EVAL_5290;
  assign _EVAL_2166 = _EVAL_5413 > _EVAL_1688;
  assign _EVAL_852 = 3'h4 | _EVAL_3064;
  assign _EVAL_4136 = _EVAL_4116 ? _EVAL_673 : _EVAL_4349;
  assign _EVAL_5203 = _EVAL_5068[664];
  assign _EVAL_1013 = {{6'd0}, _EVAL_6016};
  assign _EVAL_5432 = _EVAL_3255 & _EVAL_673;
  assign _EVAL_4816 = _EVAL_1135 ? _EVAL_1414 : _EVAL_853;
  assign _EVAL_4902 = _EVAL_5806 ? _EVAL_673 : _EVAL_4012;
  assign _EVAL_3096 = 2'h2 | _EVAL_4642;
  assign _EVAL_5683 = _EVAL_995 > _EVAL_4354;
  assign _EVAL_4959 = _EVAL_1825 & _EVAL_2756;
  assign _EVAL_1184 = _EVAL_5202[3:0];
  assign _EVAL_163 = 10'h200 == _EVAL_5757;
  assign _EVAL_3318 = _EVAL_1132 & _EVAL_673;
  assign _EVAL_5095 = _EVAL_3419 ? _EVAL_3482 : _EVAL_2319;
  assign _EVAL_1857 = _EVAL_3921 ? _EVAL_1220 : _EVAL_3395;
  assign _EVAL_5145 = _EVAL_3131 > _EVAL_1576;
  assign _EVAL_5487 = {1'h0,_EVAL_4955};
  assign _EVAL_718 = {{6'd0}, _EVAL_3017};
  assign _EVAL_4995 = _EVAL_2714 ? _EVAL_3102 : _EVAL_3452;
  assign _EVAL_1883 = {1'h0,_EVAL_3580};
  assign _EVAL_3273 = _EVAL_5951 & _EVAL_1762;
  assign _EVAL_2415 = {{6'd0}, _EVAL_5746};
  assign _EVAL_5333 = {1'h0,_EVAL_1187};
  assign _EVAL_5322 = _EVAL_4769 ? _EVAL_3726 : _EVAL_4858;
  assign _EVAL_2508 = {{6'd0}, _EVAL_186};
  assign _EVAL_3775 = _EVAL_5951 & _EVAL_2693;
  assign _EVAL_3915 = {1'h0,_EVAL_2825,_EVAL_4098};
  assign _EVAL_5140 = _EVAL_5777 ? {{8'd0}, _EVAL_605} : _EVAL_2365;
  assign _EVAL_4482 = _EVAL_3317 ? {{1'd0}, _EVAL_2978} : _EVAL_5706;
  assign _EVAL_2289 = _EVAL_2633 & _EVAL_2756;
  assign _EVAL_675 = 10'h251 == _EVAL_5757;
  assign _EVAL_707 = _EVAL_4199 ? _EVAL_3045 : _EVAL_1680;
  assign _EVAL_283 = _EVAL_2621 & _EVAL_4477;
  assign _EVAL_6042 = _EVAL_6073 & _EVAL_3154;
  assign _EVAL_1308 = {_EVAL_3449,4'hf,_EVAL_5080,4'hf,_EVAL_531,4'hf,_EVAL_3005,4'hf};
  assign _EVAL_3871 = {1'h0,_EVAL_560,_EVAL_4105};
  assign _EVAL_1827 = _EVAL_1775[31:24];
  assign _EVAL_2696 = {{1'd0}, _EVAL_2029};
  assign _EVAL_2819 = {_EVAL_3094,_EVAL_2561};
  assign _EVAL_4878 = _EVAL_5608 & _EVAL_3589;
  assign _EVAL_5719 = _EVAL_2638 ? _EVAL_3144 : _EVAL_4026;
  assign _EVAL_4523 = 10'h222 == _EVAL_5757;
  assign _EVAL_4015 = 10'h20e == _EVAL_5757;
  assign _EVAL_1791 = {1'h0,_EVAL_3456,_EVAL_525};
  assign _EVAL_4195 = {1'h0,_EVAL_2154,_EVAL_2996};
  assign _EVAL_2004 = 3'h4 | _EVAL_2696;
  assign _EVAL_5989 = _EVAL_5768 | _EVAL_4708;
  assign _EVAL_2330 = {1'h0,_EVAL_4053,_EVAL_4954};
  assign _EVAL_3355 = {{6'd0}, _EVAL_5859};
  assign _EVAL_5109 = _EVAL_1054 ? _EVAL_673 : _EVAL_1154;
  assign _EVAL_3623 = _EVAL_1935 ? _EVAL_3115 : _EVAL_2447;
  assign _EVAL_2094 = {{6'd0}, _EVAL_232};
  assign _EVAL_4973 = {_EVAL_2503,_EVAL_5518};
  assign _EVAL_2206 = {_EVAL_737,4'hf,_EVAL_2629,4'hf,_EVAL_5665,4'hf,_EVAL_5039,4'hf};
  assign _EVAL_5870 = _EVAL_988 ? _EVAL_986 : _EVAL_255;
  assign _EVAL_1465 = _EVAL_5068[661];
  assign _EVAL_2765 = {1'h0,_EVAL_5369};
  assign _EVAL_5453 = _EVAL_4127 ? _EVAL_6079 : _EVAL_3623;
  assign _EVAL_5350 = _EVAL_3814 & _EVAL_2756;
  assign _EVAL_1744 = {1'h0,_EVAL_3133,_EVAL_3343};
  assign _EVAL_724 = _EVAL_796 & _EVAL_3154;
  assign _EVAL_2864 = _EVAL_5068[650];
  assign _EVAL_824 = _EVAL_5315 & _EVAL_2291;
  assign _EVAL_4849 = _EVAL_2046 ? _EVAL_673 : _EVAL_5143;
  assign _EVAL_2813 = _EVAL_3325 ? 1'h0 : 1'h1;
  assign _EVAL_2701 = _EVAL_1630 & _EVAL_673;
  assign _EVAL_6052 = _EVAL_611 & _EVAL_673;
  assign _EVAL_5871 = _EVAL_3048 == 8'hff;
  assign _EVAL_6025 = 10'h20d == _EVAL_5757;
  assign _EVAL_1659 = _EVAL_5951 & _EVAL_1714;
  assign _EVAL_5263 = _EVAL_3717 ? _EVAL_4376 : _EVAL_295;
  assign _EVAL_4992 = _EVAL_5068[603];
  assign _EVAL_359 = Queue__EVAL_4[0];
  assign _EVAL_5577 = _EVAL_5951 & _EVAL_4167;
  assign _EVAL_4578 = _EVAL_2473 ? _EVAL_673 : _EVAL_2779;
  assign _EVAL_5463 = _EVAL_3317 ? _EVAL_349 : _EVAL_3393;
  assign _EVAL_5462 = _EVAL_160 ? _EVAL_673 : _EVAL_2477;
  assign _EVAL_918 = {1'h0,_EVAL_2360,_EVAL_5031};
  assign _EVAL_1693 = {1'h0,_EVAL_4965,_EVAL_4490};
  assign _EVAL_3438 = _EVAL_1726 & _EVAL_3487;
  assign _EVAL_4340 = _EVAL_5951 & _EVAL_4441;
  assign _EVAL_1790 = _EVAL_5472 & _EVAL_673;
  assign _EVAL_5334 = _EVAL_5751 ? _EVAL_3906 : _EVAL_2805;
  assign _EVAL_677 = {1'h0,_EVAL_1301,_EVAL_5934};
  assign _EVAL_4622 = {{6'd0}, _EVAL_3885};
  assign _EVAL_4003 = _EVAL_1866 ? 1'h0 : 1'h1;
  assign _EVAL_174 = _EVAL_5339 & _EVAL_847;
  assign _EVAL_4466 = _EVAL_2852 ? _EVAL_673 : 1'h1;
  assign _EVAL_3383 = 2'h2 | _EVAL_2559;
  assign _EVAL_2943 = _EVAL_1486 ? _EVAL_673 : _EVAL_3304;
  assign _EVAL_1834 = _EVAL_2155 & _EVAL_2350;
  assign _EVAL_4197 = {{6'd0}, _EVAL_3254};
  assign _EVAL_5519 = Queue__EVAL_4[1];
  assign _EVAL_245 = _EVAL_1147 & _EVAL_4065;
  assign _EVAL_4262 = _EVAL_3397 ? {{1'd0}, _EVAL_311} : _EVAL_4321;
  assign _EVAL_1011 = _EVAL_2218[7:0];
  assign _EVAL_518 = {{6'd0}, _EVAL_4763};
  assign _EVAL_902 = _EVAL_1135 ? {{1'd0}, _EVAL_3428} : _EVAL_1123;
  assign _EVAL_5174 = _EVAL_960 & _EVAL_1333;
  assign _EVAL_426 = {1'h0,_EVAL_1240};
  assign _EVAL_158 = _EVAL_5314 & _EVAL_847;
  assign _EVAL_1997 = {_EVAL_2130,_EVAL_3256};
  assign _EVAL_5875 = {1'h0,_EVAL_2009,_EVAL_3549};
  assign _EVAL_2797 = {{6'd0}, _EVAL_5658};
  assign _EVAL_1577 = _EVAL_501 ? _EVAL_285 : _EVAL_3023;
  assign _EVAL_1435 = _EVAL_4015 ? _EVAL_1617 : _EVAL_4446;
  assign _EVAL_602 = {_EVAL_245,_EVAL_1828};
  assign _EVAL_4650 = _EVAL_2701 & _EVAL_2756;
  assign _EVAL_3541 = {{1'd0}, _EVAL_3324};
  assign _EVAL_1749 = _EVAL_4448 ? _EVAL_673 : _EVAL_2461;
  assign _EVAL_1430 = _EVAL_1216 > _EVAL_5504;
  assign _EVAL_2400 = _EVAL_5758 & _EVAL_847;
  assign _EVAL_5377 = {{6'd0}, _EVAL_3806};
  assign _EVAL_2109 = {{1'd0}, _EVAL_992};
  assign _EVAL_1192 = {{6'd0}, _EVAL_4256};
  assign _EVAL_5949 = {{6'd0}, _EVAL_1886};
  assign _EVAL_2549 = {{6'd0}, _EVAL_5533};
  assign _EVAL_2635 = _EVAL_597 & _EVAL_3154;
  assign _EVAL_3752 = _EVAL_4827 > _EVAL_3469;
  assign _EVAL_2737 = _EVAL_4734 & _EVAL_1937;
  assign _EVAL_1637 = _EVAL_4588 & _EVAL_5345;
  assign _EVAL_1886 = {1'h0,_EVAL_5985};
  assign _EVAL_960 = _EVAL_5951 & _EVAL_5800;
  assign _EVAL_1228 = _EVAL_4064 > _EVAL_1904;
  assign intsink__EVAL_1 = _EVAL_24;
  assign _EVAL_624 = _EVAL_4338 & _EVAL_5735;
  assign _EVAL_3039 = 10'h28f == _EVAL_5757;
  assign _EVAL_2244 = _EVAL_4653 & _EVAL_847;
  assign _EVAL_782 = _EVAL_4735 | _EVAL_3390;
  assign _EVAL_232 = {1'h0,_EVAL_5249,_EVAL_4905};
  assign _EVAL_1178 = _EVAL_5924 & _EVAL_3789;
  assign _EVAL_1524 = _EVAL_690 & _EVAL_1301;
  assign _EVAL_990 = 4'h8 | _EVAL_2948;
  assign _EVAL_2587 = _EVAL_743 > _EVAL_445;
  assign _EVAL_178 = {{6'd0}, _EVAL_4541};
  assign _EVAL_4719 = {{1'd0}, _EVAL_3929};
  assign _EVAL_2202 = _EVAL_5222 & _EVAL_2756;
  assign _EVAL_2227 = {_EVAL_281,_EVAL_2920};
  assign _EVAL_1216 = {_EVAL_5966,_EVAL_1672};
  assign _EVAL_3092 = _EVAL_3879 & _EVAL_673;
  assign _EVAL_4657 = {_EVAL_2311,_EVAL_3673};
  assign _EVAL_1763 = Queue__EVAL[4:1];
  assign _EVAL_1646 = _EVAL_1248 ? _EVAL_2853 : _EVAL_2248;
  assign _EVAL_5044 = _EVAL_4820 ? _EVAL_2467 : _EVAL_1354;
  assign _EVAL_822 = _EVAL_1336 > _EVAL_5364;
  assign _EVAL_4546 = {{6'd0}, _EVAL_2396};
  assign _EVAL_5579 = {_EVAL_2711,_EVAL_3108};
  assign _EVAL_3726 = _EVAL_795 ? _EVAL_4169 : _EVAL_602;
  assign _EVAL_3779 = {1'h0,_EVAL_3213};
  assign _EVAL_5024 = _EVAL_4807 & _EVAL_2993;
  assign _EVAL_5469 = _EVAL_1761 & _EVAL_4477;
  assign _EVAL_890 = {{1'd0}, _EVAL_5983};
  assign _EVAL_3064 = {{1'd0}, _EVAL_1264};
  assign _EVAL_3230 = _EVAL_5068[594];
  assign _EVAL_5749 = {{6'd0}, _EVAL_1110};
  assign _EVAL_4638 = {{1'd0}, _EVAL_5403};
  assign _EVAL_3051 = _EVAL_5928 & _EVAL_2350;
  assign _EVAL_805 = _EVAL_2958 ? {{1'd0}, _EVAL_6018} : _EVAL_5171;
  assign _EVAL_3319 = _EVAL_5951 & _EVAL_3535;
  assign _EVAL_5065 = {{6'd0}, _EVAL_2894};
  assign _EVAL_3947 = {{6'd0}, _EVAL_1939};
  assign _EVAL_5995 = 10'h20c == _EVAL_5757;
  assign _EVAL_1923 = {1'h0,_EVAL_4119};
  assign _EVAL_1732 = _EVAL_5951 & _EVAL_1465;
  assign _EVAL_717 = {{6'd0}, _EVAL_2353};
  assign _EVAL_681 = _EVAL_2218[15:8];
  assign _EVAL_2198 = _EVAL_1608 & _EVAL_847;
  assign _EVAL_3419 = 10'h25d == _EVAL_5757;
  assign _EVAL_667 = {1'h0,_EVAL_5558,_EVAL_5378};
  assign _EVAL_5794 = {_EVAL_317,_EVAL_296};
  assign _EVAL_1023 = {_EVAL_2914,_EVAL_2462};
  assign _EVAL_5266 = _EVAL_5068[653];
  assign _EVAL_3732 = {_EVAL_2393,28'hf000000};
  assign _EVAL_1276 = {1'h0,_EVAL_1287,_EVAL_4640};
  assign _EVAL_2591 = 2'h2 | _EVAL_3541;
  assign _EVAL_5013 = _EVAL_4452 ? _EVAL_673 : _EVAL_2764;
  assign _EVAL_3466 = _EVAL_5068[662];
  assign _EVAL_5111 = _EVAL_3450 & _EVAL_3327;
  assign _EVAL_4549 = _EVAL_2566 ? _EVAL_673 : _EVAL_4902;
  assign _EVAL_278 = 10'h203 == _EVAL_5757;
  assign _EVAL_2642 = _EVAL_898 ? {{1'd0}, _EVAL_4687} : _EVAL_1397;
  assign _EVAL_517 = _EVAL_3731 ? 1'h0 : 1'h1;
  assign _EVAL_1271 = _EVAL_1252 ? {{1'd0}, _EVAL_2928} : _EVAL_1417;
  assign _EVAL_5907 = _EVAL_4486 & _EVAL_417;
  assign _EVAL_4458 = _EVAL_2979 ? _EVAL_3128 : _EVAL_3046;
  assign _EVAL_4758 = {1'h0,_EVAL_1041,_EVAL_4426};
  assign _EVAL_5505 = _EVAL_4352 > _EVAL_4657;
  assign _EVAL_4384 = _EVAL_1018 ? _EVAL_673 : _EVAL_3110;
  assign _EVAL_5615 = _EVAL_2189 & _EVAL_673;
  assign _EVAL_3891 = _EVAL_5551 > _EVAL_4474;
  assign _EVAL_472 = _EVAL_2161 ? _EVAL_673 : _EVAL_3233;
  assign _EVAL_4819 = _EVAL_1347 & _EVAL_4477;
  assign _EVAL_5824 = _EVAL_2568 ? _EVAL_763 : _EVAL_3526;
  assign _EVAL_756 = _EVAL_3989 & _EVAL_4477;
  assign _EVAL_2933 = _EVAL_4637 ? _EVAL_673 : _EVAL_3900;
  assign _EVAL_2812 = {_EVAL_1827,_EVAL_166,_EVAL_3674,_EVAL_1282};
  assign _EVAL_2105 = _EVAL_3318 & _EVAL_3487;
  assign _EVAL_1220 = {_EVAL_2462,4'hf,_EVAL_4911,4'hf,_EVAL_1828,4'hf,_EVAL_1442,4'hf};
  assign _EVAL_5348 = _EVAL_5096 & _EVAL_3487;
  assign _EVAL_1496 = {1'h0,_EVAL_644};
  assign _EVAL_733 = {_EVAL_813,_EVAL_2537};
  assign _EVAL_4763 = {1'h0,_EVAL_1671,_EVAL_1759};
  assign _EVAL_5047 = 2'h2 | _EVAL_1124;
  assign _EVAL_3661 = _EVAL_4626 ? _EVAL_3356 : _EVAL_5191;
  assign _EVAL_2176 = _EVAL_5068[601];
  assign _EVAL_3554 = {1'h0,_EVAL_1314,_EVAL_753};
  assign _EVAL_4026 = {_EVAL_3290,_EVAL_3464};
  assign _EVAL_919 = _EVAL_4318 ? _EVAL_276 : _EVAL_4055;
  assign _EVAL_1378 = _EVAL_3496 & _EVAL_673;
  assign _EVAL_5771 = _EVAL_1860 & _EVAL_3154;
  assign _EVAL_5717 = _EVAL_3099 ? _EVAL_673 : _EVAL_1115;
  assign _EVAL_4159 = 10'h210 == _EVAL_5757;
  assign _EVAL_156 = _EVAL_5468 & _EVAL_1937;
  assign _EVAL_2703 = 10'h247 == _EVAL_5757;
  assign _EVAL_687 = _EVAL_4789 ? _EVAL_1738 : _EVAL_4483;
  assign _EVAL_1382 = 10'h246 == _EVAL_5757;
  assign _EVAL_2845 = {1'h0,_EVAL_506,_EVAL_2061};
  assign _EVAL_5637 = _EVAL_5068[515];
  assign _EVAL_2211 = {{6'd0}, _EVAL_6019};
  assign _EVAL_1087 = _EVAL_5068[597];
  assign _EVAL_4445 = 5'h10 | _EVAL_4000;
  assign _EVAL_2590 = _EVAL_1191 ? {{1'd0}, _EVAL_4131} : _EVAL_1970;
  assign _EVAL_5939 = 10'h242 == _EVAL_5757;
  assign _EVAL_1630 = _EVAL_5951 & _EVAL_3985;
  assign _EVAL_4064 = _EVAL_2719 ? _EVAL_2188 : _EVAL_2332;
  assign _EVAL_3642 = _EVAL_4734 & _EVAL_2756;
  assign _EVAL_993 = _EVAL_297 ? {{1'd0}, _EVAL_2212} : _EVAL_5366;
  assign _EVAL_5181 = {1'h0,_EVAL_1510,_EVAL_211};
  assign _EVAL_1292 = _EVAL_3058 == 8'hff;
  assign _EVAL_5062 = _EVAL_5636 ? _EVAL_673 : _EVAL_5563;
  assign _EVAL_1304 = 3'h4 | _EVAL_4249;
  assign _EVAL_3011 = {1'h0,_EVAL_5878,_EVAL_2586};
  assign _EVAL_4476 = _EVAL_5314 & _EVAL_4477;
  assign _EVAL_4198 = Queue__EVAL_8[2];
  assign _EVAL_2747 = _EVAL_1321 ? _EVAL_4663 : _EVAL_1796;
  assign _EVAL_1132 = _EVAL_5951 & _EVAL_234;
  assign _EVAL_5864 = {{6'd0}, _EVAL_2671};
  assign _EVAL_6100 = {_EVAL_4440,_EVAL_899};
  assign _EVAL_2074 = _EVAL_5068[593];
  assign _EVAL_4998 = 2'h2 | _EVAL_4935;
  assign _EVAL_3971 = {1'h0,_EVAL_3887,_EVAL_4718};
  assign _EVAL_5406 = {1'h0,_EVAL_1730,_EVAL_2951};
  assign _EVAL_3016 = _EVAL_5397 ? _EVAL_673 : _EVAL_4549;
  assign _EVAL_4752 = _EVAL_5674 ? {{1'd0}, _EVAL_4945} : _EVAL_4445;
  assign _EVAL_1939 = {1'h0,_EVAL_5002,_EVAL_4919};
  assign _EVAL_4789 = _EVAL_1738 > _EVAL_4483;
  assign _EVAL_3169 = _EVAL_2312 & _EVAL_5300;
  assign _EVAL_4705 = _EVAL_2499 ? _EVAL_1035 : _EVAL_4741;
  assign _EVAL_1829 = _EVAL_2587 ? {{1'd0}, _EVAL_841} : _EVAL_5581;
  assign _EVAL_3576 = {{6'd0}, _EVAL_4360};
  assign _EVAL_1813 = _EVAL_5108 ? _EVAL_6067 : _EVAL_1011;
  assign _EVAL_5759 = _EVAL_1753 & _EVAL_3154;
  assign _EVAL_524 = _EVAL_1614 ? _EVAL_673 : _EVAL_185;
  assign _EVAL_4634 = _EVAL_2568 ? 1'h0 : 1'h1;
  assign _EVAL_5818 = _EVAL_3629 & _EVAL_5309;
  assign _EVAL_230 = _EVAL_795 ? 1'h0 : 1'h1;
  assign _EVAL_1698 = _EVAL_333 ? _EVAL_2801 : _EVAL_1623;
  assign _EVAL_1441 = {_EVAL_4382,_EVAL_3467};
  assign _EVAL_1035 = Queue__EVAL[23:16];
  assign _EVAL_3094 = _EVAL_5741 & _EVAL_2825;
  assign _EVAL_2104 = _EVAL_5763 > _EVAL_4913;
  assign _EVAL_3578 = _EVAL_4469 ? _EVAL_4421 : _EVAL_6082;
  assign _EVAL_664 = _EVAL_4746 ? _EVAL_3465 : _EVAL_5183;
  assign _EVAL_1279 = _EVAL_4863 ? _EVAL_1372 : _EVAL_5770;
  assign _EVAL_4815 = _EVAL_5386 & _EVAL_4443;
  assign _EVAL_3561 = _EVAL_2784 & _EVAL_2350;
  assign _EVAL_1952 = {{6'd0}, _EVAL_5553};
  assign _EVAL_1680 = _EVAL_5256 ? _EVAL_438 : _EVAL_6058;
  assign _EVAL_674 = {_EVAL_4878,_EVAL_3429};
  assign _EVAL_3855 = 3'h4 | _EVAL_1275;
  assign _EVAL_788 = _EVAL_1075 & _EVAL_2350;
  assign _EVAL_4089 = _EVAL_3618 ? _EVAL_1560 : _EVAL_903;
  assign _EVAL_4008 = _EVAL_2595 & _EVAL_2756;
  assign _EVAL_2714 = _EVAL_2728 & _EVAL_3043;
  assign _EVAL_4005 = _EVAL_2233 & _EVAL_1342;
  assign _EVAL_2481 = _EVAL_4835 & _EVAL_673;
  assign _EVAL_848 = {{6'd0}, _EVAL_3612};
  assign _EVAL_2579 = _EVAL_5337 ? _EVAL_2085 : {{17'd0}, _EVAL_3838};
  assign _EVAL_2757 = _EVAL_5951 & _EVAL_4566;
  assign _EVAL_615 = _EVAL_3088 ? 1'h0 : 1'h1;
  assign _EVAL_4734 = _EVAL_3775 & _EVAL_673;
  assign _EVAL_3861 = _EVAL_2486 & _EVAL_2350;
  assign _EVAL_2173 = _EVAL_1321 ? _EVAL_673 : _EVAL_2374;
  assign _EVAL_1416 = {{1'd0}, _EVAL_5967};
  assign _EVAL_3168 = {1'h0,_EVAL_4336,_EVAL_1952};
  assign _EVAL_3120 = {1'h0,_EVAL_2580};
  assign _EVAL_5340 = _EVAL_2857 & _EVAL_4477;
  assign _EVAL_2727 = _EVAL_5939 ? _EVAL_4546 : _EVAL_3291;
  assign _EVAL_3254 = {1'h0,_EVAL_5396,24'h0};
  assign _EVAL_772 = {_EVAL_2141,_EVAL_4040};
  assign _EVAL_5164 = _EVAL_4015 ? _EVAL_673 : _EVAL_2201;
  assign _EVAL_2429 = {{1'd0}, _EVAL_533};
  assign _EVAL_3715 = {1'h0,_EVAL_5163,_EVAL_1740};
  assign _EVAL_4010 = _EVAL_336 & _EVAL_673;
  assign _EVAL_1760 = {{6'd0}, _EVAL_5388};
  assign _EVAL_4266 = {_EVAL_4876,_EVAL_1822};
  assign _EVAL_1498 = _EVAL_4940 ? 1'h0 : 1'h1;
  assign _EVAL_3150 = _EVAL_5951 & _EVAL_5491;
  assign _EVAL_794 = {1'h0,1'h0,_EVAL_5864};
  assign _EVAL_5644 = _EVAL_4252 & _EVAL_673;
  assign _EVAL_6012 = _EVAL_5605 ? _EVAL_673 : _EVAL_4539;
  assign _EVAL_2851 = _EVAL_1765 & _EVAL_3213;
  assign _EVAL_1168 = _EVAL_5873 ? 1'h0 : 1'h1;
  assign _EVAL_916 = _EVAL_5540 & _EVAL_417;
  assign _EVAL_5715 = _EVAL_4606 ? 1'h0 : 1'h1;
  assign _EVAL_3430 = _EVAL_1020 ? _EVAL_772 : _EVAL_1950;
  assign _EVAL_5906 = _EVAL_569 > _EVAL_189;
  assign _EVAL_3717 = _EVAL_4376 > _EVAL_295;
  assign _EVAL_3668 = _EVAL_5951 & _EVAL_2952;
  assign _EVAL_4221 = {1'h0,_EVAL_4291,_EVAL_3330};
  assign _EVAL_929 = {{6'd0}, _EVAL_4860};
  assign _EVAL_3291 = _EVAL_160 ? _EVAL_2279 : _EVAL_5117;
  assign _EVAL_2346 = _EVAL_606 & _EVAL_3912;
  assign _EVAL_1236 = Queue__EVAL_8[8];
  assign _EVAL_2231 = Queue__EVAL[7:4];
  assign _EVAL_2348 = {_EVAL_3479,_EVAL_3743};
  assign _EVAL_2122 = {{6'd0}, _EVAL_4123};
  assign _EVAL_1532 = _EVAL_1477 & _EVAL_3154;
  assign _EVAL_2829 = _EVAL_1378 & _EVAL_2756;
  assign _EVAL_5460 = _EVAL_1382 ? _EVAL_2618 : _EVAL_2143;
  assign _EVAL_1690 = {{6'd0}, _EVAL_1113};
  assign _EVAL_988 = 10'h29e == _EVAL_5757;
  assign _EVAL_593 = {{6'd0}, _EVAL_1258};
  assign _EVAL_4301 = _EVAL_4742 & _EVAL_4397;
  assign _EVAL_3682 = {{6'd0}, _EVAL_4076};
  assign _EVAL_1073 = _EVAL_5928 & _EVAL_2756;
  assign _EVAL_1157 = {2'h0,_EVAL_3945,_EVAL_484};
  assign _EVAL_995 = _EVAL_1654 ? _EVAL_1997 : _EVAL_1221;
  assign _EVAL_1048 = {{6'd0}, _EVAL_5783};
  assign _EVAL_1374 = Queue__EVAL[24];
  assign _EVAL_979 = {1'h0,_EVAL_5940,_EVAL_1208};
  assign _EVAL_3532 = _EVAL_4345 ? {{1'd0}, _EVAL_5323} : 3'h7;
  assign _EVAL_4318 = _EVAL_276 > _EVAL_4055;
  assign _EVAL_4290 = {1'h0,_EVAL_4397,_EVAL_2794};
  assign _EVAL_436 = {1'h0,_EVAL_2918,_EVAL_3355};
  assign _EVAL_4122 = {{1'd0}, _EVAL_4582};
  assign _EVAL_4489 = _EVAL_2929 ? _EVAL_2492 : _EVAL_1827;
  assign _EVAL_892 = _EVAL_5151 & _EVAL_417;
  assign _EVAL_3950 = {{6'd0}, _EVAL_2283};
  assign _EVAL_1112 = _EVAL_782 | _EVAL_1537;
  assign _EVAL_3941 = 10'h289 == _EVAL_5757;
  assign _EVAL_5011 = _EVAL_5815 ? _EVAL_3431 : _EVAL_685;
  assign _EVAL_1503 = {{6'd0}, _EVAL_304};
  assign _EVAL_2081 = _EVAL_4374 & _EVAL_3594;
  assign _EVAL_1678 = _EVAL_675 ? _EVAL_5026 : _EVAL_732;
  assign Queue__EVAL_5 = _EVAL_124;
  assign _EVAL_3191 = {_EVAL_1059,_EVAL_834};
  assign _EVAL_313 = _EVAL_4402 ? _EVAL_4542 : _EVAL_3970;
  assign _EVAL_2951 = {{6'd0}, _EVAL_426};
  assign _EVAL_337 = {1'h0,_EVAL_3196,_EVAL_977};
  assign _EVAL_3222 = Queue__EVAL[16];
  assign _EVAL_903 = _EVAL_1780 ? _EVAL_483 : _EVAL_3937;
  assign _EVAL_1056 = {1'h0,_EVAL_2717,_EVAL_614};
  assign _EVAL_3431 = _EVAL_5505 ? _EVAL_4352 : _EVAL_4657;
  assign _EVAL_349 = _EVAL_3848 ? _EVAL_883 : _EVAL_5359;
  assign _EVAL_3056 = _EVAL_4584 & _EVAL_6098;
  assign _EVAL_5108 = _EVAL_5174 & _EVAL_1292;
  assign _EVAL_4835 = _EVAL_5951 & _EVAL_1352;
  assign _EVAL_2331 = _EVAL_4614 ? 1'h0 : 1'h1;
  assign _EVAL_4646 = {_EVAL_1637,_EVAL_3722};
  assign _EVAL_5324 = _EVAL_5093 ? _EVAL_5106 : _EVAL_1678;
  assign _EVAL_1520 = _EVAL_5617 ? _EVAL_5545 : _EVAL_5373;
  assign _EVAL_4179 = {{6'd0}, _EVAL_5638};
  assign _EVAL_2940 = {{6'd0}, _EVAL_2997};
  assign _EVAL_2417 = _EVAL_2155 & _EVAL_1937;
  assign _EVAL_2047 = {1'h0,_EVAL_3946};
  assign _EVAL_3635 = _EVAL_5951 & _EVAL_4246;
  assign _EVAL_2407 = _EVAL_1726 & _EVAL_3154;
  assign _EVAL_1100 = _EVAL_2474 & _EVAL_2756;
  assign _EVAL_3297 = {{6'd0}, _EVAL_5526};
  assign _EVAL_640 = _EVAL_5185 > _EVAL_238;
  assign _EVAL_199 = _EVAL_5221 ? _EVAL_2492 : _EVAL_4884;
  assign _EVAL_1900 = _EVAL_5011 > _EVAL_3037;
  assign _EVAL_4174 = _EVAL_3318 & _EVAL_847;
  assign _EVAL_2130 = _EVAL_2422 & _EVAL_6030;
  assign _EVAL_759 = _EVAL_1761 & _EVAL_3487;
  assign _EVAL_840 = 2'h2 | _EVAL_5513;
  assign _EVAL_3193 = _EVAL_2177 & _EVAL_1942;
  assign _EVAL_567 = _EVAL_4895 ? _EVAL_2697 : _EVAL_3791;
  assign _EVAL_6044 = {{6'd0}, _EVAL_437};
  assign _EVAL_465 = _EVAL_3215 & _EVAL_1937;
  assign _EVAL_1587 = {4'h0,_EVAL_5311,4'hf};
  assign _EVAL_3416 = {{1'd0}, _EVAL_1885};
  assign _EVAL_3567 = {1'h0,_EVAL_5781};
  assign _EVAL_2470 = _EVAL_459 > _EVAL_2348;
  assign _EVAL_250 = {1'h0,_EVAL_3914,_EVAL_5961};
  assign _EVAL_3934 = _EVAL_5951 & _EVAL_786;
  assign _EVAL_3372 = _EVAL_642 > _EVAL_466;
  assign _EVAL_791 = _EVAL_3983 & _EVAL_1929;
  assign _EVAL_3334 = {{6'd0}, _EVAL_1276};
  assign _EVAL_1967 = Queue__EVAL[8];
  assign _EVAL_1120 = {_EVAL_658,_EVAL_4571};
  assign _EVAL_3756 = _EVAL_3341 & _EVAL_673;
  assign _EVAL_1150 = _EVAL_2912 & _EVAL_2350;
  assign _EVAL_5905 = _EVAL_1159[23:20];
  assign _EVAL_715 = {_EVAL_4571,4'hf,_EVAL_4908,4'hf,_EVAL_1797,4'hf,_EVAL_3538,4'hf};
  assign _EVAL_1569 = _EVAL_5951 & _EVAL_6004;
  assign _EVAL_1817 = 3'h4 | _EVAL_1583;
  assign _EVAL_2056 = {{6'd0}, _EVAL_4036};
  assign _EVAL_5068 = 1024'h1 << _EVAL_5757;
  assign _EVAL_5849 = {1'h0,_EVAL_1602,_EVAL_1771};
  assign _EVAL_4055 = _EVAL_822 ? _EVAL_1336 : _EVAL_5364;
  assign _EVAL_5787 = _EVAL_5951 & _EVAL_3230;
  assign _EVAL_1554 = _EVAL_1020 ? 1'h0 : 1'h1;
  assign _EVAL_2944 = _EVAL_2034 ? _EVAL_2206 : _EVAL_2882;
  assign _EVAL_2997 = {1'h0,_EVAL_5696};
  assign _EVAL_5681 = {_EVAL_2578,_EVAL_4390};
  assign _EVAL_2050 = 10'h24f == _EVAL_5757;
  assign _EVAL_2467 = _EVAL_4606 ? _EVAL_2787 : _EVAL_5325;
  assign _EVAL_4021 = _EVAL_3408 ? {{1'd0}, _EVAL_4534} : _EVAL_4611;
  assign _EVAL_448 = _EVAL_5906 ? {{1'd0}, _EVAL_2120} : _EVAL_3824;
  assign _EVAL_5049 = _EVAL_919 > _EVAL_4816;
  assign _EVAL_1999 = _EVAL_4367 & _EVAL_1188;
  assign _EVAL_2457 = _EVAL_1493 & _EVAL_5985;
  assign _EVAL_138 = {{2'd0}, _EVAL_4791};
  assign _EVAL_5554 = {{6'd0}, _EVAL_1744};
  assign _EVAL_3460 = _EVAL_822 ? {{1'd0}, _EVAL_4752} : _EVAL_1495;
  assign _EVAL_4893 = {_EVAL_1484,4'hf,_EVAL_561,4'hf,_EVAL_2557,4'hf,_EVAL_1676,4'hf};
  assign _EVAL_468 = _EVAL_5794 > _EVAL_4178;
  assign _EVAL_1935 = 10'h21b == _EVAL_5757;
  assign _EVAL_3047 = _EVAL_1159[4:1];
  assign _EVAL_1842 = _EVAL_468 ? 1'h0 : 1'h1;
  assign _EVAL_4580 = {1'h0,_EVAL_2366,_EVAL_1549};
  assign _EVAL_1381 = _EVAL_329 > _EVAL_4530;
  assign _EVAL_4131 = _EVAL_219 ? 1'h0 : 1'h1;
  assign _EVAL_795 = _EVAL_4169 > _EVAL_602;
  assign _EVAL_2398 = _EVAL_278 ? _EVAL_673 : _EVAL_3405;
  assign _EVAL_4267 = {{6'd0}, _EVAL_2418};
  assign _EVAL_1156 = _EVAL_5951 & _EVAL_1699;
  assign _EVAL_2157 = {{6'd0}, _EVAL_794};
  assign _EVAL_1665 = _EVAL_5068[608];
  assign _EVAL_1644 = _EVAL_4250 ? _EVAL_1308 : _EVAL_915;
  assign _EVAL_4403 = _EVAL_943 & _EVAL_236;
  assign _EVAL_3686 = _EVAL_4789 ? 1'h0 : 1'h1;
  assign _EVAL_3330 = {{6'd0}, _EVAL_4147};
  assign _EVAL_4490 = {{6'd0}, _EVAL_4328};
  assign _EVAL_5751 = _EVAL_3906 > _EVAL_2805;
  assign _EVAL_3838 = _EVAL_2852 ? _EVAL_1157 : 7'h0;
  assign _EVAL_5677 = _EVAL_501 ? 1'h0 : 1'h1;
  assign _EVAL_5301 = {1'h0,_EVAL_783};
  assign _EVAL_3763 = _EVAL_5951 & _EVAL_289;
  assign _EVAL_4251 = {{6'd0}, _EVAL_2878};
  assign _EVAL_4919 = {{6'd0}, _EVAL_3907};
  assign _EVAL_576 = _EVAL_2667 & _EVAL_5104;
  assign _EVAL_286 = {1'h0,_EVAL_4612,_EVAL_324};
  assign _EVAL_2139 = {1'h0,_EVAL_2778};
  assign _EVAL_5833 = _EVAL_5113 & _EVAL_2350;
  assign _EVAL_3587 = {{1'd0}, _EVAL_993};
  assign _EVAL_4658 = 3'h4 | _EVAL_736;
  assign _EVAL_5777 = 10'h223 == _EVAL_5757;
  assign _EVAL_443 = {1'h0,_EVAL_3783,_EVAL_5146};
  assign _EVAL_2336 = {1'h0,_EVAL_5101,_EVAL_2122};
  assign _EVAL_4004 = {1'h0,_EVAL_690,_EVAL_1461};
  assign _EVAL_4718 = {{6'd0}, _EVAL_1481};
  assign _EVAL_2020 = _EVAL_2857 & _EVAL_3487;
  assign _EVAL_2856 = {{1'd0}, _EVAL_1164};
  assign _EVAL_3311 = _EVAL_5125 & _EVAL_2350;
  assign _EVAL_3046 = _EVAL_297 ? _EVAL_3796 : _EVAL_700;
  assign _EVAL_165 = {{6'd0}, _EVAL_3733};
  assign _EVAL_5288 = _EVAL_5821 & _EVAL_3487;
  assign _EVAL_430 = _EVAL_5435 ? 5'h10 : _EVAL_5297;
  assign _EVAL_3498 = 10'h280 == _EVAL_5757;
  assign _EVAL_4958 = _EVAL_1668 ? {{1'd0}, _EVAL_4482} : _EVAL_1508;
  assign _EVAL_2228 = {_EVAL_3603,_EVAL_5537};
  assign _EVAL_5716 = _EVAL_5951 & _EVAL_2884;
  assign _EVAL_218 = _EVAL_5429 & _EVAL_673;
  assign _EVAL_3439 = _EVAL_1806 & _EVAL_3154;
  assign _EVAL_1325 = _EVAL_3215 & _EVAL_2756;
  assign _EVAL_853 = _EVAL_4728 ? _EVAL_192 : _EVAL_2522;
  assign _EVAL_5269 = _EVAL_5068[643];
  assign _EVAL_3619 = _EVAL_835 ? _EVAL_673 : _EVAL_3667;
  assign _EVAL_2421 = _EVAL_5052 & _EVAL_4477;
  assign _EVAL_5769 = _EVAL_5951 & _EVAL_5782;
  assign _EVAL_942 = _EVAL_4633 > _EVAL_2610;
  assign _EVAL_5030 = _EVAL_4486 & _EVAL_1937;
  assign _EVAL_4414 = _EVAL_2621 & _EVAL_3154;
  assign _EVAL_4088 = Queue__EVAL[15:12];
  assign _EVAL_1956 = _EVAL_5951 & _EVAL_5269;
  assign _EVAL_2929 = _EVAL_2683 & _EVAL_5871;
  assign _EVAL_2188 = {_EVAL_3644,_EVAL_4786};
  assign _EVAL_5426 = {{1'd0}, _EVAL_2331};
  assign _EVAL_2287 = _EVAL_4412 ? 1'h0 : 1'h1;
  assign _EVAL_4012 = _EVAL_4337 ? _EVAL_673 : _EVAL_5872;
  assign _EVAL_406 = _EVAL_1121 & _EVAL_5916;
  assign _EVAL_5748 = _EVAL_4944 & _EVAL_4103;
  assign _EVAL_1101 = {{6'd0}, _EVAL_2139};
  assign _EVAL_2779 = _EVAL_1382 ? _EVAL_673 : _EVAL_5332;
  assign _EVAL_3788 = _EVAL_3146 ? _EVAL_5749 : _EVAL_3606;
  assign _EVAL_3405 = _EVAL_3146 ? _EVAL_673 : _EVAL_472;
  assign _EVAL_1113 = {1'h0,_EVAL_5521,_EVAL_5467};
  assign _EVAL_4148 = {{6'd0}, _EVAL_4237};
  assign _EVAL_5899 = {_EVAL_3193,_EVAL_5009};
  assign _EVAL_3848 = _EVAL_883 > _EVAL_5359;
  assign _EVAL_1901 = _EVAL_5222 & _EVAL_417;
  assign _EVAL_2190 = 10'h28e == _EVAL_5757;
  assign _EVAL_5468 = _EVAL_850 & _EVAL_673;
  assign _EVAL_5294 = _EVAL_1347 & _EVAL_3487;
  assign _EVAL_3149 = {{6'd0}, _EVAL_693};
  assign _EVAL_5801 = _EVAL_5951 & _EVAL_3564;
  assign _EVAL_5557 = _EVAL_2728 & _EVAL_1292;
  assign _EVAL_5612 = _EVAL_3899 ? _EVAL_2492 : _EVAL_1106;
  assign _EVAL_4805 = _EVAL_4116 ? _EVAL_2024 : _EVAL_1644;
  assign _EVAL_3872 = _EVAL_4626 ? _EVAL_673 : _EVAL_432;
  assign _EVAL_6101 = _EVAL_4620 & _EVAL_560;
  assign _EVAL_1410 = _EVAL_393 ? _EVAL_673 : _EVAL_4384;
  assign _EVAL_49 = intsink__EVAL_0;
  assign _EVAL_1354 = _EVAL_1437 ? _EVAL_368 : _EVAL_5098;
  assign _EVAL_1551 = _EVAL_356 & _EVAL_1671;
  assign _EVAL_823 = _EVAL_5515 > _EVAL_1566;
  assign _EVAL_485 = _EVAL_5951 & _EVAL_5405;
  assign _EVAL_3102 = Queue__EVAL[15:8];
  assign _EVAL_5089 = 10'h258 == _EVAL_5757;
  assign _EVAL_5113 = _EVAL_3217 & _EVAL_673;
  assign _EVAL_1409 = _EVAL_4556 & _EVAL_417;
  assign _EVAL_3895 = _EVAL_4177 ? {{1'd0}, _EVAL_1129} : _EVAL_1298;
  assign _EVAL_3128 = _EVAL_5120 ? _EVAL_5952 : _EVAL_5503;
  assign _EVAL_3977 = _EVAL_5068[657];
  assign _EVAL_3625 = {{1'd0}, _EVAL_6078};
  assign _EVAL_315 = _EVAL_3092 & _EVAL_2350;
  assign _EVAL_5373 = {_EVAL_1215,_EVAL_3173};
  assign _EVAL_958 = _EVAL_3498 ? _EVAL_2234 : _EVAL_1315;
  assign _EVAL_3428 = _EVAL_2166 ? {{1'd0}, _EVAL_4829} : _EVAL_1662;
  assign _EVAL_3442 = _EVAL_6025 ? _EVAL_673 : _EVAL_5164;
  assign _EVAL_2788 = {_EVAL_5748,_EVAL_561};
  assign _EVAL_1032 = _EVAL_3191 > _EVAL_2115;
  assign _EVAL_3865 = _EVAL_5777 ? _EVAL_673 : _EVAL_4401;
  assign _EVAL_5619 = _EVAL_2954 & _EVAL_3487;
  assign _EVAL_3637 = _EVAL_1248 ? _EVAL_673 : _EVAL_2823;
  assign _EVAL_4941 = {1'h0,_EVAL_3234,_EVAL_2337};
  assign _EVAL_2477 = _EVAL_4778 ? _EVAL_673 : _EVAL_4578;
  assign _EVAL_5166 = {_EVAL_4255,_EVAL_531};
  assign _EVAL_2895 = _EVAL_4007 & _EVAL_1641;
  assign _EVAL_2802 = _EVAL_4396 ? _EVAL_1643 : _EVAL_3059;
  assign _EVAL_4337 = 10'h25c == _EVAL_5757;
  assign _EVAL_1397 = 4'h8 | _EVAL_1433;
  assign _EVAL_6092 = _EVAL_5540 & _EVAL_2756;
  assign _EVAL_689 = _EVAL_912 ? 1'h0 : 1'h1;
  assign _EVAL_2365 = _EVAL_2101 ? _EVAL_718 : _EVAL_4906;
  assign _EVAL_5359 = _EVAL_3905 ? _EVAL_3877 : _EVAL_1914;
  assign _EVAL_969 = 4'h8 | _EVAL_5918;
  assign _EVAL_4913 = _EVAL_2342 ? _EVAL_4387 : _EVAL_3893;
  assign Queue__EVAL_13 = _EVAL_24;
  assign _EVAL_5188 = _EVAL_3756 & _EVAL_2756;
  assign _EVAL_3275 = _EVAL_5335 ? _EVAL_3851 : _EVAL_5480;
  assign _EVAL_697 = _EVAL_5125 & _EVAL_2756;
  assign _EVAL_4566 = _EVAL_5068[704];
  assign _EVAL_1359 = _EVAL_1866 ? _EVAL_1074 : _EVAL_6100;
  assign _EVAL_4081 = {1'h0,_EVAL_4828,24'h0};
  assign _EVAL_3351 = _EVAL_2707 ? _EVAL_673 : _EVAL_5013;
  assign _EVAL_2978 = _EVAL_3848 ? {{1'd0}, _EVAL_3532} : _EVAL_990;
  assign _EVAL_766 = {1'h0,_EVAL_546};
  assign _EVAL_3599 = {_EVAL_1907,_EVAL_5670};
  assign _EVAL_3683 = _EVAL_762 & _EVAL_2350;
  assign _EVAL_3883 = {1'h0,_EVAL_4014,_EVAL_4172};
  assign _EVAL_1780 = _EVAL_483 > _EVAL_3937;
  assign _EVAL_4929 = _EVAL_5675 & _EVAL_5396;
  assign _EVAL_2515 = _EVAL_5068[670];
  assign _EVAL_5910 = {{6'd0}, _EVAL_811};
  assign _EVAL_4600 = _EVAL_3772 ? {{1'd0}, _EVAL_3205} : _EVAL_3111;
  assign _EVAL_5597 = _EVAL_6053 & _EVAL_2350;
  assign _EVAL_655 = {{1'd0}, _EVAL_3513};
  assign _EVAL_3444 = {_EVAL_3518,4'hf};
  assign _EVAL_5061 = {1'h0,_EVAL_2341,_EVAL_1048};
  assign _EVAL_192 = _EVAL_3891 ? _EVAL_5551 : _EVAL_4474;
  assign _EVAL_4401 = _EVAL_2101 ? _EVAL_673 : _EVAL_3378;
  assign _EVAL_4770 = {_EVAL_2249,_EVAL_780};
  assign _EVAL_2848 = _EVAL_3786 ? _EVAL_4636 : _EVAL_5441;
  assign _EVAL_3765 = _EVAL_720 > _EVAL_2869;
  assign _EVAL_2026 = _EVAL_559 ? _EVAL_2056 : _EVAL_1646;
  assign _EVAL_4677 = 2'h2 | _EVAL_1141;
  assign _EVAL_1864 = _EVAL_1211 & _EVAL_603;
  assign _EVAL_3798 = _EVAL_1520 > _EVAL_3126;
  assign _EVAL_4735 = _EVAL_4840 | _EVAL_2929;
  assign _EVAL_5674 = _EVAL_901 > _EVAL_1534;
  assign _EVAL_4115 = _EVAL_6073 & _EVAL_3487;
  assign _EVAL_2046 = 10'h281 == _EVAL_5757;
  assign _EVAL_4799 = _EVAL_5762 ? _EVAL_2932 : _EVAL_866;
  assign _EVAL_1473 = {{6'd0}, _EVAL_2776};
  assign _EVAL_2324 = _EVAL_4336 & _EVAL_3234;
  assign _EVAL_5026 = {{6'd0}, _EVAL_2240};
  assign _EVAL_2016 = {{6'd0}, _EVAL_2047};
  assign _EVAL_2578 = _EVAL_4779 & _EVAL_5255;
  assign _EVAL_2058 = _EVAL_3150 & _EVAL_673;
  assign _EVAL_1143 = _EVAL_2091 ? _EVAL_1035 : _EVAL_3289;
  assign _EVAL_5929 = _EVAL_3585 > _EVAL_5058;
  assign _EVAL_5435 = 5'h10 > _EVAL_5297;
  assign _EVAL_2374 = _EVAL_4204 ? _EVAL_673 : _EVAL_1237;
  assign _EVAL_3272 = {1'h0,_EVAL_1593,_EVAL_5237};
  assign _EVAL_3141 = {{6'd0}, _EVAL_5712};
  assign _EVAL_4478 = _EVAL_5951 & _EVAL_2300;
  assign _EVAL_281 = _EVAL_3652 & _EVAL_3607;
  assign _EVAL_2915 = _EVAL_516 & _EVAL_847;
  assign _EVAL_3344 = _EVAL_5579 > _EVAL_4864;
  assign _EVAL_5523 = {{6'd0}, _EVAL_1379};
  assign _EVAL_2749 = {1'h0,_EVAL_2444};
  assign _EVAL_274 = _EVAL_4142 ? {{1'd0}, _EVAL_2786} : _EVAL_5690;
  assign _EVAL_4500 = _EVAL_2096 & _EVAL_2589;
  assign _EVAL_5960 = 10'hff == _EVAL_5757;
  assign _EVAL_1706 = _EVAL_5068[659];
  assign _EVAL_5231 = _EVAL_5145 ? _EVAL_3131 : _EVAL_1576;
  assign _EVAL_3393 = _EVAL_4177 ? _EVAL_3685 : _EVAL_2359;
  assign _EVAL_4676 = _EVAL_1825 & _EVAL_2350;
  assign _EVAL_5279 = {_EVAL_4700,4'hf,_EVAL_3767,4'hf,_EVAL_2546,4'hf,_EVAL_861,4'hf};
  assign _EVAL_2878 = {1'h0,_EVAL_3129,_EVAL_4933};
  assign _EVAL_2994 = {{1'd0}, _EVAL_1271};
  assign _EVAL_1280 = _EVAL_1674[15:4];
  assign _EVAL_4532 = _EVAL_2912 & _EVAL_2756;
  assign _EVAL_5918 = {{1'd0}, _EVAL_4526};
  assign _EVAL_5546 = _EVAL_1860 & _EVAL_3487;
  assign _EVAL_3189 = _EVAL_5751 ? 1'h0 : 1'h1;
  assign _EVAL_5800 = _EVAL_5068[254];
  assign _EVAL_4837 = {1'h0,_EVAL_1408,_EVAL_4056};
  assign _EVAL_5180 = {{1'd0}, _EVAL_5204};
  assign _EVAL_592 = _EVAL_3615 ? {{1'd0}, _EVAL_3686} : _EVAL_1357;
  assign _EVAL_4696 = _EVAL_5064 & _EVAL_417;
  assign _EVAL_1668 = _EVAL_5463 > _EVAL_4953;
  assign _EVAL_5898 = _EVAL_5951 & _EVAL_5169;
  assign _EVAL_4167 = _EVAL_5068[591];
  assign _EVAL_2057 = _EVAL_5064 & _EVAL_2350;
  assign _EVAL_4456 = _EVAL_5951 & _EVAL_923;
  assign _EVAL_4885 = {1'h0,_EVAL_4045,_EVAL_5499};
  assign _EVAL_2751 = {_EVAL_4297,_EVAL_4911};
  assign _EVAL_2568 = _EVAL_763 > _EVAL_3526;
  assign _EVAL_3441 = _EVAL_2058 & _EVAL_2756;
  assign _EVAL_1762 = _EVAL_5068[576];
  assign _EVAL_4708 = {{1'd0}, _EVAL_1092};
  assign _EVAL_4070 = {{1'd0}, _EVAL_3460};
  assign _EVAL_113 = _EVAL_4828;
  assign _EVAL_333 = 10'h202 == _EVAL_5757;
  assign _EVAL_3504 = _EVAL_1775[55:48];
  assign _EVAL_417 = _EVAL_5913 == 4'hf;
  assign _EVAL_498 = {{6'd0}, _EVAL_3883};
  assign _EVAL_847 = _EVAL_1159[24];
  assign _EVAL_2197 = 10'h20a == _EVAL_5757;
  assign _EVAL_1961 = {1'h0,_EVAL_6021,_EVAL_382};
  assign _EVAL_431 = {_EVAL_1551,_EVAL_737};
  assign _EVAL_4441 = _EVAL_5068[585];
  assign _EVAL_1492 = _EVAL_308 ? 1'h0 : 1'h1;
  assign _EVAL_3435 = _EVAL_3215 & _EVAL_417;
  assign _EVAL_3472 = _EVAL_2595 & _EVAL_1937;
  assign _EVAL_1768 = _EVAL_5960 ? _EVAL_1333 : _EVAL_3890;
  assign _EVAL_5197 = {{6'd0}, _EVAL_706};
  assign _EVAL_2586 = {{6'd0}, _EVAL_1239};
  assign _EVAL_4921 = _EVAL_1614 ? _EVAL_498 : _EVAL_416;
  assign _EVAL_3905 = _EVAL_3877 > _EVAL_1914;
  assign _EVAL_2201 = _EVAL_5258 ? _EVAL_673 : _EVAL_5374;
  assign _EVAL_5728 = _EVAL_2743 ? _EVAL_4176 : _EVAL_632;
  assign _EVAL_4840 = _EVAL_3036 | _EVAL_4956;
  assign _EVAL_2180 = _EVAL_5725 > _EVAL_5793;
  assign _EVAL_5952 = _EVAL_1758 ? _EVAL_3119 : _EVAL_2054;
  assign _EVAL_1688 = _EVAL_3772 ? _EVAL_5547 : _EVAL_4182;
  assign _EVAL_3067 = {_EVAL_5860,_EVAL_4908};
  assign _EVAL_543 = _EVAL_5068[642];
  assign _EVAL_3570 = {1'h0,_EVAL_5232};
  assign _EVAL_2852 = 10'h2c0 == _EVAL_5757;
  assign _EVAL_2979 = _EVAL_3128 > _EVAL_3046;
  assign _EVAL_2968 = 10'h282 == _EVAL_5757;
  assign _EVAL_2488 = {{6'd0}, _EVAL_4290};
  assign _EVAL_4637 = 10'h28d == _EVAL_5757;
  assign _EVAL_3410 = _EVAL_2277 & _EVAL_2360;
  assign _EVAL_5884 = 3'h4 | _EVAL_4889;
  assign _EVAL_872 = _EVAL_2112 ? _EVAL_220 : _EVAL_2385;
  assign _EVAL_2528 = _EVAL_5125 & _EVAL_417;
  assign _EVAL_1713 = _EVAL_5951 & _EVAL_2074;
  assign _EVAL_5171 = 4'h8 | _EVAL_5626;
  assign _EVAL_5058 = _EVAL_468 ? _EVAL_5794 : _EVAL_4178;
  assign _EVAL_1398 = {{6'd0}, _EVAL_337};
  assign _EVAL_2300 = _EVAL_5068[646];
  assign _EVAL_2487 = {{6'd0}, _EVAL_1056};
  assign _EVAL_6023 = _EVAL_5096 & _EVAL_4477;
  assign _EVAL_5375 = _EVAL_5505 ? 1'h0 : 1'h1;
  assign _EVAL_6049 = _EVAL_1613 & _EVAL_673;
  assign _EVAL_3834 = {_EVAL_2081,_EVAL_1356};
  assign _EVAL_3697 = {1'h0,_EVAL_2876,_EVAL_5156};
  assign _EVAL_4260 = _EVAL_2707 ? _EVAL_981 : _EVAL_1821;
  assign _EVAL_2706 = _EVAL_5068[256];
  assign _EVAL_1190 = {{6'd0}, _EVAL_3012};
  assign _EVAL_3145 = _EVAL_796 & _EVAL_847;
  assign _EVAL_5086 = _EVAL_2474 & _EVAL_1937;
  assign _EVAL_4170 = _EVAL_5929 ? {{1'd0}, _EVAL_1908} : _EVAL_1874;
  assign _EVAL_419 = {1'h0,_EVAL_2589};
  assign _EVAL_5915 = {{6'd0}, _EVAL_648};
  assign _EVAL_5441 = _EVAL_2855 ? _EVAL_733 : _EVAL_647;
  assign _EVAL_3975 = {1'h0,_EVAL_1388};
  assign _EVAL_3806 = {1'h0,_EVAL_4103,_EVAL_5318};
  assign _EVAL_5828 = {{6'd0}, _EVAL_2113};
  assign _EVAL_4614 = _EVAL_4603 > _EVAL_3380;
  assign _EVAL_2099 = _EVAL_4159 ? _EVAL_2840 : _EVAL_2026;
  assign _EVAL_5965 = _EVAL_3039 ? _EVAL_673 : _EVAL_5628;
  assign _EVAL_3750 = _EVAL_640 ? _EVAL_5185 : _EVAL_238;
  assign _EVAL_2495 = _EVAL_2486 & _EVAL_1937;
  assign _EVAL_1464 = _EVAL_5068[606];
  assign _EVAL_3164 = _EVAL_2428 ? _EVAL_673 : _EVAL_2048;
  assign _EVAL_1020 = _EVAL_772 > _EVAL_1950;
  assign _EVAL_2641 = {{6'd0}, _EVAL_4173};
  assign _EVAL_2225 = _EVAL_4370 | _EVAL_5557;
  assign _EVAL_5225 = _EVAL_5369 & _EVAL_546;
  assign _EVAL_511 = _EVAL_4980 & _EVAL_673;
  assign _EVAL_1026 = {{6'd0}, _EVAL_5522};
  assign _EVAL_5220 = _EVAL_1737 ? _EVAL_5899 : _EVAL_858;
  assign _EVAL_962 = {1'h0,_EVAL_5890,_EVAL_4826};
  assign _EVAL_5410 = {1'h0,_EVAL_381,_EVAL_2970};
  assign _EVAL_4515 = {{2'd0}, _EVAL_5876};
  assign _EVAL_3356 = {{6'd0}, _EVAL_3259};
  assign _EVAL_864 = _EVAL_1761 & _EVAL_847;
  assign _EVAL_3423 = _EVAL_2218 + 64'h1;
  assign _EVAL_5859 = {1'h0,_EVAL_3001};
  assign _EVAL_5556 = _EVAL_5068[596];
  assign _EVAL_3921 = 10'h299 == _EVAL_5757;
  assign _EVAL_5638 = {1'h0,_EVAL_3962};
  assign _EVAL_2132 = {1'h0,_EVAL_3639,_EVAL_3832};
  assign _EVAL_3105 = _EVAL_1217 ? _EVAL_673 : _EVAL_6000;
  assign _EVAL_5872 = _EVAL_3419 ? _EVAL_673 : _EVAL_2880;
  assign _EVAL_1461 = {{6'd0}, _EVAL_2132};
  assign _EVAL_291 = {{6'd0}, _EVAL_5669};
  assign _EVAL_1164 = _EVAL_1228 ? {{1'd0}, _EVAL_5494} : 2'h2;
  assign _EVAL_1451 = _EVAL_5064 & _EVAL_2756;
  assign _EVAL_6078 = _EVAL_1815 ? 1'h0 : 1'h1;
  assign _EVAL_173 = {{6'd0}, _EVAL_264};
  assign _EVAL_300 = _EVAL_5113 & _EVAL_2756;
  assign _EVAL_5891 = {{6'd0}, _EVAL_6034};
  assign _EVAL_1712 = {_EVAL_3310,4'hf,_EVAL_1318,4'hf,_EVAL_1427,4'hf,_EVAL_3429,4'hf};
  assign _EVAL_2668 = _EVAL_783 & _EVAL_5600;
  assign _EVAL_2152 = {{6'd0}, _EVAL_1177};
  assign _EVAL_1163 = _EVAL_1240 & _EVAL_1187;
  assign _EVAL_5757 = {_EVAL_5475,_EVAL_1705,_EVAL_5520,_EVAL_1236,_EVAL_2111,_EVAL_1681,_EVAL_4377,_EVAL_4198,_EVAL_3810,_EVAL_5931};
  assign _EVAL_1885 = _EVAL_5045 ? 1'h0 : 1'h1;
  assign _EVAL_5029 = _EVAL_1436 & _EVAL_847;
  assign _EVAL_4632 = _EVAL_1815 ? _EVAL_4266 : _EVAL_863;
  assign _EVAL_4839 = _EVAL_6052 & _EVAL_847;
  assign _EVAL_5636 = 10'h24d == _EVAL_5757;
  assign _EVAL_5112 = _EVAL_3870[3:0];
  assign _EVAL_5034 = _EVAL_2784 & _EVAL_417;
  assign _EVAL_1970 = 2'h2 | _EVAL_2959;
  assign _EVAL_4562 = 10'h28a == _EVAL_5757;
  assign _EVAL_1135 = _EVAL_1414 > _EVAL_853;
  assign _EVAL_4025 = _EVAL_606 & _EVAL_3487;
  assign _EVAL_452 = {1'h0,_EVAL_3294};
  assign _EVAL_3906 = {_EVAL_4005,_EVAL_2183};
  assign _EVAL_5448 = _EVAL_1751 & _EVAL_2350;
  assign _EVAL_5792 = 10'h285 == _EVAL_5757;
  assign _EVAL_5984 = _EVAL_5068[665];
  assign _EVAL_1204 = {{6'd0}, _EVAL_4977};
  assign _EVAL_3229 = {{6'd0}, _EVAL_5875};
  assign _EVAL_1054 = 10'h101 == _EVAL_5757;
  assign _EVAL_4747 = _EVAL_1780 ? 1'h0 : 1'h1;
  assign _EVAL_2003 = {_EVAL_1163,_EVAL_4416};
  assign _EVAL_1983 = {_EVAL_2324,_EVAL_1863};
  assign _EVAL_1295 = {{6'd0}, _EVAL_3779};
  assign _EVAL_1098 = _EVAL_4124 ? 1'h0 : 1'h1;
  assign _EVAL_5645 = {{1'd0}, _EVAL_1805};
  assign _EVAL_5247 = {_EVAL_199,_EVAL_1143,_EVAL_4995,_EVAL_1238,_EVAL_5612,_EVAL_4705,_EVAL_5287,_EVAL_1813};
  assign _EVAL_4275 = {1'h0,_EVAL_2828,_EVAL_2016};
  assign _EVAL_170 = 2'h2 | _EVAL_728;
  assign _EVAL_2948 = {{1'd0}, _EVAL_3819};
  assign _EVAL_1796 = _EVAL_4204 ? _EVAL_3297 : _EVAL_784;
  assign _EVAL_1859 = {{6'd0}, _EVAL_4417};
  assign _EVAL_6082 = _EVAL_2042 ? _EVAL_5742 : _EVAL_707;
  assign _EVAL_6053 = _EVAL_1138 & _EVAL_673;
  assign _EVAL_5165 = {_EVAL_1864,_EVAL_2030};
  assign _EVAL_4728 = _EVAL_192 > _EVAL_2522;
  assign _EVAL_753 = {{6'd0}, _EVAL_5244};
  assign _EVAL_741 = {{6'd0}, _EVAL_4846};
  assign _EVAL_3125 = 3'h4 | _EVAL_2639;
  assign _EVAL_4303 = _EVAL_4895 ? _EVAL_673 : _EVAL_5595;
  assign _EVAL_2954 = _EVAL_3934 & _EVAL_673;
  assign _EVAL_2611 = _EVAL_1378 & _EVAL_2350;
  assign _EVAL_2697 = {{6'd0}, _EVAL_4969};
  assign _EVAL_1738 = {_EVAL_2668,_EVAL_558};
  assign _EVAL_3126 = _EVAL_2128 ? _EVAL_6063 : _EVAL_3963;
  assign _EVAL_3615 = _EVAL_687 > _EVAL_4632;
  assign _EVAL_5699 = _EVAL_4010 & _EVAL_847;
  assign _EVAL_3944 = _EVAL_5068[581];
  assign _EVAL_4041 = {1'h0,_EVAL_943,_EVAL_4313};
  assign _EVAL_5325 = {_EVAL_4480,_EVAL_1891};
  assign _EVAL_167 = {{1'd0}, _EVAL_517};
  assign _EVAL_4215 = _EVAL_5951 & _EVAL_3944;
  assign _EVAL_3903 = {_EVAL_824,_EVAL_861};
  assign _EVAL_1438 = _EVAL_5951 & _EVAL_2052;
  assign _EVAL_3627 = _EVAL_5617 ? 1'h0 : 1'h1;
  assign _EVAL_1030 = 10'h290 == _EVAL_5757;
  assign _EVAL_329 = _EVAL_4415 ? _EVAL_1339 : _EVAL_3599;
  assign _EVAL_2894 = {1'h0,_EVAL_4065,_EVAL_575};
  assign _EVAL_3814 = _EVAL_5716 & _EVAL_673;
  assign _EVAL_1982 = _EVAL_5836 & _EVAL_2756;
  assign _EVAL_1892 = {{6'd0}, _EVAL_5333};
  assign _EVAL_5248 = {_EVAL_3693,4'hf,_EVAL_2183,4'hf,_EVAL_1720,4'hf,_EVAL_6040,4'hf};
  assign _EVAL_3080 = _EVAL_4410 ? _EVAL_673 : _EVAL_3164;
  assign _EVAL_1377 = _EVAL_5951 & _EVAL_1087;
  assign _EVAL_455 = _EVAL_2486 & _EVAL_2756;
  assign _EVAL_4883 = {_EVAL_2013,_EVAL_4574};
  assign _EVAL_471 = _EVAL_1761 & _EVAL_3154;
  assign _EVAL_1904 = {_EVAL_1524,_EVAL_4631};
  assign _EVAL_907 = _EVAL_5951 & _EVAL_550;
  assign _EVAL_4776 = _EVAL_942 ? _EVAL_4633 : _EVAL_2610;
  assign _EVAL_2543 = {_EVAL_412,28'hf000000};
  assign _EVAL_3465 = _EVAL_2587 ? _EVAL_743 : _EVAL_445;
  assign _EVAL_3918 = {{6'd0}, _EVAL_4221};
  assign _EVAL_4824 = {4'h0,_EVAL_344};
  assign _EVAL_2959 = {{1'd0}, _EVAL_4548};
  assign _EVAL_1758 = _EVAL_3119 > _EVAL_2054;
  assign _EVAL_2085 = {_EVAL_4631,4'hf,_EVAL_5727,4'hf,_EVAL_4786,4'hf};
  assign _EVAL_5860 = _EVAL_2148 & _EVAL_4810;
  assign _EVAL_4400 = {1'h0,_EVAL_2766,_EVAL_5926};
  assign _EVAL_5584 = _EVAL_5806 ? _EVAL_2178 : _EVAL_4665;
  assign _EVAL_1080 = _EVAL_2980 ? 8'hff : 8'h0;
  assign _EVAL_176 = _EVAL_218 & _EVAL_3487;
  assign _EVAL_2263 = {_EVAL_164,4'hf,_EVAL_4181,4'hf,_EVAL_3173,4'hf,_EVAL_2889,4'hf};
  assign _EVAL_5244 = {1'h0,_EVAL_2177};
  assign _EVAL_2102 = {1'h0,_EVAL_2616,_EVAL_1927};
  assign _EVAL_6014 = _EVAL_1311 & _EVAL_487;
  assign _EVAL_1573 = {{6'd0}, _EVAL_924};
  assign _EVAL_3762 = _EVAL_1032 ? 1'h0 : 1'h1;
  assign _EVAL_6006 = _EVAL_5089 ? _EVAL_3797 : _EVAL_3332;
  assign _EVAL_4640 = {{6'd0}, _EVAL_419};
  assign _EVAL_288 = {{6'd0}, _EVAL_1552};
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_164 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_212 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_236 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_272 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_277 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_296 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_355 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_356 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_381 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_404 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_412 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_454 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_484 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_487 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_493 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_506 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_507 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_531 = _RAND_17[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_542 = _RAND_18[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_546 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_558 = _RAND_20[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_560 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_561 = _RAND_22[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_563 = _RAND_23[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_582 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_603 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_607 = _RAND_26[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_616 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_643 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_644 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_653 = _RAND_30[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_661 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_666 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_690 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_702 = _RAND_34[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_703 = _RAND_35[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_727 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_737 = _RAND_37[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _EVAL_780 = _RAND_38[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _EVAL_783 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _EVAL_834 = _RAND_40[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _EVAL_861 = _RAND_41[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _EVAL_880 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _EVAL_887 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _EVAL_891 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _EVAL_896 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _EVAL_899 = _RAND_46[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _EVAL_906 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _EVAL_943 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _EVAL_994 = _RAND_49[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _EVAL_1028 = _RAND_50[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _EVAL_1040 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _EVAL_1041 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _EVAL_1052 = _RAND_53[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _EVAL_1057 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _EVAL_1121 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _EVAL_1131 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _EVAL_1147 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _EVAL_1166 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _EVAL_1186 = _RAND_59[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _EVAL_1187 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _EVAL_1188 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _EVAL_1206 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _EVAL_1211 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _EVAL_1229 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _EVAL_1235 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _EVAL_1240 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _EVAL_1245 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _EVAL_1273 = _RAND_68[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _EVAL_1286 = _RAND_69[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _EVAL_1287 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _EVAL_1288 = _RAND_71[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _EVAL_1289 = _RAND_72[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _EVAL_1293 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _EVAL_1301 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _EVAL_1311 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _EVAL_1314 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _EVAL_1318 = _RAND_77[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _EVAL_1331 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _EVAL_1342 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _EVAL_1351 = _RAND_80[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _EVAL_1356 = _RAND_81[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _EVAL_1383 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _EVAL_1388 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _EVAL_1396 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _EVAL_1407 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _EVAL_1408 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _EVAL_1427 = _RAND_87[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _EVAL_1440 = _RAND_88[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _EVAL_1442 = _RAND_89[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _EVAL_1484 = _RAND_90[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _EVAL_1493 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _EVAL_1506 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _EVAL_1510 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _EVAL_1515 = _RAND_94[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _EVAL_1544 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _EVAL_1581 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _EVAL_1593 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _EVAL_1602 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _EVAL_1610 = _RAND_99[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _EVAL_1618 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _EVAL_1629 = _RAND_101[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _EVAL_1641 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _EVAL_1645 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _EVAL_1664 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _EVAL_1670 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _EVAL_1671 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _EVAL_1672 = _RAND_107[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _EVAL_1676 = _RAND_108[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _EVAL_1686 = _RAND_109[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _EVAL_1720 = _RAND_110[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _EVAL_1730 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _EVAL_1746 = _RAND_112[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _EVAL_1765 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {2{`RANDOM}};
  _EVAL_1775 = _RAND_114[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _EVAL_1777 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _EVAL_1797 = _RAND_116[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _EVAL_1820 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _EVAL_1822 = _RAND_118[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _EVAL_1826 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _EVAL_1828 = _RAND_120[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _EVAL_1831 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _EVAL_1863 = _RAND_122[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _EVAL_1875 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _EVAL_1880 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _EVAL_1882 = _RAND_125[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _EVAL_1891 = _RAND_126[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _EVAL_1917 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _EVAL_1929 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _EVAL_1942 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _EVAL_2009 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _EVAL_2030 = _RAND_131[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _EVAL_2065 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _EVAL_2086 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _EVAL_2096 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _EVAL_2148 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _EVAL_2154 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _EVAL_2162 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _EVAL_2177 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _EVAL_2183 = _RAND_139[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _EVAL_2203 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _EVAL_2215 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {2{`RANDOM}};
  _EVAL_2218 = _RAND_142[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _EVAL_2229 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _EVAL_2233 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _EVAL_2247 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _EVAL_2277 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _EVAL_2291 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _EVAL_2293 = _RAND_148[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _EVAL_2301 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _EVAL_2307 = _RAND_150[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _EVAL_2308 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _EVAL_2312 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _EVAL_2339 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _EVAL_2341 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _EVAL_2357 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _EVAL_2360 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _EVAL_2366 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _EVAL_2381 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _EVAL_2393 = _RAND_159[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _EVAL_2422 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _EVAL_2444 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _EVAL_2462 = _RAND_162[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _EVAL_2484 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _EVAL_2490 = _RAND_164[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _EVAL_2493 = _RAND_165[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _EVAL_2516 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _EVAL_2537 = _RAND_167[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _EVAL_2546 = _RAND_168[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _EVAL_2557 = _RAND_169[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _EVAL_2561 = _RAND_170[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _EVAL_2580 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _EVAL_2583 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _EVAL_2589 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _EVAL_2616 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _EVAL_2626 = _RAND_175[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _EVAL_2629 = _RAND_176[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _EVAL_2667 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _EVAL_2669 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _EVAL_2690 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _EVAL_2717 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _EVAL_2766 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _EVAL_2778 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _EVAL_2781 = _RAND_183[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _EVAL_2782 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _EVAL_2806 = _RAND_185[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _EVAL_2825 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _EVAL_2827 = _RAND_187[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _EVAL_2828 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _EVAL_2837 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _EVAL_2847 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _EVAL_2876 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _EVAL_2889 = _RAND_192[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _EVAL_2905 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _EVAL_2910 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _EVAL_2918 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _EVAL_2920 = _RAND_196[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _EVAL_2984 = _RAND_197[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _EVAL_2988 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _EVAL_2993 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _EVAL_3001 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _EVAL_3005 = _RAND_201[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _EVAL_3040 = _RAND_202[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _EVAL_3062 = _RAND_203[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _EVAL_3108 = _RAND_204[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _EVAL_3129 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _EVAL_3133 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _EVAL_3152 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _EVAL_3171 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _EVAL_3172 = _RAND_209[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _EVAL_3173 = _RAND_210[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _EVAL_3181 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _EVAL_3194 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _EVAL_3196 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _EVAL_3197 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _EVAL_3203 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _EVAL_3213 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _EVAL_3225 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _EVAL_3234 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _EVAL_3256 = _RAND_219[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _EVAL_3280 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _EVAL_3286 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _EVAL_3294 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _EVAL_3310 = _RAND_223[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _EVAL_3327 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _EVAL_3363 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _EVAL_3374 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _EVAL_3384 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _EVAL_3404 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _EVAL_3429 = _RAND_229[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _EVAL_3449 = _RAND_230[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _EVAL_3450 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _EVAL_3456 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _EVAL_3464 = _RAND_233[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _EVAL_3467 = _RAND_234[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _EVAL_3538 = _RAND_235[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _EVAL_3580 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _EVAL_3584 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _EVAL_3589 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _EVAL_3594 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _EVAL_3607 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _EVAL_3609 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _EVAL_3629 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _EVAL_3634 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _EVAL_3639 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _EVAL_3652 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _EVAL_3673 = _RAND_246[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _EVAL_3676 = _RAND_247[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _EVAL_3692 = _RAND_248[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _EVAL_3693 = _RAND_249[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _EVAL_3722 = _RAND_250[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _EVAL_3743 = _RAND_251[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _EVAL_3767 = _RAND_252[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _EVAL_3771 = _RAND_253[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _EVAL_3783 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _EVAL_3789 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _EVAL_3843 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _EVAL_3847 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _EVAL_3857 = _RAND_258[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _EVAL_3866 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _EVAL_3887 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _EVAL_3914 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _EVAL_3940 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _EVAL_3945 = _RAND_263[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _EVAL_3946 = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _EVAL_3962 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _EVAL_3965 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _EVAL_3983 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _EVAL_3986 = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _EVAL_4007 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _EVAL_4014 = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _EVAL_4019 = _RAND_271[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _EVAL_4040 = _RAND_272[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _EVAL_4045 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _EVAL_4051 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _EVAL_4053 = _RAND_275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _EVAL_4065 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _EVAL_4080 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _EVAL_4085 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _EVAL_4087 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _EVAL_4103 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _EVAL_4119 = _RAND_281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _EVAL_4181 = _RAND_282[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _EVAL_4184 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _EVAL_4233 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _EVAL_4264 = _RAND_285[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _EVAL_4291 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _EVAL_4304 = _RAND_287[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _EVAL_4308 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _EVAL_4336 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _EVAL_4338 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _EVAL_4348 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _EVAL_4367 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _EVAL_4374 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _EVAL_4390 = _RAND_294[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _EVAL_4397 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _EVAL_4398 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _EVAL_4404 = _RAND_297[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _EVAL_4416 = _RAND_298[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _EVAL_4443 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _EVAL_4479 = _RAND_300[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _EVAL_4518 = _RAND_301[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _EVAL_4571 = _RAND_302[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _EVAL_4572 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _EVAL_4574 = _RAND_304[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _EVAL_4584 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _EVAL_4588 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _EVAL_4612 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _EVAL_4620 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _EVAL_4624 = _RAND_309[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _EVAL_4631 = _RAND_310[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _EVAL_4700 = _RAND_311[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _EVAL_4711 = _RAND_312[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _EVAL_4732 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _EVAL_4738 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _EVAL_4742 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _EVAL_4779 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _EVAL_4785 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _EVAL_4786 = _RAND_318[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _EVAL_4807 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _EVAL_4808 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _EVAL_4810 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _EVAL_4828 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _EVAL_4843 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _EVAL_4908 = _RAND_324[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _EVAL_4911 = _RAND_325[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _EVAL_4922 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _EVAL_4927 = _RAND_327[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _EVAL_4932 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _EVAL_4944 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _EVAL_4955 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _EVAL_4965 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _EVAL_4997 = _RAND_332[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _EVAL_5002 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _EVAL_5008 = _RAND_334[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _EVAL_5009 = _RAND_335[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _EVAL_5039 = _RAND_336[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _EVAL_5080 = _RAND_337[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _EVAL_5101 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _EVAL_5104 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _EVAL_5139 = _RAND_340[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _EVAL_5142 = _RAND_341[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _EVAL_5147 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _EVAL_5163 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _EVAL_5190 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _EVAL_5232 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _EVAL_5249 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _EVAL_5255 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _EVAL_5293 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _EVAL_5300 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _EVAL_5307 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _EVAL_5309 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _EVAL_5311 = _RAND_352[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _EVAL_5315 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _EVAL_5345 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _EVAL_5369 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _EVAL_5386 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _EVAL_5389 = _RAND_357[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _EVAL_5396 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _EVAL_5409 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _EVAL_5411 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _EVAL_5479 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _EVAL_5484 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _EVAL_5518 = _RAND_363[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _EVAL_5521 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _EVAL_5535 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _EVAL_5537 = _RAND_366[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _EVAL_5558 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _EVAL_5600 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _EVAL_5606 = _RAND_369[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _EVAL_5608 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _EVAL_5609 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _EVAL_5623 = _RAND_372[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _EVAL_5624 = _RAND_373[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _EVAL_5629 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _EVAL_5635 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _EVAL_5665 = _RAND_376[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _EVAL_5667 = _RAND_377[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _EVAL_5670 = _RAND_378[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _EVAL_5675 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _EVAL_5684 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _EVAL_5696 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _EVAL_5697 = _RAND_382[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _EVAL_5713 = _RAND_383[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _EVAL_5727 = _RAND_384[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _EVAL_5735 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _EVAL_5741 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _EVAL_5743 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _EVAL_5765 = _RAND_388[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _EVAL_5781 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _EVAL_5846 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _EVAL_5878 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _EVAL_5890 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _EVAL_5916 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _EVAL_5924 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _EVAL_5940 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _EVAL_5962 = _RAND_396[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _EVAL_5981 = _RAND_397[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _EVAL_5985 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _EVAL_6021 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _EVAL_6030 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _EVAL_6040 = _RAND_401[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _EVAL_6098 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_106) begin
    if (_EVAL_306) begin
      _EVAL_164 <= _EVAL_3709;
    end
    _EVAL_212 <= _EVAL_9;
    if (_EVAL_5603) begin
      _EVAL_236 <= _EVAL_1374;
    end
    if (_EVAL_465) begin
      _EVAL_272 <= _EVAL_2231;
    end
    _EVAL_277 <= _EVAL_128;
    if (_EVAL_3861) begin
      _EVAL_296 <= _EVAL_4709;
    end
    if (_EVAL_4242) begin
      _EVAL_355 <= _EVAL_338;
    end
    _EVAL_356 <= _EVAL_75;
    _EVAL_381 <= _EVAL_66;
    if (_EVAL_4030) begin
      _EVAL_404 <= 8'h0;
    end else begin
      _EVAL_404 <= _EVAL_1976;
    end
    if (_EVAL_5188) begin
      _EVAL_412 <= _EVAL_3709;
    end
    if (_EVAL_4414) begin
      _EVAL_454 <= _EVAL_1967;
    end
    if (_EVAL_24) begin
      _EVAL_484 <= 1'h0;
    end else if (_EVAL_4025) begin
      _EVAL_484 <= _EVAL_338;
    end
    if (_EVAL_553) begin
      _EVAL_487 <= _EVAL_3222;
    end
    if (_EVAL_4406) begin
      _EVAL_493 <= _EVAL_4088;
    end
    if (_EVAL_2922) begin
      _EVAL_506 <= _EVAL_3222;
    end
    if (_EVAL_3336) begin
      _EVAL_507 <= _EVAL_1967;
    end
    if (_EVAL_3501) begin
      _EVAL_531 <= _EVAL_4088;
    end
    if (_EVAL_3646) begin
      _EVAL_542 <= _EVAL_3709;
    end
    if (_EVAL_4096) begin
      _EVAL_546 <= _EVAL_338;
    end
    if (_EVAL_5730) begin
      _EVAL_558 <= _EVAL_2231;
    end
    if (_EVAL_5745) begin
      _EVAL_560 <= _EVAL_1374;
    end
    if (_EVAL_3266) begin
      _EVAL_561 <= _EVAL_4709;
    end
    if (_EVAL_3158) begin
      _EVAL_563 <= _EVAL_2231;
    end
    if (_EVAL_1666) begin
      _EVAL_582 <= _EVAL_1374;
    end
    if (_EVAL_3493) begin
      _EVAL_603 <= _EVAL_3222;
    end
    if (_EVAL_2239) begin
      _EVAL_607 <= _EVAL_2231;
    end
    _EVAL_616 <= _EVAL_127;
    if (_EVAL_3854) begin
      _EVAL_643 <= _EVAL_338;
    end
    _EVAL_644 <= _EVAL_95;
    if (_EVAL_2417) begin
      _EVAL_653 <= _EVAL_2231;
    end
    if (_EVAL_3939) begin
      _EVAL_661 <= _EVAL_1967;
    end
    if (_EVAL_2198) begin
      _EVAL_666 <= _EVAL_1374;
    end
    _EVAL_690 <= _EVAL_43;
    if (_EVAL_5131) begin
      _EVAL_702 <= _EVAL_4088;
    end
    if (_EVAL_2577) begin
      _EVAL_703 <= _EVAL_2231;
    end
    _EVAL_727 <= _EVAL_31;
    if (_EVAL_2598) begin
      _EVAL_737 <= _EVAL_3709;
    end
    if (_EVAL_300) begin
      _EVAL_780 <= _EVAL_3709;
    end
    _EVAL_783 <= _EVAL_57;
    if (_EVAL_1367) begin
      _EVAL_834 <= _EVAL_2231;
    end
    if (_EVAL_1250) begin
      _EVAL_861 <= _EVAL_2231;
    end
    _EVAL_880 <= _EVAL_82;
    if (_EVAL_5759) begin
      _EVAL_887 <= _EVAL_1967;
    end
    _EVAL_891 <= _EVAL_134;
    if (_EVAL_2168) begin
      _EVAL_896 <= _EVAL_3222;
    end
    if (_EVAL_3441) begin
      _EVAL_899 <= _EVAL_3709;
    end
    if (_EVAL_6023) begin
      _EVAL_906 <= _EVAL_3222;
    end
    _EVAL_943 <= _EVAL_85;
    if (_EVAL_4753) begin
      _EVAL_994 <= _EVAL_4709;
    end
    if (_EVAL_601) begin
      _EVAL_1028 <= _EVAL_3709;
    end
    _EVAL_1040 <= _EVAL_40;
    if (_EVAL_3758) begin
      _EVAL_1041 <= _EVAL_1374;
    end
    if (_EVAL_1871) begin
      _EVAL_1052 <= _EVAL_2231;
    end
    _EVAL_1057 <= _EVAL_121;
    _EVAL_1121 <= _EVAL_50;
    if (_EVAL_4819) begin
      _EVAL_1131 <= _EVAL_3222;
    end
    _EVAL_1147 <= _EVAL_115;
    if (_EVAL_1261) begin
      _EVAL_1166 <= _EVAL_1967;
    end
    if (_EVAL_3422) begin
      _EVAL_1186 <= _EVAL_2231;
    end
    if (_EVAL_759) begin
      _EVAL_1187 <= _EVAL_338;
    end
    if (_EVAL_2108) begin
      _EVAL_1188 <= _EVAL_1374;
    end
    _EVAL_1206 <= _EVAL_42;
    _EVAL_1211 <= _EVAL_136;
    _EVAL_1229 <= _EVAL_20;
    _EVAL_1235 <= _EVAL_17;
    _EVAL_1240 <= _EVAL_1;
    if (_EVAL_4839) begin
      _EVAL_1245 <= _EVAL_1374;
    end
    if (_EVAL_3435) begin
      _EVAL_1273 <= _EVAL_4088;
    end
    if (_EVAL_5049) begin
      _EVAL_1286 <= {{1'd0}, _EVAL_4990};
    end else begin
      _EVAL_1286 <= _EVAL_4685;
    end
    if (_EVAL_3087) begin
      _EVAL_1287 <= _EVAL_1967;
    end
    if (_EVAL_1150) begin
      _EVAL_1288 <= _EVAL_4709;
    end
    if (_EVAL_5909) begin
      _EVAL_1289 <= _EVAL_3709;
    end
    if (_EVAL_397) begin
      _EVAL_1293 <= _EVAL_1374;
    end
    if (_EVAL_5012) begin
      _EVAL_1301 <= _EVAL_3222;
    end
    _EVAL_1311 <= _EVAL_74;
    _EVAL_1314 <= _EVAL_64;
    if (_EVAL_2022) begin
      _EVAL_1318 <= _EVAL_4709;
    end
    if (_EVAL_1844) begin
      _EVAL_1331 <= _EVAL_1374;
    end
    if (_EVAL_3285) begin
      _EVAL_1342 <= _EVAL_3222;
    end
    if (_EVAL_2523) begin
      _EVAL_1351 <= _EVAL_3709;
    end
    if (_EVAL_2495) begin
      _EVAL_1356 <= _EVAL_2231;
    end
    if (_EVAL_765) begin
      _EVAL_1383 <= _EVAL_1374;
    end
    if (_EVAL_5627) begin
      _EVAL_1388 <= _EVAL_338;
    end
    _EVAL_1396 <= _EVAL_141;
    if (_EVAL_2244) begin
      _EVAL_1407 <= _EVAL_1374;
    end
    _EVAL_1408 <= _EVAL_30;
    if (_EVAL_5907) begin
      _EVAL_1427 <= _EVAL_4088;
    end
    if (_EVAL_844) begin
      _EVAL_1440 <= _EVAL_4088;
    end
    if (_EVAL_5086) begin
      _EVAL_1442 <= _EVAL_2231;
    end
    if (_EVAL_4008) begin
      _EVAL_1484 <= _EVAL_3709;
    end
    _EVAL_1493 <= _EVAL_144;
    if (_EVAL_471) begin
      _EVAL_1506 <= _EVAL_1967;
    end
    if (_EVAL_5421) begin
      _EVAL_1510 <= _EVAL_1374;
    end
    if (_EVAL_2202) begin
      _EVAL_1515 <= _EVAL_3709;
    end
    if (_EVAL_948) begin
      _EVAL_1544 <= _EVAL_338;
    end
    _EVAL_1581 <= _EVAL_2218 >= _EVAL_1775;
    _EVAL_1593 <= _EVAL_147;
    if (_EVAL_4437) begin
      _EVAL_1602 <= _EVAL_3222;
    end
    if (_EVAL_3051) begin
      _EVAL_1610 <= _EVAL_4709;
    end
    if (_EVAL_5150) begin
      _EVAL_1618 <= _EVAL_3222;
    end
    if (_EVAL_4339) begin
      _EVAL_1629 <= _EVAL_4709;
    end
    if (_EVAL_5294) begin
      _EVAL_1641 <= _EVAL_338;
    end
    if (_EVAL_978) begin
      _EVAL_1645 <= _EVAL_1374;
    end
    _EVAL_1664 <= _EVAL_98;
    if (_EVAL_2758) begin
      _EVAL_1670 <= _EVAL_1967;
    end
    if (_EVAL_158) begin
      _EVAL_1671 <= _EVAL_1374;
    end
    if (_EVAL_3799) begin
      _EVAL_1672 <= _EVAL_2231;
    end
    if (_EVAL_3472) begin
      _EVAL_1676 <= _EVAL_2231;
    end
    _EVAL_1686 <= _EVAL_3444[7:0];
    if (_EVAL_2528) begin
      _EVAL_1720 <= _EVAL_4088;
    end
    _EVAL_1730 <= _EVAL_116;
    if (_EVAL_24) begin
      _EVAL_1746 <= 4'h0;
    end else begin
      _EVAL_1746 <= _EVAL_3945;
    end
    _EVAL_1765 <= _EVAL_56;
    if (_EVAL_4721) begin
      _EVAL_1775 <= _EVAL_4725;
    end
    if (_EVAL_197) begin
      _EVAL_1777 <= _EVAL_1967;
    end
    if (_EVAL_2119) begin
      _EVAL_1797 <= _EVAL_4088;
    end
    if (_EVAL_5326) begin
      _EVAL_1820 <= _EVAL_1967;
    end
    if (_EVAL_5597) begin
      _EVAL_1822 <= _EVAL_4709;
    end
    if (_EVAL_5646) begin
      _EVAL_1826 <= _EVAL_1374;
    end
    if (_EVAL_1454) begin
      _EVAL_1828 <= _EVAL_4088;
    end
    if (_EVAL_1565) begin
      _EVAL_1831 <= _EVAL_1967;
    end
    if (_EVAL_6092) begin
      _EVAL_1863 <= _EVAL_3709;
    end
    _EVAL_1875 <= _EVAL_132;
    if (_EVAL_5771) begin
      _EVAL_1880 <= _EVAL_1967;
    end
    if (_EVAL_3795) begin
      _EVAL_1882 <= _EVAL_4088;
    end
    if (_EVAL_1005) begin
      _EVAL_1891 <= _EVAL_4088;
    end
    _EVAL_1917 <= _EVAL_90;
    if (_EVAL_489) begin
      _EVAL_1929 <= _EVAL_3222;
    end
    if (_EVAL_5619) begin
      _EVAL_1942 <= _EVAL_338;
    end
    _EVAL_2009 <= _EVAL_36;
    if (_EVAL_934) begin
      _EVAL_2030 <= _EVAL_4709;
    end
    _EVAL_2065 <= _EVAL_16;
    _EVAL_2086 <= _EVAL_54;
    _EVAL_2096 <= _EVAL_13;
    _EVAL_2148 <= _EVAL_45;
    _EVAL_2154 <= _EVAL_93;
    if (_EVAL_2400) begin
      _EVAL_2162 <= _EVAL_1374;
    end
    _EVAL_2177 <= _EVAL_51;
    if (_EVAL_3311) begin
      _EVAL_2183 <= _EVAL_4709;
    end
    if (_EVAL_1592) begin
      _EVAL_2203 <= _EVAL_3222;
    end
    _EVAL_2215 <= _EVAL_0;
    if (_EVAL_24) begin
      _EVAL_2218 <= 64'h0;
    end else if (_EVAL_5903) begin
      _EVAL_2218 <= _EVAL_5247;
    end else if (_EVAL_101) begin
      _EVAL_2218 <= _EVAL_2237;
    end
    _EVAL_2229 <= _EVAL_73;
    _EVAL_2233 <= _EVAL_81;
    _EVAL_2247 <= _EVAL_5;
    _EVAL_2277 <= _EVAL_38;
    if (_EVAL_2741) begin
      _EVAL_2291 <= _EVAL_338;
    end
    if (_EVAL_618) begin
      _EVAL_2293 <= _EVAL_2231;
    end
    if (_EVAL_5699) begin
      _EVAL_2301 <= _EVAL_1374;
    end
    if (_EVAL_916) begin
      _EVAL_2307 <= _EVAL_4088;
    end
    _EVAL_2308 <= _EVAL_111;
    _EVAL_2312 <= _EVAL_146;
    _EVAL_2339 <= _EVAL_125;
    _EVAL_2341 <= _EVAL_58;
    if (_EVAL_5041) begin
      _EVAL_2357 <= _EVAL_1967;
    end
    if (_EVAL_3439) begin
      _EVAL_2360 <= _EVAL_1967;
    end
    _EVAL_2366 <= _EVAL_33;
    if (_EVAL_3705) begin
      _EVAL_2381 <= _EVAL_1374;
    end
    if (_EVAL_2289) begin
      _EVAL_2393 <= _EVAL_3709;
    end
    _EVAL_2422 <= _EVAL_102;
    _EVAL_2444 <= _EVAL_10;
    if (_EVAL_1100) begin
      _EVAL_2462 <= _EVAL_3709;
    end
    _EVAL_2484 <= _EVAL_71;
    if (_EVAL_203) begin
      _EVAL_2490 <= _EVAL_4088;
    end
    if (_EVAL_1589) begin
      _EVAL_2493 <= _EVAL_2231;
    end
    _EVAL_2516 <= _EVAL_84;
    if (_EVAL_2804) begin
      _EVAL_2537 <= _EVAL_4709;
    end
    if (_EVAL_5591) begin
      _EVAL_2546 <= _EVAL_4088;
    end
    if (_EVAL_4610) begin
      _EVAL_2557 <= _EVAL_4088;
    end
    if (_EVAL_2605) begin
      _EVAL_2561 <= _EVAL_4088;
    end
    if (_EVAL_889) begin
      _EVAL_2580 <= _EVAL_338;
    end
    _EVAL_2583 <= _EVAL_53;
    if (_EVAL_1225) begin
      _EVAL_2589 <= _EVAL_338;
    end
    _EVAL_2616 <= _EVAL_80;
    if (_EVAL_1682) begin
      _EVAL_2626 <= _EVAL_4709;
    end
    if (_EVAL_3683) begin
      _EVAL_2629 <= _EVAL_4709;
    end
    if (_EVAL_24) begin
      _EVAL_2667 <= 1'h0;
    end else if (_EVAL_691) begin
      _EVAL_2667 <= _EVAL_338;
    end
    if (_EVAL_874) begin
      _EVAL_2669 <= _EVAL_1967;
    end
    if (_EVAL_3911) begin
      _EVAL_2690 <= _EVAL_1967;
    end
    _EVAL_2717 <= _EVAL_118;
    if (_EVAL_4684) begin
      _EVAL_2766 <= _EVAL_1967;
    end
    _EVAL_2778 <= _EVAL_6;
    if (_EVAL_696) begin
      _EVAL_2781 <= _EVAL_3709;
    end
    _EVAL_2782 <= _EVAL_62;
    if (_EVAL_1669) begin
      _EVAL_2806 <= _EVAL_2231;
    end
    if (_EVAL_2259) begin
      _EVAL_2825 <= _EVAL_1967;
    end
    if (_EVAL_4547) begin
      _EVAL_2827 <= _EVAL_2231;
    end
    if (_EVAL_2407) begin
      _EVAL_2828 <= _EVAL_1967;
    end
    if (_EVAL_4554) begin
      _EVAL_2837 <= _EVAL_338;
    end
    if (_EVAL_2521) begin
      _EVAL_2847 <= _EVAL_3222;
    end
    _EVAL_2876 <= _EVAL_76;
    if (_EVAL_3748) begin
      _EVAL_2889 <= _EVAL_2231;
    end
    _EVAL_2905 <= _EVAL_97;
    _EVAL_2910 <= _EVAL_69;
    if (_EVAL_628) begin
      _EVAL_2918 <= _EVAL_1967;
    end
    if (_EVAL_2057) begin
      _EVAL_2920 <= _EVAL_4709;
    end
    if (_EVAL_4937) begin
      _EVAL_2984 <= _EVAL_3709;
    end
    _EVAL_2988 <= _EVAL_72;
    if (_EVAL_4476) begin
      _EVAL_2993 <= _EVAL_3222;
    end
    if (_EVAL_2265) begin
      _EVAL_3001 <= _EVAL_338;
    end
    if (_EVAL_3530) begin
      _EVAL_3005 <= _EVAL_2231;
    end
    if (_EVAL_5993) begin
      _EVAL_3040 <= _EVAL_4709;
    end
    if (_EVAL_4959) begin
      _EVAL_3062 <= _EVAL_3709;
    end
    if (_EVAL_4676) begin
      _EVAL_3108 <= _EVAL_4709;
    end
    if (_EVAL_5340) begin
      _EVAL_3129 <= _EVAL_3222;
    end
    if (_EVAL_724) begin
      _EVAL_3133 <= _EVAL_1967;
    end
    _EVAL_3152 <= _EVAL_19;
    _EVAL_3171 <= _EVAL_91;
    if (_EVAL_455) begin
      _EVAL_3172 <= _EVAL_3709;
    end
    if (_EVAL_5034) begin
      _EVAL_3173 <= _EVAL_4088;
    end
    _EVAL_3181 <= _EVAL_46;
    if (_EVAL_864) begin
      _EVAL_3194 <= _EVAL_1374;
    end
    if (_EVAL_2660) begin
      _EVAL_3196 <= _EVAL_3222;
    end
    _EVAL_3197 <= _EVAL_96;
    if (_EVAL_2489) begin
      _EVAL_3203 <= _EVAL_1967;
    end
    if (_EVAL_6060) begin
      _EVAL_3213 <= _EVAL_338;
    end
    _EVAL_3225 <= _EVAL_153;
    if (_EVAL_1877) begin
      _EVAL_3234 <= _EVAL_1374;
    end
    if (_EVAL_1851) begin
      _EVAL_3256 <= _EVAL_2231;
    end
    if (_EVAL_5172) begin
      _EVAL_3280 <= _EVAL_3222;
    end
    if (_EVAL_6009) begin
      _EVAL_3286 <= _EVAL_1374;
    end
    if (_EVAL_2020) begin
      _EVAL_3294 <= _EVAL_338;
    end
    if (_EVAL_5022) begin
      _EVAL_3310 <= _EVAL_3709;
    end
    if (_EVAL_5348) begin
      _EVAL_3327 <= _EVAL_338;
    end
    _EVAL_3363 <= _EVAL_133;
    if (_EVAL_367) begin
      _EVAL_3374 <= _EVAL_3222;
    end
    if (_EVAL_5029) begin
      _EVAL_3384 <= _EVAL_1374;
    end
    _EVAL_3404 <= _EVAL_107;
    if (_EVAL_5030) begin
      _EVAL_3429 <= _EVAL_2231;
    end
    if (_EVAL_4013) begin
      _EVAL_3449 <= _EVAL_3709;
    end
    _EVAL_3450 <= _EVAL_114;
    _EVAL_3456 <= _EVAL_149;
    if (_EVAL_1073) begin
      _EVAL_3464 <= _EVAL_3709;
    end
    if (_EVAL_3735) begin
      _EVAL_3467 <= _EVAL_2231;
    end
    if (_EVAL_3389) begin
      _EVAL_3538 <= _EVAL_2231;
    end
    if (_EVAL_3831) begin
      _EVAL_3580 <= _EVAL_338;
    end
    if (_EVAL_5195) begin
      _EVAL_3584 <= _EVAL_3222;
    end
    if (_EVAL_571) begin
      _EVAL_3589 <= _EVAL_338;
    end
    if (_EVAL_5288) begin
      _EVAL_3594 <= _EVAL_338;
    end
    if (_EVAL_4236) begin
      _EVAL_3607 <= _EVAL_3222;
    end
    _EVAL_3609 <= _EVAL_4;
    _EVAL_3629 <= _EVAL_94;
    if (_EVAL_444) begin
      _EVAL_3634 <= _EVAL_1967;
    end
    _EVAL_3639 <= _EVAL_109;
    _EVAL_3652 <= _EVAL_32;
    if (_EVAL_1409) begin
      _EVAL_3673 <= _EVAL_4088;
    end
    if (_EVAL_4696) begin
      _EVAL_3676 <= _EVAL_4088;
    end
    if (_EVAL_4822) begin
      _EVAL_3692 <= _EVAL_4088;
    end
    if (_EVAL_697) begin
      _EVAL_3693 <= _EVAL_3709;
    end
    if (_EVAL_1307) begin
      _EVAL_3722 <= _EVAL_4709;
    end
    if (_EVAL_2829) begin
      _EVAL_3743 <= _EVAL_3709;
    end
    if (_EVAL_968) begin
      _EVAL_3767 <= _EVAL_4709;
    end
    if (_EVAL_1934) begin
      _EVAL_3771 <= _EVAL_4088;
    end
    _EVAL_3783 <= _EVAL_119;
    if (_EVAL_4797) begin
      _EVAL_3789 <= _EVAL_1967;
    end
    _EVAL_3843 <= _EVAL_122;
    _EVAL_3847 <= _EVAL_27;
    if (_EVAL_4449) begin
      _EVAL_3857 <= _EVAL_4088;
    end
    _EVAL_3866 <= _EVAL_3;
    _EVAL_3887 <= _EVAL_23;
    if (_EVAL_4174) begin
      _EVAL_3914 <= _EVAL_1374;
    end
    if (_EVAL_1415) begin
      _EVAL_3940 <= _EVAL_1967;
    end
    if (_EVAL_24) begin
      _EVAL_3945 <= 4'h0;
    end else if (_EVAL_2346) begin
      if (_EVAL_5168) begin
        _EVAL_3945 <= _EVAL_1763;
      end else begin
        _EVAL_3945 <= 4'h8;
      end
    end
    if (_EVAL_3438) begin
      _EVAL_3946 <= _EVAL_338;
    end
    if (_EVAL_2105) begin
      _EVAL_3962 <= _EVAL_338;
    end
    _EVAL_3965 <= _EVAL_44;
    _EVAL_3983 <= _EVAL_14;
    _EVAL_3986 <= _EVAL_35;
    _EVAL_4007 <= _EVAL_139;
    _EVAL_4014 <= _EVAL_70;
    if (_EVAL_3642) begin
      _EVAL_4019 <= _EVAL_3709;
    end
    if (_EVAL_315) begin
      _EVAL_4040 <= _EVAL_4709;
    end
    _EVAL_4045 <= _EVAL_129;
    if (_EVAL_3145) begin
      _EVAL_4051 <= _EVAL_1374;
    end
    _EVAL_4053 <= _EVAL_108;
    if (_EVAL_3590) begin
      _EVAL_4065 <= _EVAL_1967;
    end
    _EVAL_4080 <= _EVAL_65;
    _EVAL_4085 <= _EVAL_148;
    if (_EVAL_5481) begin
      _EVAL_4087 <= _EVAL_1374;
    end
    if (_EVAL_6043) begin
      _EVAL_4103 <= _EVAL_3222;
    end
    if (_EVAL_5894) begin
      _EVAL_4119 <= _EVAL_338;
    end
    if (_EVAL_3561) begin
      _EVAL_4181 <= _EVAL_4709;
    end
    if (_EVAL_3537) begin
      _EVAL_4184 <= _EVAL_3222;
    end
    if (_EVAL_2530) begin
      _EVAL_4233 <= _EVAL_338;
    end
    if (_EVAL_4662) begin
      _EVAL_4264 <= _EVAL_4088;
    end
    _EVAL_4291 <= _EVAL_151;
    if (_EVAL_556) begin
      _EVAL_4304 <= _EVAL_4709;
    end
    _EVAL_4308 <= _EVAL_29;
    _EVAL_4336 <= _EVAL_89;
    _EVAL_4338 <= _EVAL_137;
    if (_EVAL_4117) begin
      _EVAL_4348 <= _EVAL_1374;
    end
    _EVAL_4367 <= _EVAL_99;
    _EVAL_4374 <= _EVAL_21;
    if (_EVAL_3542) begin
      _EVAL_4390 <= _EVAL_4709;
    end
    if (_EVAL_2575) begin
      _EVAL_4397 <= _EVAL_1967;
    end
    if (_EVAL_2861) begin
      _EVAL_4398 <= _EVAL_1967;
    end
    if (_EVAL_488) begin
      _EVAL_4404 <= _EVAL_4709;
    end
    if (_EVAL_3517) begin
      _EVAL_4416 <= _EVAL_2231;
    end
    if (_EVAL_557) begin
      _EVAL_4443 <= _EVAL_3222;
    end
    if (_EVAL_2737) begin
      _EVAL_4479 <= _EVAL_2231;
    end
    if (_EVAL_5833) begin
      _EVAL_4518 <= _EVAL_4709;
    end
    if (_EVAL_5841) begin
      _EVAL_4571 <= _EVAL_3709;
    end
    if (_EVAL_24) begin
      _EVAL_4572 <= 1'h0;
    end else begin
      _EVAL_4572 <= _EVAL_484;
    end
    if (_EVAL_4532) begin
      _EVAL_4574 <= _EVAL_3709;
    end
    _EVAL_4584 <= _EVAL;
    _EVAL_4588 <= _EVAL_104;
    _EVAL_4612 <= _EVAL_110;
    _EVAL_4620 <= _EVAL_41;
    if (_EVAL_1901) begin
      _EVAL_4624 <= _EVAL_4088;
    end
    if (_EVAL_5448) begin
      _EVAL_4631 <= _EVAL_4709;
    end
    if (_EVAL_1982) begin
      _EVAL_4700 <= _EVAL_3709;
    end
    if (_EVAL_2740) begin
      _EVAL_4711 <= _EVAL_4709;
    end
    if (_EVAL_2413) begin
      _EVAL_4732 <= _EVAL_338;
    end
    if (_EVAL_756) begin
      _EVAL_4738 <= _EVAL_3222;
    end
    _EVAL_4742 <= _EVAL_79;
    _EVAL_4779 <= _EVAL_105;
    _EVAL_4785 <= _EVAL_22;
    if (_EVAL_4282) begin
      _EVAL_4786 <= _EVAL_2231;
    end
    _EVAL_4807 <= _EVAL_52;
    if (_EVAL_2421) begin
      _EVAL_4808 <= _EVAL_3222;
    end
    if (_EVAL_5014) begin
      _EVAL_4810 <= _EVAL_3222;
    end
    if (_EVAL_24) begin
      _EVAL_4828 <= 1'h0;
    end else if (_EVAL_2674) begin
      _EVAL_4828 <= _EVAL_1374;
    end else if (_EVAL_176) begin
      _EVAL_4828 <= _EVAL_338;
    end
    _EVAL_4843 <= _EVAL_92;
    if (_EVAL_788) begin
      _EVAL_4908 <= _EVAL_4709;
    end
    if (_EVAL_2935) begin
      _EVAL_4911 <= _EVAL_4709;
    end
    if (_EVAL_6042) begin
      _EVAL_4922 <= _EVAL_1967;
    end
    if (_EVAL_3358) begin
      _EVAL_4927 <= _EVAL_4709;
    end
    if (_EVAL_5539) begin
      _EVAL_4932 <= _EVAL_1374;
    end
    _EVAL_4944 <= _EVAL_152;
    _EVAL_4955 <= _EVAL_48;
    _EVAL_4965 <= _EVAL_117;
    if (_EVAL_1462) begin
      _EVAL_4997 <= _EVAL_3709;
    end
    _EVAL_5002 <= _EVAL_37;
    if (_EVAL_1834) begin
      _EVAL_5008 <= _EVAL_4709;
    end
    if (_EVAL_2622) begin
      _EVAL_5009 <= _EVAL_2231;
    end
    if (_EVAL_3892) begin
      _EVAL_5039 <= _EVAL_2231;
    end
    if (_EVAL_1575) begin
      _EVAL_5080 <= _EVAL_4709;
    end
    if (_EVAL_1949) begin
      _EVAL_5101 <= _EVAL_1374;
    end
    if (_EVAL_810) begin
      _EVAL_5104 <= _EVAL_338;
    end
    if (_EVAL_3030) begin
      _EVAL_5139 <= _EVAL_4088;
    end
    if (_EVAL_5350) begin
      _EVAL_5142 <= _EVAL_3709;
    end
    _EVAL_5147 <= _EVAL_130;
    _EVAL_5163 <= _EVAL_8;
    if (_EVAL_1809) begin
      _EVAL_5190 <= _EVAL_1374;
    end
    if (_EVAL_2510) begin
      _EVAL_5232 <= _EVAL_338;
    end
    _EVAL_5249 <= _EVAL_39;
    if (_EVAL_2025) begin
      _EVAL_5255 <= _EVAL_3222;
    end
    _EVAL_5293 <= _EVAL_7;
    if (_EVAL_283) begin
      _EVAL_5300 <= _EVAL_3222;
    end
    if (_EVAL_4168) begin
      _EVAL_5307 <= _EVAL_338;
    end
    if (_EVAL_678) begin
      _EVAL_5309 <= _EVAL_3222;
    end
    if (_EVAL_5154) begin
      _EVAL_5311 <= _EVAL_2231;
    end
    _EVAL_5315 <= _EVAL_87;
    if (_EVAL_5469) begin
      _EVAL_5345 <= _EVAL_3222;
    end
    _EVAL_5369 <= _EVAL_100;
    _EVAL_5386 <= _EVAL_12;
    if (_EVAL_1325) begin
      _EVAL_5389 <= _EVAL_3709;
    end
    if (_EVAL_2755) begin
      _EVAL_5396 <= _EVAL_1374;
    end
    if (_EVAL_5851) begin
      _EVAL_5409 <= _EVAL_3222;
    end
    _EVAL_5411 <= _EVAL_103;
    if (_EVAL_527) begin
      _EVAL_5479 <= _EVAL_1967;
    end
    if (_EVAL_5802) begin
      _EVAL_5484 <= _EVAL_338;
    end
    if (_EVAL_1451) begin
      _EVAL_5518 <= _EVAL_3709;
    end
    _EVAL_5521 <= _EVAL_63;
    if (_EVAL_3716) begin
      _EVAL_5535 <= _EVAL_3222;
    end
    if (_EVAL_6046) begin
      _EVAL_5537 <= _EVAL_3709;
    end
    if (_EVAL_1532) begin
      _EVAL_5558 <= _EVAL_1967;
    end
    if (_EVAL_2519) begin
      _EVAL_5600 <= _EVAL_338;
    end
    if (_EVAL_156) begin
      _EVAL_5606 <= _EVAL_2231;
    end
    _EVAL_5608 <= _EVAL_2;
    _EVAL_5609 <= _EVAL_83;
    if (_EVAL_892) begin
      _EVAL_5623 <= _EVAL_4088;
    end
    if (_EVAL_4650) begin
      _EVAL_5624 <= _EVAL_3709;
    end
    _EVAL_5629 <= _EVAL_55;
    if (_EVAL_174) begin
      _EVAL_5635 <= _EVAL_1374;
    end
    if (_EVAL_3636) begin
      _EVAL_5665 <= _EVAL_4088;
    end
    if (_EVAL_2611) begin
      _EVAL_5667 <= _EVAL_4709;
    end
    if (_EVAL_3967) begin
      _EVAL_5670 <= _EVAL_4088;
    end
    _EVAL_5675 <= _EVAL_2218 >= _EVAL_1775;
    _EVAL_5684 <= _EVAL_59;
    if (_EVAL_4115) begin
      _EVAL_5696 <= _EVAL_338;
    end
    if (_EVAL_3620) begin
      _EVAL_5697 <= _EVAL_4088;
    end
    if (_EVAL_5331) begin
      _EVAL_5713 <= _EVAL_2231;
    end
    if (_EVAL_1111) begin
      _EVAL_5727 <= _EVAL_4088;
    end
    if (_EVAL_2915) begin
      _EVAL_5735 <= _EVAL_1374;
    end
    _EVAL_5741 <= _EVAL_150;
    _EVAL_5743 <= _EVAL_123;
    if (_EVAL_650) begin
      _EVAL_5765 <= _EVAL_3709;
    end
    if (_EVAL_5957) begin
      _EVAL_5781 <= _EVAL_338;
    end
    _EVAL_5846 <= _EVAL_28;
    if (_EVAL_547) begin
      _EVAL_5878 <= _EVAL_1374;
    end
    _EVAL_5890 <= _EVAL_61;
    if (_EVAL_3104) begin
      _EVAL_5916 <= _EVAL_1374;
    end
    _EVAL_5924 <= _EVAL_143;
    _EVAL_5940 <= _EVAL_126;
    if (_EVAL_463) begin
      _EVAL_5962 <= _EVAL_4088;
    end
    if (_EVAL_6081) begin
      _EVAL_5981 <= _EVAL_4088;
    end
    if (_EVAL_3737) begin
      _EVAL_5985 <= _EVAL_338;
    end
    _EVAL_6021 <= _EVAL_135;
    if (_EVAL_5546) begin
      _EVAL_6030 <= _EVAL_338;
    end
    if (_EVAL_669) begin
      _EVAL_6040 <= _EVAL_2231;
    end
    if (_EVAL_2635) begin
      _EVAL_6098 <= _EVAL_1967;
    end
  end
endmodule
