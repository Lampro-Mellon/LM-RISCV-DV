//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_164_assert(
  input  [2:0]  _EVAL,
  input  [3:0]  _EVAL_0,
  input  [31:0] _EVAL_6,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_15,
  input         _EVAL_19,
  input         _EVAL_21,
  input         _EVAL_24,
  input  [3:0]  _EVAL_25,
  input  [3:0]  _EVAL_26,
  input  [31:0] _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_31,
  input         _EVAL_34,
  input  [1:0]  _EVAL_39,
  input         _EVAL_40,
  input         _EVAL_41,
  input         _EVAL_44,
  input         _EVAL_45,
  input  [2:0]  _EVAL_48,
  input         _EVAL_58,
  input  [3:0]  _EVAL_61,
  input         _EVAL_62,
  input         _EVAL_66,
  input         _EVAL_67,
  input  [2:0]  _EVAL_72,
  input  [1:0]  _EVAL_82,
  input  [3:0]  _EVAL_84,
  input         _EVAL_85,
  input         _EVAL_90,
  input         _EVAL_91,
  input  [2:0]  _EVAL_94,
  input         _EVAL_96,
  input  [3:0]  _EVAL_100,
  input         _EVAL_103,
  input         _EVAL_105,
  input         _EVAL_106
);
  wire  TLMonitor_1__EVAL;
  wire  TLMonitor_1__EVAL_0;
  wire  TLMonitor_1__EVAL_1;
  wire [2:0] TLMonitor_1__EVAL_2;
  wire [2:0] TLMonitor_1__EVAL_3;
  wire [1:0] TLMonitor_1__EVAL_4;
  wire [31:0] TLMonitor_1__EVAL_5;
  wire [3:0] TLMonitor_1__EVAL_6;
  wire  TLMonitor_1__EVAL_7;
  wire  TLMonitor_1__EVAL_8;
  wire  TLMonitor_1__EVAL_9;
  wire  TLMonitor_1__EVAL_10;
  wire  TLMonitor_1__EVAL_11;
  wire [3:0] TLMonitor_1__EVAL_12;
  wire  TLMonitor_1__EVAL_13;
  wire [3:0] TLMonitor_1__EVAL_14;
  wire [2:0] TLMonitor_1__EVAL_15;
  wire  TLMonitor_1__EVAL_16;
  wire  TLMonitor_1__EVAL_17;
  wire  TLMonitor_1__EVAL_18;
  wire  TLMonitor__EVAL;
  wire  TLMonitor__EVAL_0;
  wire  TLMonitor__EVAL_1;
  wire [2:0] TLMonitor__EVAL_2;
  wire [2:0] TLMonitor__EVAL_3;
  wire [1:0] TLMonitor__EVAL_4;
  wire [31:0] TLMonitor__EVAL_5;
  wire [3:0] TLMonitor__EVAL_6;
  wire  TLMonitor__EVAL_7;
  wire  TLMonitor__EVAL_8;
  wire  TLMonitor__EVAL_9;
  wire  TLMonitor__EVAL_10;
  wire  TLMonitor__EVAL_11;
  wire [3:0] TLMonitor__EVAL_12;
  wire  TLMonitor__EVAL_13;
  wire [3:0] TLMonitor__EVAL_14;
  wire [2:0] TLMonitor__EVAL_15;
  wire  TLMonitor__EVAL_16;
  wire  TLMonitor__EVAL_17;
  wire  TLMonitor__EVAL_18;
  _EVAL_163_assert TLMonitor_1 (
    ._EVAL(TLMonitor_1__EVAL),
    ._EVAL_0(TLMonitor_1__EVAL_0),
    ._EVAL_1(TLMonitor_1__EVAL_1),
    ._EVAL_2(TLMonitor_1__EVAL_2),
    ._EVAL_3(TLMonitor_1__EVAL_3),
    ._EVAL_4(TLMonitor_1__EVAL_4),
    ._EVAL_5(TLMonitor_1__EVAL_5),
    ._EVAL_6(TLMonitor_1__EVAL_6),
    ._EVAL_7(TLMonitor_1__EVAL_7),
    ._EVAL_8(TLMonitor_1__EVAL_8),
    ._EVAL_9(TLMonitor_1__EVAL_9),
    ._EVAL_10(TLMonitor_1__EVAL_10),
    ._EVAL_11(TLMonitor_1__EVAL_11),
    ._EVAL_12(TLMonitor_1__EVAL_12),
    ._EVAL_13(TLMonitor_1__EVAL_13),
    ._EVAL_14(TLMonitor_1__EVAL_14),
    ._EVAL_15(TLMonitor_1__EVAL_15),
    ._EVAL_16(TLMonitor_1__EVAL_16),
    ._EVAL_17(TLMonitor_1__EVAL_17),
    ._EVAL_18(TLMonitor_1__EVAL_18)
  );
  _EVAL_163_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14),
    ._EVAL_15(TLMonitor__EVAL_15),
    ._EVAL_16(TLMonitor__EVAL_16),
    ._EVAL_17(TLMonitor__EVAL_17),
    ._EVAL_18(TLMonitor__EVAL_18)
  );
  assign TLMonitor_1__EVAL_11 = _EVAL_105;
  assign TLMonitor_1__EVAL_3 = _EVAL_94;
  assign TLMonitor__EVAL_14 = _EVAL_61;
  assign TLMonitor_1__EVAL_12 = _EVAL_0;
  assign TLMonitor__EVAL_5 = _EVAL_6;
  assign TLMonitor__EVAL_18 = _EVAL_85;
  assign TLMonitor_1__EVAL_6 = _EVAL_26;
  assign TLMonitor__EVAL_11 = _EVAL_105;
  assign TLMonitor_1__EVAL_8 = _EVAL_31;
  assign TLMonitor__EVAL_2 = _EVAL_15;
  assign TLMonitor_1__EVAL_0 = _EVAL_34;
  assign TLMonitor__EVAL_12 = _EVAL_25;
  assign TLMonitor_1__EVAL_15 = _EVAL_72;
  assign TLMonitor_1__EVAL_10 = _EVAL_66;
  assign TLMonitor_1__EVAL_4 = _EVAL_39;
  assign TLMonitor_1__EVAL = _EVAL_45;
  assign TLMonitor_1__EVAL_16 = _EVAL_106;
  assign TLMonitor__EVAL_15 = _EVAL_10;
  assign TLMonitor__EVAL_3 = _EVAL;
  assign TLMonitor_1__EVAL_1 = _EVAL_28;
  assign TLMonitor__EVAL_4 = _EVAL_82;
  assign TLMonitor__EVAL_8 = _EVAL_96;
  assign TLMonitor_1__EVAL_2 = _EVAL_48;
  assign TLMonitor__EVAL_16 = _EVAL_103;
  assign TLMonitor__EVAL_9 = _EVAL_41;
  assign TLMonitor__EVAL_1 = _EVAL_62;
  assign TLMonitor__EVAL_17 = _EVAL_19;
  assign TLMonitor__EVAL_10 = _EVAL_91;
  assign TLMonitor_1__EVAL_18 = _EVAL_85;
  assign TLMonitor_1__EVAL_17 = _EVAL_67;
  assign TLMonitor_1__EVAL_5 = _EVAL_27;
  assign TLMonitor__EVAL_6 = _EVAL_84;
  assign TLMonitor__EVAL_0 = _EVAL_24;
  assign TLMonitor__EVAL = _EVAL_90;
  assign TLMonitor__EVAL_7 = _EVAL_11;
  assign TLMonitor_1__EVAL_14 = _EVAL_100;
  assign TLMonitor_1__EVAL_7 = _EVAL_40;
  assign TLMonitor__EVAL_13 = _EVAL_58;
  assign TLMonitor_1__EVAL_9 = _EVAL_44;
  assign TLMonitor_1__EVAL_13 = _EVAL_21;

endmodule
