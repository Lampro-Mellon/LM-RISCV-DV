//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module SiFive_MemTap(
  output [31:0] mem_0,
  output [31:0] mem_1,
  output [31:0] mem_2,
  output [31:0] mem_3,
  output [31:0] mem_4,
  output [31:0] mem_5,
  output [31:0] mem_6,
  output [31:0] mem_7,
  output [31:0] mem_8,
  output [31:0] mem_9,
  output [31:0] mem_10,
  output [31:0] mem_11,
  output [31:0] mem_12,
  output [31:0] mem_13,
  output [31:0] mem_14,
  output [31:0] mem_15,
  output [31:0] mem_16,
  output [31:0] mem_17,
  output [31:0] mem_18,
  output [31:0] mem_19,
  output [31:0] mem_20,
  output [31:0] mem_21,
  output [31:0] mem_22,
  output [31:0] mem_23,
  output [31:0] mem_24,
  output [31:0] mem_25,
  output [31:0] mem_26,
  output [31:0] mem_27,
  output [31:0] mem_28,
  output [31:0] mem_29,
  output [31:0] mem_30
);
  assign mem_0 = tile.core.rf._EVAL_7[0];
  assign mem_1 = tile.core.rf._EVAL_7[1];
  assign mem_2 = tile.core.rf._EVAL_7[2];
  assign mem_3 = tile.core.rf._EVAL_7[3];
  assign mem_4 = tile.core.rf._EVAL_7[4];
  assign mem_5 = tile.core.rf._EVAL_7[5];
  assign mem_6 = tile.core.rf._EVAL_7[6];
  assign mem_7 = tile.core.rf._EVAL_7[7];
  assign mem_8 = tile.core.rf._EVAL_7[8];
  assign mem_9 = tile.core.rf._EVAL_7[9];
  assign mem_10 = tile.core.rf._EVAL_7[10];
  assign mem_11 = tile.core.rf._EVAL_7[11];
  assign mem_12 = tile.core.rf._EVAL_7[12];
  assign mem_13 = tile.core.rf._EVAL_7[13];
  assign mem_14 = tile.core.rf._EVAL_7[14];
  assign mem_15 = tile.core.rf._EVAL_7[15];
  assign mem_16 = tile.core.rf._EVAL_7[16];
  assign mem_17 = tile.core.rf._EVAL_7[17];
  assign mem_18 = tile.core.rf._EVAL_7[18];
  assign mem_19 = tile.core.rf._EVAL_7[19];
  assign mem_20 = tile.core.rf._EVAL_7[20];
  assign mem_21 = tile.core.rf._EVAL_7[21];
  assign mem_22 = tile.core.rf._EVAL_7[22];
  assign mem_23 = tile.core.rf._EVAL_7[23];
  assign mem_24 = tile.core.rf._EVAL_7[24];
  assign mem_25 = tile.core.rf._EVAL_7[25];
  assign mem_26 = tile.core.rf._EVAL_7[26];
  assign mem_27 = tile.core.rf._EVAL_7[27];
  assign mem_28 = tile.core.rf._EVAL_7[28];
  assign mem_29 = tile.core.rf._EVAL_7[29];
  assign mem_30 = tile.core.rf._EVAL_7[30];
endmodule
