//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_53_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input  [1:0]  _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input  [3:0]  _EVAL_12,
  input  [2:0]  _EVAL_13,
  input  [3:0]  _EVAL_14,
  input         _EVAL_15,
  input  [31:0] _EVAL_16,
  input  [2:0]  _EVAL_17,
  input  [3:0]  _EVAL_18
);
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  reg [31:0] _EVAL_25;
  reg [31:0] _RAND_0;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire [32:0] _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire [3:0] _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire [1:0] _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire [32:0] _EVAL_59;
  wire [32:0] _EVAL_60;
  wire  _EVAL_61;
  wire [32:0] _EVAL_62;
  wire  _EVAL_63;
  wire [5:0] _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire [7:0] _EVAL_69;
  wire [31:0] _EVAL_70;
  wire  _EVAL_71;
  wire [5:0] _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  reg  _EVAL_76;
  reg [31:0] _RAND_1;
  wire  _EVAL_77;
  wire [1:0] _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire [7:0] _EVAL_81;
  wire  _EVAL_82;
  reg [2:0] _EVAL_83;
  reg [31:0] _RAND_2;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire [32:0] _EVAL_87;
  wire  _EVAL_88;
  wire [32:0] _EVAL_89;
  wire  _EVAL_90;
  wire [3:0] _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire [31:0] _EVAL_112;
  wire [31:0] _EVAL_113;
  wire  _EVAL_114;
  reg [2:0] _EVAL_115;
  reg [31:0] _RAND_3;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire [1:0] _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  reg [5:0] _EVAL_122;
  reg [31:0] _RAND_4;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_129;
  wire [7:0] _EVAL_131;
  wire [32:0] _EVAL_132;
  wire  _EVAL_133;
  reg [31:0] _EVAL_134;
  reg [31:0] _RAND_5;
  wire [1:0] _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire [32:0] _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [31:0] _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  reg [3:0] _EVAL_148;
  reg [31:0] _RAND_6;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire [6:0] _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire [32:0] _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  reg  _EVAL_169;
  reg [31:0] _RAND_7;
  wire [32:0] _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [32:0] _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire [32:0] _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire [22:0] _EVAL_191;
  wire  _EVAL_193;
  wire [22:0] _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire [5:0] _EVAL_199;
  wire [32:0] _EVAL_200;
  wire [32:0] _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire [31:0] _EVAL_208;
  wire [32:0] _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire [32:0] _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire [32:0] _EVAL_222;
  wire  _EVAL_223;
  wire [5:0] _EVAL_224;
  reg [1:0] _EVAL_225;
  reg [31:0] _RAND_8;
  wire  _EVAL_226;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire [5:0] _EVAL_233;
  wire  _EVAL_234;
  wire [31:0] _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire [1:0] _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire [6:0] _EVAL_244;
  reg  _EVAL_245;
  reg [31:0] _RAND_9;
  reg  _EVAL_246;
  reg [31:0] _RAND_10;
  wire [32:0] _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire [1:0] _EVAL_252;
  wire  _EVAL_253;
  reg [5:0] _EVAL_254;
  reg [31:0] _RAND_11;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  reg [5:0] _EVAL_258;
  reg [31:0] _RAND_12;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire [7:0] _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  reg [2:0] _EVAL_271;
  reg [31:0] _RAND_13;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  reg  _EVAL_281;
  reg [31:0] _RAND_14;
  wire  _EVAL_282;
  wire [6:0] _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_290;
  wire [32:0] _EVAL_291;
  wire  _EVAL_292;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_293;
  reg [5:0] _EVAL_294;
  reg [31:0] _RAND_15;
  wire  _EVAL_295;
  reg [3:0] _EVAL_296;
  reg [31:0] _RAND_16;
  wire [31:0] _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire [6:0] _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire [3:0] _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire [5:0] _EVAL_310;
  wire  _EVAL_311;
  wire [3:0] _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire [31:0] _EVAL_320;
  wire  _EVAL_321;
  wire  _EVAL_322;
  wire  _EVAL_323;
  wire  _EVAL_324;
  wire  _EVAL_325;
  wire  _EVAL_326;
  wire  _EVAL_328;
  wire  _EVAL_329;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_257 = _EVAL_123 | _EVAL_11;
  assign _EVAL_54 = _EVAL_120 & _EVAL_75;
  assign _EVAL_164 = ~_EVAL_234;
  assign _EVAL_98 = ~_EVAL_49;
  assign _EVAL_273 = _EVAL_23 | _EVAL_11;
  assign _EVAL_174 = $signed(_EVAL_170) & -33'sh1000000;
  assign _EVAL_163 = ~_EVAL_93;
  assign _EVAL_232 = _EVAL_167 | _EVAL_11;
  assign _EVAL_211 = ~_EVAL_107;
  assign _EVAL_68 = ~_EVAL_5;
  assign _EVAL_63 = _EVAL & _EVAL_61;
  assign _EVAL_259 = _EVAL_10 == _EVAL_83;
  assign _EVAL_65 = ~_EVAL_126;
  assign _EVAL_158 = _EVAL_323 | _EVAL_11;
  assign _EVAL_312 = ~_EVAL_306;
  assign _EVAL_146 = _EVAL_277 | _EVAL_216;
  assign _EVAL_133 = _EVAL_108 | _EVAL_11;
  assign _EVAL_103 = _EVAL_329 | _EVAL_41;
  assign _EVAL_190 = ~_EVAL_243;
  assign _EVAL_110 = _EVAL_228 | _EVAL_11;
  assign _EVAL_50 = 2'h1 << _EVAL_166;
  assign _EVAL_20 = _EVAL_122 == 6'h0;
  assign _EVAL_153 = _EVAL_13 <= 3'h1;
  assign _EVAL_295 = _EVAL_293 | _EVAL_11;
  assign _EVAL_200 = _EVAL_174;
  assign _EVAL_171 = _EVAL & _EVAL_88;
  assign _EVAL_89 = {1'b0,$signed(_EVAL_320)};
  assign _EVAL_293 = _EVAL_17 <= 3'h6;
  assign _EVAL_97 = ~_EVAL_282;
  assign _EVAL_309 = _EVAL_12 <= 4'h2;
  assign _EVAL_161 = _EVAL_17[0];
  assign _EVAL_256 = _EVAL_314 | _EVAL_11;
  assign _EVAL_40 = _EVAL_304 | _EVAL_11;
  assign _EVAL_290 = ~_EVAL_142;
  assign _EVAL_121 = $signed(_EVAL_200) == 33'sh0;
  assign _EVAL_72 = _EVAL_154[5:0];
  assign _EVAL_108 = _EVAL_51 | _EVAL_292;
  assign _EVAL_215 = _EVAL_1 == _EVAL_281;
  assign _EVAL_325 = $signed(_EVAL_87) == 33'sh0;
  assign _EVAL_287 = _EVAL_230 | _EVAL_11;
  assign _EVAL_113 = _EVAL_16 ^ 32'h80000000;
  assign _EVAL_278 = ~_EVAL_308;
  assign _EVAL_106 = _EVAL_98 & _EVAL_217;
  assign _EVAL_241 = ~_EVAL_298;
  assign _EVAL_207 = _EVAL_10 == 3'h0;
  assign _EVAL_313 = _EVAL_252[0];
  assign _EVAL_228 = _EVAL_17 == _EVAL_115;
  assign _EVAL_39 = _EVAL_178 & _EVAL_27;
  assign _EVAL_111 = _EVAL_86 | _EVAL_210;
  assign _EVAL_269 = _EVAL_13 == _EVAL_271;
  assign _EVAL_255 = ~_EVAL_82;
  assign _EVAL_288 = ~_EVAL_24;
  assign _EVAL_51 = _EVAL_309 & _EVAL_275;
  assign _EVAL_262 = _EVAL_206 | _EVAL_11;
  assign _EVAL_88 = _EVAL_10 == 3'h7;
  assign _EVAL_36 = _EVAL_49 & _EVAL_217;
  assign _EVAL_55 = ~_EVAL_92;
  assign _EVAL_151 = _EVAL_309 & _EVAL_103;
  assign _EVAL_37 = _EVAL_274 | _EVAL_11;
  assign _EVAL_132 = _EVAL_60;
  assign _EVAL_267 = ~_EVAL_40;
  assign _EVAL_168 = ~_EVAL_217;
  assign _EVAL_202 = _EVAL_250 | _EVAL_11;
  assign _EVAL_311 = ~_EVAL_197;
  assign _EVAL_307 = _EVAL_8 == 2'h0;
  assign _EVAL_165 = ~_EVAL_313;
  assign _EVAL_322 = _EVAL_38 == 4'h0;
  assign _EVAL_117 = ~_EVAL_264;
  assign _EVAL_137 = _EVAL_127 | _EVAL_205;
  assign _EVAL_135 = 2'h1 << _EVAL_6;
  assign _EVAL_70 = _EVAL_16 & _EVAL_112;
  assign _EVAL_236 = _EVAL_198 | _EVAL_66;
  assign _EVAL_251 = ~_EVAL_3;
  assign _EVAL_66 = _EVAL_7 & _EVAL_4;
  assign _EVAL_35 = _EVAL_198 & _EVAL_195;
  assign _EVAL_218 = _EVAL_17 == 3'h1;
  assign _EVAL_266 = _EVAL_196 & _EVAL_288;
  assign _EVAL_73 = _EVAL_294 == 6'h0;
  assign _EVAL_27 = _EVAL_49 & _EVAL_168;
  assign _EVAL_62 = _EVAL_247;
  assign _EVAL_252 = _EVAL_266 ? _EVAL_78 : 2'h0;
  assign _EVAL_102 = _EVAL_85 | _EVAL_54;
  assign _EVAL_222 = $signed(_EVAL_209) & -33'shc000;
  assign _EVAL_243 = _EVAL_185 | _EVAL_11;
  assign _EVAL_303 = _EVAL_136 | _EVAL_11;
  assign _EVAL_205 = _EVAL_309 & _EVAL_41;
  assign _EVAL_48 = _EVAL_66 & _EVAL_67;
  assign _EVAL_157 = {1'b0,$signed(_EVAL_208)};
  assign _EVAL_270 = ~_EVAL_101;
  assign _EVAL_326 = ~_EVAL_144;
  assign _EVAL_223 = _EVAL_178 & _EVAL_106;
  assign _EVAL_69 = _EVAL_191[7:0];
  assign _EVAL_230 = _EVAL_18 == _EVAL_306;
  assign _EVAL_71 = _EVAL_25 < plusarg_reader_out;
  assign _EVAL_154 = _EVAL_294 - 6'h1;
  assign _EVAL_198 = _EVAL_9 & _EVAL;
  assign _EVAL_80 = ~_EVAL_287;
  assign _EVAL_318 = ~_EVAL_279;
  assign _EVAL_109 = _EVAL & _EVAL_261;
  assign _EVAL_56 = _EVAL_21 != _EVAL_313;
  assign _EVAL_141 = ~_EVAL_21;
  assign _EVAL_315 = _EVAL_10[2];
  assign _EVAL_156 = _EVAL_13 <= 3'h4;
  assign _EVAL_118 = _EVAL & _EVAL_44;
  assign _EVAL_261 = _EVAL_10 == 3'h5;
  assign _EVAL_320 = _EVAL_16 ^ 32'h40000000;
  assign _EVAL_216 = _EVAL_319 & _EVAL_98;
  assign _EVAL_194 = 23'hff << _EVAL_14;
  assign _EVAL_233 = _EVAL_81[7:2];
  assign _EVAL_104 = _EVAL_17 == 3'h0;
  assign _EVAL_276 = ~_EVAL_256;
  assign _EVAL_221 = _EVAL_4 & _EVAL_105;
  assign _EVAL_59 = _EVAL_25 + 32'h1;
  assign _EVAL_286 = ~_EVAL_133;
  assign _EVAL_145 = _EVAL_176 | _EVAL_11;
  assign _EVAL_177 = ~_EVAL_11;
  assign _EVAL_253 = ~_EVAL_95;
  assign _EVAL_240 = _EVAL_129 | _EVAL_121;
  assign _EVAL_52 = _EVAL_16 == _EVAL_134;
  assign _EVAL_23 = _EVAL_111 | _EVAL_71;
  assign _EVAL_46 = _EVAL_58 & _EVAL_165;
  assign _EVAL_136 = _EVAL_68 | _EVAL_15;
  assign _EVAL_248 = _EVAL_4 & _EVAL_183;
  assign _EVAL_32 = _EVAL & _EVAL_260;
  assign _EVAL_86 = ~_EVAL_246;
  assign _EVAL_107 = _EVAL_259 | _EVAL_11;
  assign _EVAL_217 = _EVAL_16[0];
  assign _EVAL_206 = _EVAL_8 <= 2'h2;
  assign _EVAL_193 = ~_EVAL_158;
  assign _EVAL_95 = _EVAL_156 | _EVAL_11;
  assign _EVAL_87 = _EVAL_291;
  assign _EVAL_74 = ~_EVAL_15;
  assign _EVAL_44 = _EVAL_10 == 3'h6;
  assign _EVAL_308 = _EVAL_151 | _EVAL_11;
  assign _EVAL_124 = ~_EVAL_202;
  assign _EVAL_324 = ~_EVAL_295;
  assign _EVAL_195 = _EVAL_258 == 6'h0;
  assign _EVAL_167 = ~_EVAL_2;
  assign _EVAL_219 = {1'b0,$signed(_EVAL_16)};
  assign _EVAL_150 = ~_EVAL_100;
  assign _EVAL_210 = plusarg_reader_out == 32'h0;
  assign _EVAL_47 = _EVAL & _EVAL_172;
  assign _EVAL_283 = _EVAL_254 - 6'h1;
  assign _EVAL_183 = _EVAL_17 == 3'h4;
  assign _EVAL_321 = _EVAL_4 & _EVAL_162;
  assign _EVAL_213 = _EVAL & _EVAL_207;
  assign _EVAL_268 = ~_EVAL_69;
  assign _EVAL_155 = _EVAL_14 >= 4'h2;
  assign _EVAL_139 = {1'b0,$signed(_EVAL_235)};
  assign _EVAL_112 = {{24'd0}, _EVAL_268};
  assign _EVAL_204 = _EVAL_10 == 3'h1;
  assign _EVAL_237 = ~_EVAL_145;
  assign _EVAL_224 = _EVAL_300[5:0];
  assign _EVAL_305 = ~_EVAL_37;
  assign _EVAL_292 = _EVAL_184 & _EVAL_325;
  assign _EVAL_22 = _EVAL_251 | _EVAL_11;
  assign _EVAL_317 = ~_EVAL_22;
  assign _EVAL_105 = _EVAL_17 == 3'h2;
  assign _EVAL_300 = _EVAL_122 - 6'h1;
  assign _EVAL_92 = _EVAL_155 | _EVAL_11;
  assign _EVAL_99 = _EVAL_30 | _EVAL_11;
  assign _EVAL_84 = ~_EVAL_67;
  assign _EVAL_170 = {1'b0,$signed(_EVAL_143)};
  assign _EVAL_316 = ~_EVAL_315;
  assign _EVAL_129 = $signed(_EVAL_201) == 33'sh0;
  assign _EVAL_209 = {1'b0,$signed(_EVAL_113)};
  assign _EVAL_244 = _EVAL_258 - 6'h1;
  assign _EVAL_38 = ~_EVAL_18;
  assign _EVAL_247 = $signed(_EVAL_89) & -33'sh2000;
  assign _EVAL_249 = _EVAL_179 | _EVAL_11;
  assign _EVAL_185 = _EVAL_56 | _EVAL_141;
  assign _EVAL_197 = _EVAL_188 | _EVAL_11;
  assign _EVAL_57 = _EVAL_325 | _EVAL_121;
  assign _EVAL_138 = _EVAL_4 & _EVAL_84;
  assign _EVAL_75 = $signed(_EVAL_62) == 33'sh0;
  assign _EVAL_196 = _EVAL_66 & _EVAL_73;
  assign _EVAL_82 = _EVAL_326 | _EVAL_11;
  assign _EVAL_166 = _EVAL_12[0];
  assign _EVAL_176 = _EVAL_13 == 3'h0;
  assign _EVAL_85 = _EVAL_309 & _EVAL_231;
  assign _EVAL_297 = _EVAL_59[31:0];
  assign _EVAL_279 = _EVAL_269 | _EVAL_11;
  assign _EVAL_61 = _EVAL_10 == 3'h2;
  assign _EVAL_186 = $signed(_EVAL_139) & -33'sh2000;
  assign _EVAL_152 = _EVAL_91 == 4'h0;
  assign _EVAL_285 = _EVAL_13 <= 3'h2;
  assign _EVAL_181 = _EVAL_146 | _EVAL_140;
  assign _EVAL_94 = _EVAL_13 != 3'h0;
  assign _EVAL_91 = _EVAL_18 & _EVAL_312;
  assign _EVAL_144 = _EVAL_246 >> _EVAL_6;
  assign _EVAL_149 = ~_EVAL_6;
  assign _EVAL_127 = _EVAL_54 | _EVAL_292;
  assign _EVAL_79 = _EVAL_277 | _EVAL_53;
  assign _EVAL_274 = _EVAL_8 != 2'h2;
  assign _EVAL_100 = _EVAL_149 | _EVAL_11;
  assign _EVAL_29 = ~_EVAL_262;
  assign _EVAL_30 = _EVAL_12 == _EVAL_148;
  assign _EVAL_19 = _EVAL_10 == 3'h4;
  assign _EVAL_328 = _EVAL_153 | _EVAL_11;
  assign _EVAL_31 = ~_EVAL_249;
  assign _EVAL_162 = _EVAL_17 == 3'h5;
  assign _EVAL_178 = _EVAL_119[0];
  assign _EVAL_299 = _EVAL_146 | _EVAL_223;
  assign _EVAL_143 = _EVAL_16 ^ 32'h2000000;
  assign _EVAL_179 = _EVAL_14 == _EVAL_296;
  assign _EVAL_191 = 23'hff << _EVAL_12;
  assign _EVAL_265 = ~_EVAL_43;
  assign _EVAL_41 = $signed(_EVAL_34) == 33'sh0;
  assign _EVAL_78 = 2'h1 << _EVAL_2;
  assign _EVAL_175 = ~_EVAL_110;
  assign _EVAL_93 = _EVAL_96 | _EVAL_11;
  assign _EVAL_53 = _EVAL_319 & _EVAL_49;
  assign _EVAL_301 = ~_EVAL_28;
  assign _EVAL_114 = ~_EVAL_232;
  assign _EVAL_284 = ~_EVAL_257;
  assign _EVAL_242 = _EVAL & _EVAL_204;
  assign _EVAL_34 = _EVAL_186;
  assign _EVAL_24 = _EVAL_17 == 3'h6;
  assign _EVAL_49 = _EVAL_16[1];
  assign _EVAL_64 = _EVAL_283[5:0];
  assign _EVAL_125 = _EVAL_4 & _EVAL_24;
  assign _EVAL_304 = _EVAL_102 | _EVAL_292;
  assign _EVAL_180 = _EVAL_98 & _EVAL_168;
  assign _EVAL_182 = _EVAL_79 | _EVAL_39;
  assign _EVAL_272 = _EVAL_198 & _EVAL_20;
  assign _EVAL_319 = _EVAL_119[1];
  assign _EVAL_282 = _EVAL_322 | _EVAL_11;
  assign _EVAL_280 = _EVAL_2 == _EVAL_76;
  assign _EVAL_229 = ~_EVAL_302;
  assign _EVAL_238 = _EVAL_35 ? _EVAL_135 : 2'h0;
  assign _EVAL_203 = ~_EVAL_220;
  assign _EVAL_96 = _EVAL_6 == _EVAL_245;
  assign _EVAL_260 = _EVAL_10 == 3'h3;
  assign _EVAL_188 = _EVAL_70 == 32'h0;
  assign _EVAL_21 = _EVAL_238[0];
  assign _EVAL_173 = _EVAL_152 | _EVAL_11;
  assign _EVAL_101 = _EVAL_137 | _EVAL_11;
  assign _EVAL_131 = _EVAL_194[7:0];
  assign _EVAL_172 = ~_EVAL_20;
  assign _EVAL_67 = _EVAL_254 == 6'h0;
  assign _EVAL_314 = _EVAL_189 >> _EVAL_2;
  assign _EVAL_264 = _EVAL_94 | _EVAL_11;
  assign _EVAL_142 = _EVAL_74 | _EVAL_11;
  assign _EVAL_214 = ~_EVAL_173;
  assign _EVAL_291 = $signed(_EVAL_157) & -33'sh1000;
  assign _EVAL_140 = _EVAL_178 & _EVAL_180;
  assign _EVAL_220 = _EVAL_215 | _EVAL_11;
  assign _EVAL_184 = _EVAL_12 <= 4'h8;
  assign _EVAL_231 = _EVAL_275 | _EVAL_41;
  assign _EVAL_28 = _EVAL_52 | _EVAL_11;
  assign _EVAL_147 = _EVAL_4 & _EVAL_218;
  assign _EVAL_199 = _EVAL_268[7:2];
  assign _EVAL_275 = _EVAL_240 | _EVAL_33;
  assign _EVAL_45 = _EVAL & _EVAL_19;
  assign _EVAL_187 = ~_EVAL_303;
  assign _EVAL_235 = _EVAL_16 ^ 32'h20000000;
  assign _EVAL_201 = _EVAL_222;
  assign _EVAL_123 = _EVAL_8 == _EVAL_225;
  assign _EVAL_212 = _EVAL_79 | _EVAL_239;
  assign _EVAL_58 = _EVAL_246 | _EVAL_21;
  assign _EVAL_116 = ~_EVAL_273;
  assign _EVAL_250 = _EVAL_13 <= 3'h3;
  assign _EVAL_329 = _EVAL_57 | _EVAL_33;
  assign _EVAL_226 = _EVAL_4 & _EVAL_104;
  assign _EVAL_302 = _EVAL_307 | _EVAL_11;
  assign _EVAL_208 = _EVAL_16 ^ 32'h3000;
  assign _EVAL_90 = ~_EVAL_99;
  assign _EVAL_234 = _EVAL_280 | _EVAL_11;
  assign _EVAL_81 = ~_EVAL_131;
  assign _EVAL_239 = _EVAL_178 & _EVAL_36;
  assign _EVAL_323 = _EVAL_5 == _EVAL_169;
  assign _EVAL_306 = {_EVAL_212,_EVAL_182,_EVAL_299,_EVAL_181};
  assign _EVAL_189 = _EVAL_21 | _EVAL_246;
  assign _EVAL_43 = _EVAL_277 | _EVAL_11;
  assign _EVAL_298 = _EVAL_285 | _EVAL_11;
  assign _EVAL_119 = _EVAL_50 | 2'h1;
  assign _EVAL_77 = ~_EVAL_328;
  assign _EVAL_310 = _EVAL_244[5:0];
  assign _EVAL_120 = _EVAL_12 <= 4'h6;
  assign _EVAL_33 = $signed(_EVAL_132) == 33'sh0;
  assign _EVAL_126 = _EVAL_68 | _EVAL_11;
  assign _EVAL_277 = _EVAL_12 >= 4'h2;
  assign _EVAL_60 = $signed(_EVAL_219) & -33'sh5000;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_25 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_76 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_83 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_115 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_122 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_134 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_148 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_169 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_225 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_245 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_246 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_254 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_258 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_271 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_281 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_294 = _RAND_15[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_296 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_0) begin
    if (_EVAL_11) begin
      _EVAL_25 <= 32'h0;
    end else if (_EVAL_236) begin
      _EVAL_25 <= 32'h0;
    end else begin
      _EVAL_25 <= _EVAL_297;
    end
    if (_EVAL_48) begin
      _EVAL_76 <= _EVAL_2;
    end
    if (_EVAL_272) begin
      _EVAL_83 <= _EVAL_10;
    end
    if (_EVAL_48) begin
      _EVAL_115 <= _EVAL_17;
    end
    if (_EVAL_11) begin
      _EVAL_122 <= 6'h0;
    end else if (_EVAL_198) begin
      if (_EVAL_20) begin
        if (_EVAL_316) begin
          _EVAL_122 <= _EVAL_199;
        end else begin
          _EVAL_122 <= 6'h0;
        end
      end else begin
        _EVAL_122 <= _EVAL_224;
      end
    end
    if (_EVAL_272) begin
      _EVAL_134 <= _EVAL_16;
    end
    if (_EVAL_272) begin
      _EVAL_148 <= _EVAL_12;
    end
    if (_EVAL_48) begin
      _EVAL_169 <= _EVAL_5;
    end
    if (_EVAL_48) begin
      _EVAL_225 <= _EVAL_8;
    end
    if (_EVAL_272) begin
      _EVAL_245 <= _EVAL_6;
    end
    if (_EVAL_11) begin
      _EVAL_246 <= 1'h0;
    end else begin
      _EVAL_246 <= _EVAL_46;
    end
    if (_EVAL_11) begin
      _EVAL_254 <= 6'h0;
    end else if (_EVAL_66) begin
      if (_EVAL_67) begin
        if (_EVAL_161) begin
          _EVAL_254 <= _EVAL_233;
        end else begin
          _EVAL_254 <= 6'h0;
        end
      end else begin
        _EVAL_254 <= _EVAL_64;
      end
    end
    if (_EVAL_11) begin
      _EVAL_258 <= 6'h0;
    end else if (_EVAL_198) begin
      if (_EVAL_195) begin
        if (_EVAL_316) begin
          _EVAL_258 <= _EVAL_199;
        end else begin
          _EVAL_258 <= 6'h0;
        end
      end else begin
        _EVAL_258 <= _EVAL_310;
      end
    end
    if (_EVAL_272) begin
      _EVAL_271 <= _EVAL_13;
    end
    if (_EVAL_48) begin
      _EVAL_281 <= _EVAL_1;
    end
    if (_EVAL_11) begin
      _EVAL_294 <= 6'h0;
    end else if (_EVAL_66) begin
      if (_EVAL_73) begin
        if (_EVAL_161) begin
          _EVAL_294 <= _EVAL_233;
        end else begin
          _EVAL_294 <= 6'h0;
        end
      end else begin
        _EVAL_294 <= _EVAL_72;
      end
    end
    if (_EVAL_48) begin
      _EVAL_296 <= _EVAL_14;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_305) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_265) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_211) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f620f4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_311) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4313905)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73048659)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d638ea3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a57d90a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bff8b648)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_311) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4ffac33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79527ee9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(249ed36b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(634bc176)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a16350da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff032235)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_311) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_31) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_255) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad625f62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be47aba3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_324) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b3b9cc4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(673a8de7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35d36280)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7047f3fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_311) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a90f547)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_311) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f12255b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_301) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcfcb16c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e205a12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdd0dddb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45b949ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_311) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97598747)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0471b4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_265) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ceeb6029)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_305) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_311) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79af1693)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46d571f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6eb91f67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_305) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b52eeb42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_31) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5379f74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b01ae8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e1ab22b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a5d0f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42741129)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_324) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13ddba57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d31ef4bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8793b5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22c3460)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_255) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eef606e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1602382)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_311) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69219bab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99edc7ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70d33460)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cef455b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4554fd86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1848bd55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(485056c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(923737d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c58e501e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_305) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffcd9843)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cab0925e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_311) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(558d7513)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c25ab55d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9af49a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3af52e82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d287d6ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5993dfa7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6e52b22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c22f48fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(830e4bc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(994e5ee3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6c5457e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_311) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(310abcd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(744627c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34b9f105)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c382d4e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_311) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d32e7053)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_311) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffdd95a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_311) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d82f152)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf36d155)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebc31213)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4a9f235)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_311) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a57d2f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbd1de7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_211) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_284) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_265) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6329dd2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae9b751a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(206d14d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_311) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b86b16f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_311) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_284) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f55fa41c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2edbdf5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec6dbcac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fea92950)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_265) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44ba9f37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2938905)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3879979d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9baf7eea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51002750)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d08a293)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_301) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a1f8a09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
