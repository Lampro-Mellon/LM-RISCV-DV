//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_145(
  output [1:0]  _EVAL,
  output [2:0]  _EVAL_0,
  output        _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  output [31:0] _EVAL_4,
  input  [2:0]  _EVAL_5,
  input  [3:0]  _EVAL_6,
  output        _EVAL_7,
  input  [2:0]  _EVAL_8,
  output        _EVAL_9,
  output        _EVAL_10,
  output [1:0]  _EVAL_11,
  output [2:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  output        _EVAL_16,
  output [8:0]  _EVAL_17,
  input  [1:0]  _EVAL_18,
  input  [8:0]  _EVAL_19,
  output        _EVAL_20,
  input  [31:0] _EVAL_21,
  input         _EVAL_22,
  output        _EVAL_23,
  input  [31:0] _EVAL_24,
  output [2:0]  _EVAL_25,
  input         _EVAL_26,
  output [31:0] _EVAL_27,
  output [3:0]  _EVAL_28
);
  wire [8:0] AsyncQueueSink__EVAL;
  wire [3:0] AsyncQueueSink__EVAL_0;
  wire [2:0] AsyncQueueSink__EVAL_1;
  wire [8:0] AsyncQueueSink__EVAL_2;
  wire [3:0] AsyncQueueSink__EVAL_3;
  wire [2:0] AsyncQueueSink__EVAL_4;
  wire  AsyncQueueSink__EVAL_5;
  wire  AsyncQueueSink__EVAL_6;
  wire [2:0] AsyncQueueSink__EVAL_7;
  wire [31:0] AsyncQueueSink__EVAL_8;
  wire [1:0] AsyncQueueSink__EVAL_9;
  wire [31:0] AsyncQueueSink__EVAL_10;
  wire  AsyncQueueSink__EVAL_11;
  wire  AsyncQueueSink__EVAL_12;
  wire  AsyncQueueSink__EVAL_13;
  wire  AsyncQueueSink__EVAL_14;
  wire  AsyncQueueSink__EVAL_15;
  wire  AsyncQueueSink__EVAL_16;
  wire  AsyncQueueSource__EVAL;
  wire  AsyncQueueSource__EVAL_0;
  wire [1:0] AsyncQueueSource__EVAL_1;
  wire [31:0] AsyncQueueSource__EVAL_2;
  wire  AsyncQueueSource__EVAL_3;
  wire  AsyncQueueSource__EVAL_4;
  wire [31:0] AsyncQueueSource__EVAL_5;
  wire  AsyncQueueSource__EVAL_6;
  wire [2:0] AsyncQueueSource__EVAL_7;
  wire [1:0] AsyncQueueSource__EVAL_8;
  wire  AsyncQueueSource__EVAL_9;
  wire  AsyncQueueSource__EVAL_10;
  wire [2:0] AsyncQueueSource__EVAL_11;
  wire  AsyncQueueSource__EVAL_12;
  _EVAL_143 AsyncQueueSink (
    ._EVAL(AsyncQueueSink__EVAL),
    ._EVAL_0(AsyncQueueSink__EVAL_0),
    ._EVAL_1(AsyncQueueSink__EVAL_1),
    ._EVAL_2(AsyncQueueSink__EVAL_2),
    ._EVAL_3(AsyncQueueSink__EVAL_3),
    ._EVAL_4(AsyncQueueSink__EVAL_4),
    ._EVAL_5(AsyncQueueSink__EVAL_5),
    ._EVAL_6(AsyncQueueSink__EVAL_6),
    ._EVAL_7(AsyncQueueSink__EVAL_7),
    ._EVAL_8(AsyncQueueSink__EVAL_8),
    ._EVAL_9(AsyncQueueSink__EVAL_9),
    ._EVAL_10(AsyncQueueSink__EVAL_10),
    ._EVAL_11(AsyncQueueSink__EVAL_11),
    ._EVAL_12(AsyncQueueSink__EVAL_12),
    ._EVAL_13(AsyncQueueSink__EVAL_13),
    ._EVAL_14(AsyncQueueSink__EVAL_14),
    ._EVAL_15(AsyncQueueSink__EVAL_15),
    ._EVAL_16(AsyncQueueSink__EVAL_16)
  );
  _EVAL_144 AsyncQueueSource (
    ._EVAL(AsyncQueueSource__EVAL),
    ._EVAL_0(AsyncQueueSource__EVAL_0),
    ._EVAL_1(AsyncQueueSource__EVAL_1),
    ._EVAL_2(AsyncQueueSource__EVAL_2),
    ._EVAL_3(AsyncQueueSource__EVAL_3),
    ._EVAL_4(AsyncQueueSource__EVAL_4),
    ._EVAL_5(AsyncQueueSource__EVAL_5),
    ._EVAL_6(AsyncQueueSource__EVAL_6),
    ._EVAL_7(AsyncQueueSource__EVAL_7),
    ._EVAL_8(AsyncQueueSource__EVAL_8),
    ._EVAL_9(AsyncQueueSource__EVAL_9),
    ._EVAL_10(AsyncQueueSource__EVAL_10),
    ._EVAL_11(AsyncQueueSource__EVAL_11),
    ._EVAL_12(AsyncQueueSource__EVAL_12)
  );
  assign _EVAL_1 = AsyncQueueSink__EVAL_13;
  assign _EVAL_4 = AsyncQueueSink__EVAL_8;
  assign AsyncQueueSource__EVAL_10 = _EVAL_15;
  assign AsyncQueueSource__EVAL_11 = _EVAL_5;
  assign _EVAL_23 = AsyncQueueSink__EVAL_5;
  assign AsyncQueueSink__EVAL_10 = _EVAL_21;
  assign _EVAL_0 = AsyncQueueSource__EVAL_7;
  assign _EVAL = AsyncQueueSink__EVAL_9;
  assign AsyncQueueSource__EVAL_6 = _EVAL_3;
  assign AsyncQueueSource__EVAL_3 = _EVAL_2;
  assign AsyncQueueSink__EVAL_3 = _EVAL_6;
  assign _EVAL_17 = AsyncQueueSink__EVAL;
  assign AsyncQueueSink__EVAL_16 = _EVAL_22;
  assign _EVAL_27 = AsyncQueueSource__EVAL_2;
  assign AsyncQueueSink__EVAL_14 = _EVAL_26;
  assign AsyncQueueSource__EVAL_8 = _EVAL_18;
  assign AsyncQueueSink__EVAL_2 = _EVAL_19;
  assign AsyncQueueSource__EVAL_5 = _EVAL_24;
  assign _EVAL_16 = AsyncQueueSource__EVAL_12;
  assign AsyncQueueSource__EVAL_4 = _EVAL_22;
  assign _EVAL_12 = AsyncQueueSink__EVAL_4;
  assign AsyncQueueSink__EVAL_11 = _EVAL_3;
  assign _EVAL_20 = AsyncQueueSource__EVAL_0;
  assign _EVAL_11 = AsyncQueueSource__EVAL_1;
  assign AsyncQueueSink__EVAL_7 = _EVAL_8;
  assign AsyncQueueSink__EVAL_6 = _EVAL_13;
  assign _EVAL_7 = AsyncQueueSink__EVAL_15;
  assign _EVAL_28 = AsyncQueueSink__EVAL_0;
  assign _EVAL_25 = AsyncQueueSink__EVAL_1;
  assign AsyncQueueSource__EVAL = _EVAL_14;
  assign _EVAL_10 = AsyncQueueSink__EVAL_12;
  assign _EVAL_9 = AsyncQueueSource__EVAL_9;
endmodule
