//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_152(
  output        _EVAL,
  input  [31:0] _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  output        _EVAL_3,
  output [31:0] _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [31:0] _EVAL_7,
  input  [3:0]  _EVAL_8
);
  wire  _EVAL_9;
  wire [1:0] _EVAL_10;
  wire [15:0] _EVAL_11;
  wire [1:0] _EVAL_12;
  wire [1:0] _EVAL_14;
  wire [62:0] _EVAL_15;
  wire [2:0] _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire [3:0] _EVAL_20;
  wire [1:0] _EVAL_22;
  wire [15:0] _EVAL_23;
  wire [1:0] _EVAL_24;
  wire [1:0] _EVAL_25;
  wire [1:0] _EVAL_26;
  wire [3:0] _EVAL_27;
  wire  _EVAL_28;
  wire [7:0] _EVAL_29;
  wire [3:0] _EVAL_31;
  wire  _EVAL_32;
  wire [1:0] _EVAL_33;
  wire [32:0] _EVAL_34;
  wire [7:0] _EVAL_35;
  wire  _EVAL_36;
  wire [1:0] _EVAL_37;
  wire [64:0] _EVAL_38;
  wire [32:0] _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire [2:0] _EVAL_45;
  reg  _EVAL_46;
  reg [31:0] _RAND_0;
  wire  _EVAL_47;
  wire [1:0] _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire [3:0] _EVAL_53;
  wire [7:0] _EVAL_54;
  wire  _EVAL_55;
  wire [1:0] _EVAL_56;
  wire [1:0] _EVAL_57;
  wire [7:0] _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire [15:0] _EVAL_62;
  wire  _EVAL_63;
  wire [1:0] _EVAL_64;
  wire [15:0] _EVAL_65;
  wire [4:0] _EVAL_66;
  wire [1:0] _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire [6:0] _EVAL_71;
  wire [3:0] _EVAL_72;
  wire  _EVAL_73;
  wire [2:0] _EVAL_74;
  wire [3:0] _EVAL_75;
  wire  _EVAL_76;
  wire [3:0] _EVAL_78;
  wire [3:0] _EVAL_80;
  wire  _EVAL_81;
  reg [32:0] _EVAL_82;
  reg [63:0] _RAND_1;
  wire  _EVAL_83;
  reg [2:0] _EVAL_84;
  reg [31:0] _RAND_2;
  wire  _EVAL_85;
  wire [32:0] _EVAL_86;
  wire [15:0] _EVAL_87;
  wire [1:0] _EVAL_88;
  wire [1:0] _EVAL_89;
  wire  _EVAL_90;
  wire [31:0] _EVAL_91;
  wire [15:0] _EVAL_92;
  wire  _EVAL_94;
  wire [1:0] _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire [1:0] _EVAL_98;
  wire [3:0] _EVAL_99;
  wire [3:0] _EVAL_100;
  wire [15:0] _EVAL_101;
  wire [1:0] _EVAL_102;
  wire [5:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire [1:0] _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire [15:0] _EVAL_109;
  wire [1:0] _EVAL_110;
  wire [1:0] _EVAL_112;
  wire [1:0] _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire [15:0] _EVAL_121;
  wire  _EVAL_122;
  wire [31:0] _EVAL_123;
  wire [1:0] _EVAL_124;
  wire [1:0] _EVAL_125;
  wire  _EVAL_126;
  wire [4:0] _EVAL_128;
  wire [3:0] _EVAL_129;
  wire  _EVAL_130;
  wire [7:0] _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_134;
  wire [1:0] _EVAL_135;
  wire  _EVAL_136;
  wire [3:0] _EVAL_137;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire [15:0] _EVAL_141;
  wire [3:0] _EVAL_142;
  wire [1:0] _EVAL_143;
  wire [3:0] _EVAL_144;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire [31:0] _EVAL_148;
  wire  _EVAL_149;
  wire [31:0] _EVAL_150;
  wire  _EVAL_151;
  wire [3:0] _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire [31:0] _EVAL_158;
  wire [31:0] _EVAL_159;
  reg [65:0] _EVAL_160;
  reg [95:0] _RAND_3;
  reg [5:0] _EVAL_161;
  reg [31:0] _RAND_4;
  wire  _EVAL_162;
  wire [2:0] _EVAL_163;
  wire  _EVAL_164;
  wire [2:0] _EVAL_165;
  wire [2:0] _EVAL_166;
  reg  _EVAL_167;
  reg [31:0] _RAND_5;
  wire  _EVAL_168;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire [4:0] _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_175;
  wire [31:0] _EVAL_176;
  wire [31:0] _EVAL_177;
  wire [1:0] _EVAL_178;
  wire [1:0] _EVAL_179;
  wire [3:0] _EVAL_180;
  wire [1:0] _EVAL_181;
  reg  _EVAL_182;
  reg [31:0] _RAND_6;
  wire [4:0] _EVAL_183;
  wire  _EVAL_184;
  wire [5:0] _EVAL_185;
  wire [3:0] _EVAL_186;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire [1:0] _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_193;
  wire [32:0] _EVAL_194;
  wire [1:0] _EVAL_195;
  wire [2:0] _EVAL_196;
  wire [7:0] _EVAL_197;
  wire [7:0] _EVAL_198;
  wire [1:0] _EVAL_199;
  wire [31:0] _EVAL_200;
  wire [3:0] _EVAL_202;
  wire [62:0] _EVAL_203;
  wire [3:0] _EVAL_204;
  wire [3:0] _EVAL_205;
  wire  _EVAL_207;
  wire [64:0] _EVAL_208;
  wire [1:0] _EVAL_209;
  wire  _EVAL_210;
  wire [2:0] _EVAL_211;
  wire [1:0] _EVAL_212;
  wire [1:0] _EVAL_213;
  wire  _EVAL_214;
  wire [1:0] _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_220;
  wire [3:0] _EVAL_221;
  wire [7:0] _EVAL_222;
  wire [1:0] _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire [2:0] _EVAL_228;
  wire [3:0] _EVAL_229;
  wire [33:0] _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire [2:0] _EVAL_234;
  wire  _EVAL_235;
  wire [3:0] _EVAL_236;
  wire [2:0] _EVAL_237;
  wire [3:0] _EVAL_238;
  wire  _EVAL_239;
  wire [1:0] _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire [1:0] _EVAL_243;
  wire  _EVAL_244;
  wire [2:0] _EVAL_245;
  wire  _EVAL_246;
  assign _EVAL_190 = _EVAL_242 ? 2'h3 : _EVAL_56;
  assign _EVAL_37 = _EVAL_227 ? 2'h2 : {{1'd0}, _EVAL_140};
  assign _EVAL_222 = _EVAL_141[15:8];
  assign _EVAL_221 = _EVAL_35[7:4];
  assign _EVAL_118 = _EVAL_154 & _EVAL_85;
  assign _EVAL_208 = _EVAL_175 ? {{2'd0}, _EVAL_15} : _EVAL_38;
  assign _EVAL_130 = _EVAL_202[3];
  assign _EVAL_244 = _EVAL_27[2];
  assign _EVAL_178 = _EVAL_76 ? 2'h3 : _EVAL_89;
  assign _EVAL_245 = {_EVAL_59,_EVAL_216};
  assign _EVAL_214 = _EVAL_39[32];
  assign _EVAL_74 = {_EVAL_114,_EVAL_106};
  assign _EVAL_29 = _EVAL_23[15:8];
  assign _EVAL_95 = _EVAL_68 ? 2'h3 : _EVAL_113;
  assign _EVAL_16 = _EVAL_69 ? _EVAL_245 : _EVAL_237;
  assign _EVAL_202 = _EVAL_197[7:4];
  assign _EVAL_56 = _EVAL_41 ? 2'h2 : {{1'd0}, _EVAL_17};
  assign _EVAL_12 = _EVAL_63 ? 2'h3 : _EVAL_125;
  assign _EVAL_150 = _EVAL_82[31:0];
  assign _EVAL_158 = _EVAL_160[31:0];
  assign _EVAL_25 = _EVAL_244 ? 2'h2 : {{1'd0}, _EVAL_120};
  assign _EVAL_128 = {_EVAL_19,_EVAL_152};
  assign _EVAL_152 = _EVAL_19 ? _EVAL_229 : _EVAL_144;
  assign _EVAL_170 = _EVAL_75[2];
  assign _EVAL_110 = _EVAL_235 ? 2'h3 : _EVAL_179;
  assign _EVAL_239 = _EVAL_31[1];
  assign _EVAL_165 = {_EVAL_9,_EVAL_22};
  assign _EVAL_151 = _EVAL_238[2];
  assign _EVAL_22 = _EVAL_9 ? _EVAL_110 : _EVAL_10;
  assign _EVAL_106 = _EVAL_114 ? _EVAL_240 : _EVAL_24;
  assign _EVAL_227 = _EVAL_129[2];
  assign _EVAL_88 = _EVAL_70 ? _EVAL_124 : _EVAL_26;
  assign _EVAL_129 = _EVAL_58[7:4];
  assign _EVAL_235 = _EVAL_142[3];
  assign _EVAL = _EVAL_84 == 3'h0;
  assign _EVAL_17 = _EVAL_186[1];
  assign _EVAL_90 = _EVAL_35 != 8'h0;
  assign _EVAL_226 = _EVAL_84 == 3'h3;
  assign _EVAL_230 = _EVAL_86 - _EVAL_82;
  assign _EVAL_104 = _EVAL_3 | _EVAL_1;
  assign _EVAL_121 = _EVAL_0[31:16];
  assign _EVAL_50 = _EVAL_84 == 3'h6;
  assign _EVAL_164 = _EVAL_23 != 16'h0;
  assign _EVAL_199 = _EVAL_147 ? _EVAL_195 : _EVAL_213;
  assign _EVAL_225 = _EVAL_202[1];
  assign _EVAL_47 = _EVAL_221[1];
  assign _EVAL_126 = _EVAL_161 == 6'h20;
  assign _EVAL_31 = _EVAL_58[3:0];
  assign _EVAL_108 = _EVAL_142[2];
  assign _EVAL_97 = _EVAL_20[1];
  assign _EVAL_86 = _EVAL_160[64:32];
  assign _EVAL_212 = _EVAL_122 ? 2'h2 : {{1'd0}, _EVAL_217};
  assign _EVAL_28 = _EVAL_197 != 8'h0;
  assign _EVAL_213 = _EVAL_40 ? 2'h3 : _EVAL_64;
  assign _EVAL_189 = _EVAL_157 != _EVAL_168;
  assign _EVAL_92 = _EVAL_7[15:0];
  assign _EVAL_11 = _EVAL_150[31:16];
  assign _EVAL_112 = _EVAL_116 ? _EVAL_143 : _EVAL_95;
  assign _EVAL_209 = _EVAL_52 ? 2'h3 : _EVAL_181;
  assign _EVAL_23 = _EVAL_158[31:16];
  assign _EVAL_205 = _EVAL_222[3:0];
  assign _EVAL_232 = _EVAL_20[2];
  assign _EVAL_42 = ~_EVAL_46;
  assign _EVAL_153 = _EVAL_157 | _EVAL_168;
  assign _EVAL_200 = _EVAL_160[63:32];
  assign _EVAL_204 = _EVAL_35[3:0];
  assign _EVAL_171 = _EVAL_31[2];
  assign _EVAL_217 = _EVAL_137[1];
  assign _EVAL_116 = _EVAL_180 != 4'h0;
  assign _EVAL_114 = _EVAL_129 != 4'h0;
  assign _EVAL_43 = _EVAL_118 & _EVAL_42;
  assign _EVAL_236 = _EVAL_164 ? _EVAL_72 : _EVAL_99;
  assign _EVAL_122 = _EVAL_137[2];
  assign _EVAL_137 = _EVAL_29[7:4];
  assign _EVAL_113 = _EVAL_136 ? 2'h2 : {{1'd0}, _EVAL_188};
  assign _EVAL_89 = _EVAL_232 ? 2'h2 : {{1'd0}, _EVAL_97};
  assign _EVAL_57 = _EVAL_151 ? 2'h2 : {{1'd0}, _EVAL_193};
  assign _EVAL_4 = {_EVAL_87,_EVAL_101};
  assign _EVAL_63 = _EVAL_80[3];
  assign _EVAL_76 = _EVAL_20[3];
  assign _EVAL_242 = _EVAL_186[3];
  assign _EVAL_20 = _EVAL_29[3:0];
  assign _EVAL_48 = _EVAL_96 ? 2'h2 : {{1'd0}, _EVAL_49};
  assign _EVAL_175 = _EVAL_173 & _EVAL_207;
  assign _EVAL_237 = {_EVAL_119,_EVAL_223};
  assign _EVAL_70 = _EVAL_202 != 4'h0;
  assign _EVAL_32 = _EVAL_78 == 4'h0;
  assign _EVAL_139 = _EVAL_160[31];
  assign _EVAL_185 = _EVAL_66 - _EVAL_128;
  assign _EVAL_210 = _EVAL_75[1];
  assign _EVAL_207 = _EVAL_172 >= 5'h1;
  assign _EVAL_36 = _EVAL_221[3];
  assign _EVAL_180 = _EVAL_198[7:4];
  assign _EVAL_54 = _EVAL_23[7:0];
  assign _EVAL_231 = _EVAL_100 == 4'h2;
  assign _EVAL_188 = _EVAL_53[1];
  assign _EVAL_159 = _EVAL_39[31:0];
  assign _EVAL_228 = {_EVAL_116,_EVAL_112};
  assign _EVAL_59 = _EVAL_137 != 4'h0;
  assign _EVAL_179 = _EVAL_108 ? 2'h2 : {{1'd0}, _EVAL_51};
  assign _EVAL_197 = _EVAL_109[15:8];
  assign _EVAL_136 = _EVAL_53[2];
  assign _EVAL_102 = _EVAL_94 ? 2'h3 : _EVAL_25;
  assign _EVAL_38 = {_EVAL_176,_EVAL_158,_EVAL_85};
  assign _EVAL_166 = _EVAL_28 ? _EVAL_163 : _EVAL_234;
  assign _EVAL_19 = _EVAL_11 != 16'h0;
  assign _EVAL_96 = _EVAL_205[2];
  assign _EVAL_186 = _EVAL_54[3:0];
  assign _EVAL_33 = _EVAL_117 ? 2'h2 : {{1'd0}, _EVAL_47};
  assign _EVAL_203 = {{31'd0}, _EVAL_158};
  assign _EVAL_52 = _EVAL_75[3];
  assign _EVAL_163 = {_EVAL_70,_EVAL_88};
  assign _EVAL_53 = _EVAL_198[3:0];
  assign _EVAL_34 = {_EVAL_168,_EVAL_62,_EVAL_92};
  assign _EVAL_141 = _EVAL_158[15:0];
  assign _EVAL_229 = {_EVAL_90,_EVAL_196};
  assign _EVAL_62 = _EVAL_7[31:16];
  assign _EVAL_81 = _EVAL & _EVAL_2;
  assign _EVAL_123 = _EVAL_182 ? _EVAL_91 : _EVAL_158;
  assign _EVAL_45 = _EVAL_60 ? _EVAL_165 : _EVAL_228;
  assign _EVAL_69 = _EVAL_29 != 8'h0;
  assign _EVAL_120 = _EVAL_27[1];
  assign _EVAL_15 = _EVAL_203 << _EVAL_172;
  assign _EVAL_72 = {_EVAL_69,_EVAL_16};
  assign _EVAL_246 = _EVAL_84 == 3'h1;
  assign _EVAL_9 = _EVAL_142 != 4'h0;
  assign _EVAL_18 = _EVAL_238[3];
  assign _EVAL_85 = ~_EVAL_214;
  assign _EVAL_181 = _EVAL_170 ? 2'h2 : {{1'd0}, _EVAL_210};
  assign _EVAL_26 = _EVAL_18 ? 2'h3 : _EVAL_57;
  assign _EVAL_87 = _EVAL_123[31:16];
  assign _EVAL_220 = _EVAL_137[3];
  assign _EVAL_183 = _EVAL_185[4:0];
  assign _EVAL_24 = _EVAL_146 ? 2'h3 : _EVAL_243;
  assign _EVAL_149 = _EVAL_84 == 3'h5;
  assign _EVAL_117 = _EVAL_221[2];
  assign _EVAL_100 = _EVAL_8 & 4'h2;
  assign _EVAL_41 = _EVAL_186[2];
  assign _EVAL_157 = _EVAL_32 & _EVAL_191;
  assign _EVAL_55 = _EVAL_7[31];
  assign _EVAL_223 = _EVAL_119 ? _EVAL_12 : _EVAL_190;
  assign _EVAL_240 = _EVAL_107 ? 2'h3 : _EVAL_37;
  assign _EVAL_156 = _EVAL_84 == 3'h7;
  assign _EVAL_148 = {_EVAL_121,_EVAL_65};
  assign _EVAL_14 = _EVAL_224 ? 2'h2 : {{1'd0}, _EVAL_225};
  assign _EVAL_195 = _EVAL_36 ? 2'h3 : _EVAL_33;
  assign _EVAL_103 = _EVAL_71[5:0];
  assign _EVAL_154 = _EVAL_161 == 6'h0;
  assign _EVAL_191 = _EVAL_0[31];
  assign _EVAL_78 = _EVAL_8 & 4'h1;
  assign _EVAL_75 = _EVAL_131[7:4];
  assign _EVAL_58 = _EVAL_11[7:0];
  assign _EVAL_65 = _EVAL_0[15:0];
  assign _EVAL_142 = _EVAL_222[7:4];
  assign _EVAL_119 = _EVAL_80 != 4'h0;
  assign _EVAL_135 = _EVAL_115 ? _EVAL_209 : _EVAL_102;
  assign _EVAL_162 = _EVAL_180[2];
  assign _EVAL_147 = _EVAL_221 != 4'h0;
  assign _EVAL_73 = _EVAL_80[2];
  assign _EVAL_49 = _EVAL_205[1];
  assign _EVAL_234 = {_EVAL_115,_EVAL_135};
  assign _EVAL_27 = _EVAL_131[3:0];
  assign _EVAL_68 = _EVAL_53[3];
  assign _EVAL_211 = {_EVAL_147,_EVAL_199};
  assign _EVAL_140 = _EVAL_129[1];
  assign _EVAL_241 = _EVAL_204[1];
  assign _EVAL_64 = _EVAL_134 ? 2'h2 : {{1'd0}, _EVAL_241};
  assign _EVAL_115 = _EVAL_75 != 4'h0;
  assign _EVAL_194 = 32'h0 - _EVAL_123;
  assign _EVAL_243 = _EVAL_171 ? 2'h2 : {{1'd0}, _EVAL_239};
  assign _EVAL_83 = _EVAL_80[1];
  assign _EVAL_184 = _EVAL_82[31];
  assign _EVAL_132 = _EVAL_205[3];
  assign _EVAL_40 = _EVAL_204[3];
  assign _EVAL_51 = _EVAL_142[1];
  assign _EVAL_3 = _EVAL_50 | _EVAL_156;
  assign _EVAL_66 = {_EVAL_164,_EVAL_236};
  assign _EVAL_143 = _EVAL_233 ? 2'h3 : _EVAL_67;
  assign _EVAL_172 = ~_EVAL_183;
  assign _EVAL_107 = _EVAL_129[3];
  assign _EVAL_98 = _EVAL_220 ? 2'h3 : _EVAL_212;
  assign _EVAL_80 = _EVAL_54[7:4];
  assign _EVAL_193 = _EVAL_238[1];
  assign _EVAL_105 = _EVAL_180[1];
  assign _EVAL_94 = _EVAL_27[3];
  assign _EVAL_173 = _EVAL_154 & _EVAL_218;
  assign _EVAL_216 = _EVAL_59 ? _EVAL_98 : _EVAL_178;
  assign _EVAL_134 = _EVAL_204[2];
  assign _EVAL_131 = _EVAL_109[7:0];
  assign _EVAL_125 = _EVAL_73 ? 2'h2 : {{1'd0}, _EVAL_83};
  assign _EVAL_10 = _EVAL_132 ? 2'h3 : _EVAL_48;
  assign _EVAL_39 = _EVAL_230[32:0];
  assign _EVAL_168 = _EVAL_32 & _EVAL_55;
  assign _EVAL_71 = _EVAL_161 + 6'h1;
  assign _EVAL_196 = _EVAL_90 ? _EVAL_211 : _EVAL_74;
  assign _EVAL_60 = _EVAL_222 != 8'h0;
  assign _EVAL_177 = _EVAL_194[31:0];
  assign _EVAL_109 = _EVAL_150[15:0];
  assign _EVAL_67 = _EVAL_162 ? 2'h2 : {{1'd0}, _EVAL_105};
  assign _EVAL_144 = {_EVAL_28,_EVAL_166};
  assign _EVAL_146 = _EVAL_31[3];
  assign _EVAL_99 = {_EVAL_60,_EVAL_45};
  assign _EVAL_218 = ~_EVAL_118;
  assign _EVAL_238 = _EVAL_197[3:0];
  assign _EVAL_224 = _EVAL_202[2];
  assign _EVAL_198 = _EVAL_141[7:0];
  assign _EVAL_233 = _EVAL_180[3];
  assign _EVAL_101 = _EVAL_123[15:0];
  assign _EVAL_91 = _EVAL_160[64:33];
  assign _EVAL_35 = _EVAL_11[15:8];
  assign _EVAL_176 = _EVAL_214 ? _EVAL_200 : _EVAL_159;
  assign _EVAL_124 = _EVAL_130 ? 2'h3 : _EVAL_14;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_46 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  _EVAL_82 = _RAND_1[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_84 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {3{`RANDOM}};
  _EVAL_160 = _RAND_3[65:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_161 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_167 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_182 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_6) begin
    if (_EVAL_81) begin
      _EVAL_46 <= _EVAL_231;
    end
    if (_EVAL_81) begin
      _EVAL_82 <= _EVAL_34;
    end else if (_EVAL_246) begin
      if (_EVAL_184) begin
        _EVAL_82 <= _EVAL_39;
      end
    end
    if (_EVAL_5) begin
      _EVAL_84 <= 3'h0;
    end else if (_EVAL_81) begin
      if (_EVAL_153) begin
        _EVAL_84 <= 3'h1;
      end else begin
        _EVAL_84 <= 3'h3;
      end
    end else if (_EVAL_104) begin
      _EVAL_84 <= 3'h0;
    end else if (_EVAL_226) begin
      if (_EVAL_126) begin
        if (_EVAL_167) begin
          _EVAL_84 <= 3'h5;
        end else begin
          _EVAL_84 <= 3'h7;
        end
      end else if (_EVAL_149) begin
        _EVAL_84 <= 3'h7;
      end else if (_EVAL_246) begin
        _EVAL_84 <= 3'h3;
      end
    end else if (_EVAL_149) begin
      _EVAL_84 <= 3'h7;
    end else if (_EVAL_246) begin
      _EVAL_84 <= 3'h3;
    end
    if (_EVAL_81) begin
      _EVAL_160 <= {{34'd0}, _EVAL_148};
    end else if (_EVAL_226) begin
      _EVAL_160 <= {{1'd0}, _EVAL_208};
    end else if (_EVAL_149) begin
      _EVAL_160 <= {{34'd0}, _EVAL_177};
    end else if (_EVAL_246) begin
      if (_EVAL_139) begin
        _EVAL_160 <= {{34'd0}, _EVAL_177};
      end
    end
    if (_EVAL_81) begin
      _EVAL_161 <= 6'h0;
    end else if (_EVAL_226) begin
      if (_EVAL_175) begin
        _EVAL_161 <= {{1'd0}, _EVAL_172};
      end else begin
        _EVAL_161 <= _EVAL_103;
      end
    end
    if (_EVAL_81) begin
      if (_EVAL_231) begin
        _EVAL_167 <= _EVAL_157;
      end else begin
        _EVAL_167 <= _EVAL_189;
      end
    end else if (_EVAL_226) begin
      if (_EVAL_43) begin
        _EVAL_167 <= 1'h0;
      end
    end
    if (_EVAL_81) begin
      _EVAL_182 <= 1'h0;
    end else if (_EVAL_226) begin
      if (_EVAL_126) begin
        _EVAL_182 <= _EVAL_46;
      end else if (_EVAL_149) begin
        _EVAL_182 <= 1'h0;
      end
    end else if (_EVAL_149) begin
      _EVAL_182 <= 1'h0;
    end
  end
endmodule
