//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_121_assert(
  input  [6:0]  _EVAL_1,
  input         _EVAL_3,
  input         _EVAL_5,
  input         _EVAL_10,
  input         _EVAL_15,
  input  [2:0]  _EVAL_16,
  input  [3:0]  _EVAL_20,
  input         _EVAL_30,
  input         _EVAL_43,
  input         _EVAL_48,
  input         _EVAL_61,
  input         _EVAL_64,
  input         _EVAL_66,
  input         _EVAL_67,
  input         _EVAL_69,
  input         _EVAL_70,
  input         _EVAL_78,
  input         _EVAL_80,
  input         _EVAL_82,
  input         _EVAL_97,
  input  [31:0] _EVAL_101
);
  wire  _EVAL_22;
  wire  TLMonitor__EVAL;
  wire  TLMonitor__EVAL_0;
  wire [3:0] TLMonitor__EVAL_1;
  wire  TLMonitor__EVAL_2;
  wire [2:0] TLMonitor__EVAL_3;
  wire [6:0] TLMonitor__EVAL_4;
  wire [2:0] TLMonitor__EVAL_5;
  wire  TLMonitor__EVAL_6;
  wire  TLMonitor__EVAL_7;
  wire  TLMonitor__EVAL_8;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_35;
  wire  _EVAL_37;
  wire  _EVAL_40;
  wire  _EVAL_45;
  wire  _EVAL_47;
  wire  _EVAL_54;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_63;
  wire  _EVAL_85;
  wire  _EVAL_87;
  wire [8:0] _EVAL_88;
  wire  _EVAL_96;
  wire  _EVAL_102;
  wire [11:0] _EVAL_105;
  wire  _EVAL_107;
  wire  _EVAL_108;
  _EVAL_120_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8)
  );
  assign _EVAL_40 = _EVAL_101[26];
  assign _EVAL_63 = _EVAL_57 & _EVAL_107;
  assign _EVAL_32 = _EVAL_101[29];
  assign _EVAL_45 = _EVAL_57 & _EVAL_67;
  assign _EVAL_54 = ~_EVAL_22;
  assign _EVAL_31 = _EVAL_101[27];
  assign _EVAL_57 = _EVAL_56 & _EVAL_78;
  assign TLMonitor__EVAL = _EVAL_5;
  assign _EVAL_35 = _EVAL_57 & _EVAL_47;
  assign TLMonitor__EVAL_0 = _EVAL_15;
  assign _EVAL_85 = _EVAL_57 & _EVAL_37;
  assign _EVAL_96 = _EVAL_57 & _EVAL_31;
  assign _EVAL_47 = _EVAL_105 != 12'h0;
  assign _EVAL_56 = _EVAL_66 & _EVAL_80;
  assign _EVAL_33 = _EVAL_57 & _EVAL_48;
  assign _EVAL_88 = _EVAL_101[25:17];
  assign _EVAL_107 = _EVAL_101[16];
  assign _EVAL_105 = _EVAL_101[15:4];
  assign _EVAL_87 = _EVAL_57 & _EVAL_32;
  assign TLMonitor__EVAL_5 = _EVAL_16;
  assign _EVAL_37 = _EVAL_88 != 9'h0;
  assign TLMonitor__EVAL_8 = _EVAL_10;
  assign _EVAL_22 = _EVAL_3;
  assign TLMonitor__EVAL_7 = _EVAL_15;
  assign TLMonitor__EVAL_3 = {{2'd0}, _EVAL_80};
  assign TLMonitor__EVAL_4 = _EVAL_1;
  assign _EVAL_108 = _EVAL_57 & _EVAL_40;
  assign TLMonitor__EVAL_2 = _EVAL_5;
  assign TLMonitor__EVAL_6 = _EVAL_3;
  assign TLMonitor__EVAL_1 = _EVAL_20;
  assign _EVAL_102 = _EVAL_57 & _EVAL_30;
  always @(posedge _EVAL_10) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b48c4cb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1d2687e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66e56038)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f072f23f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d241a9cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(890d3ef1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bce6af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec8940c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45d9949e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e526471)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5679099)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f4fca16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39fbe06b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ade4fa1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f7bf715)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad970284)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(633557b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(849417eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2850a86f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(397a6e57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
