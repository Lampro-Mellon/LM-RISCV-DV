//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_103_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input  [3:0]  _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input  [3:0]  _EVAL_8,
  input         _EVAL_9,
  input  [3:0]  _EVAL_10,
  input  [1:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [29:0] _EVAL_13,
  input  [2:0]  _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18
);
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire [29:0] _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire [30:0] _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire [30:0] _EVAL_39;
  wire [5:0] _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  reg [3:0] _EVAL_47;
  reg [31:0] _RAND_0;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  reg [2:0] _EVAL_53;
  reg [31:0] _RAND_1;
  wire [30:0] _EVAL_54;
  wire [32:0] _EVAL_55;
  wire [6:0] _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  reg [5:0] _EVAL_59;
  reg [31:0] _RAND_2;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire [30:0] _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire [4:0] _EVAL_76;
  wire  _EVAL_78;
  reg [2:0] _EVAL_79;
  reg [31:0] _RAND_3;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire [1:0] _EVAL_89;
  wire [7:0] _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_93;
  wire [5:0] _EVAL_94;
  wire [29:0] _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire [3:0] _EVAL_101;
  wire [3:0] _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire [31:0] _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire [30:0] _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire [7:0] _EVAL_117;
  reg  _EVAL_118;
  reg [31:0] _RAND_4;
  wire  _EVAL_119;
  reg [2:0] _EVAL_120;
  reg [31:0] _RAND_5;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire [1:0] _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire [4:0] _EVAL_130;
  wire [7:0] _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire [5:0] _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire [3:0] _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire [22:0] _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire [7:0] _EVAL_155;
  wire  _EVAL_156;
  wire [4:0] _EVAL_157;
  wire [5:0] _EVAL_158;
  wire [4:0] _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  reg [2:0] _EVAL_168;
  reg [31:0] _RAND_6;
  wire [3:0] _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire [29:0] _EVAL_175;
  wire  _EVAL_176;
  wire [7:0] _EVAL_177;
  wire [30:0] _EVAL_178;
  wire [1:0] _EVAL_179;
  wire [30:0] _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire [5:0] _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire [4:0] _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire [6:0] _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire [4:0] _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire [1:0] _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_205;
  wire  _EVAL_206;
  reg [2:0] _EVAL_207;
  reg [31:0] _RAND_7;
  wire [30:0] _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  reg [5:0] _EVAL_212;
  reg [31:0] _RAND_8;
  wire  _EVAL_213;
  wire  _EVAL_214;
  reg [1:0] _EVAL_215;
  reg [31:0] _RAND_9;
  reg [5:0] _EVAL_216;
  reg [31:0] _RAND_10;
  wire  _EVAL_217;
  wire  _EVAL_218;
  reg  _EVAL_219;
  reg [31:0] _RAND_11;
  wire  _EVAL_220;
  wire [29:0] _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire [22:0] _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_231;
  reg [3:0] _EVAL_232;
  reg [31:0] _RAND_12;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire [30:0] _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  reg [29:0] _EVAL_246;
  reg [31:0] _RAND_13;
  wire  _EVAL_247;
  wire  _EVAL_249;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire [7:0] _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire [4:0] _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire [7:0] _EVAL_260;
  wire  _EVAL_261;
  reg [4:0] _EVAL_262;
  reg [31:0] _RAND_14;
  wire  _EVAL_263;
  wire [30:0] _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire [6:0] _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire [30:0] _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire [29:0] _EVAL_293;
  wire [7:0] _EVAL_294;
  reg [5:0] _EVAL_295;
  reg [31:0] _RAND_15;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire [4:0] _EVAL_302;
  reg [31:0] _EVAL_303;
  reg [31:0] _RAND_16;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire [5:0] _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire [30:0] _EVAL_320;
  wire  _EVAL_321;
  wire  _EVAL_322;
  wire  _EVAL_323;
  wire [6:0] _EVAL_324;
  wire  _EVAL_325;
  wire  _EVAL_326;
  wire  _EVAL_327;
  wire  _EVAL_328;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_293 = _EVAL_13 ^ 30'h2000000;
  assign _EVAL_30 = _EVAL_10 == _EVAL_102;
  assign _EVAL_91 = _EVAL_4[0];
  assign _EVAL_290 = $signed(_EVAL_264) == 31'sh0;
  assign _EVAL_282 = _EVAL_303 < plusarg_reader_out;
  assign _EVAL_268 = _EVAL_108 | _EVAL_213;
  assign _EVAL_163 = ~_EVAL_15;
  assign _EVAL_228 = _EVAL_5 <= 3'h2;
  assign _EVAL_210 = _EVAL_153 | _EVAL_74;
  assign _EVAL_318 = ~_EVAL_317;
  assign _EVAL_121 = _EVAL_6 & _EVAL_88;
  assign _EVAL_80 = _EVAL_295 == 6'h0;
  assign _EVAL_110 = _EVAL_55[31:0];
  assign _EVAL_60 = _EVAL_153 | _EVAL_287;
  assign _EVAL_296 = _EVAL_28 | _EVAL_3;
  assign _EVAL_126 = _EVAL_313 & _EVAL_29;
  assign _EVAL_208 = $signed(_EVAL_180) & -31'sh5000;
  assign _EVAL_309 = ~_EVAL_217;
  assign _EVAL_223 = _EVAL_95 == 30'h0;
  assign _EVAL_85 = _EVAL_6 & _EVAL_135;
  assign _EVAL_312 = _EVAL_167 | _EVAL_3;
  assign _EVAL_78 = ~_EVAL_18;
  assign _EVAL_308 = _EVAL_8 >= 4'h2;
  assign _EVAL_58 = _EVAL_122 | _EVAL_3;
  assign _EVAL_218 = ~_EVAL_291;
  assign _EVAL_239 = ~_EVAL_313;
  assign _EVAL_76 = _EVAL_262 | _EVAL_157;
  assign _EVAL_179 = _EVAL_89 | 2'h1;
  assign _EVAL_29 = ~_EVAL_112;
  assign _EVAL_71 = ~_EVAL_199;
  assign _EVAL_157 = _EVAL_155[4:0];
  assign _EVAL_150 = _EVAL_202 & _EVAL_152;
  assign _EVAL_66 = $signed(_EVAL_54) & -31'sh1000000;
  assign _EVAL_127 = ~_EVAL_319;
  assign _EVAL_201 = _EVAL_0 == 3'h1;
  assign _EVAL_270 = ~_EVAL_132;
  assign _EVAL_292 = _EVAL_255 | _EVAL_3;
  assign _EVAL_141 = _EVAL_251 | _EVAL_81;
  assign _EVAL_101 = ~_EVAL_102;
  assign _EVAL_285 = _EVAL_186 | _EVAL_281;
  assign _EVAL_297 = _EVAL_306 | _EVAL_103;
  assign _EVAL_180 = {1'b0,$signed(_EVAL_13)};
  assign _EVAL_249 = _EVAL_142 & _EVAL_198;
  assign _EVAL_225 = 23'hff << _EVAL_8;
  assign _EVAL_267 = _EVAL_46 | _EVAL_3;
  assign _EVAL_253 = _EVAL_225[7:0];
  assign _EVAL_140 = _EVAL_4 == 3'h2;
  assign _EVAL_72 = _EVAL_5 <= 3'h1;
  assign _EVAL_19 = _EVAL_188 | _EVAL_3;
  assign _EVAL_200 = _EVAL_14[2:1];
  assign _EVAL_117 = ~_EVAL_253;
  assign _EVAL_243 = _EVAL_301 | _EVAL_3;
  assign _EVAL_244 = ~_EVAL_292;
  assign _EVAL_289 = plusarg_reader_out == 32'h0;
  assign _EVAL_222 = _EVAL_142 & _EVAL_226;
  assign _EVAL_119 = ~_EVAL_138;
  assign _EVAL_286 = ~_EVAL_206;
  assign _EVAL_229 = ~_EVAL_152;
  assign _EVAL_184 = _EVAL_117[7:2];
  assign _EVAL_274 = ~_EVAL_259;
  assign _EVAL_160 = _EVAL_313 & _EVAL_112;
  assign _EVAL_145 = _EVAL_202 & _EVAL_93;
  assign _EVAL_41 = _EVAL_247 | _EVAL_3;
  assign _EVAL_137 = _EVAL_9 & _EVAL_201;
  assign _EVAL_220 = _EVAL_173 | _EVAL_3;
  assign _EVAL_90 = _EVAL_96 ? _EVAL_294 : 8'h0;
  assign _EVAL_87 = _EVAL_189 & _EVAL_80;
  assign _EVAL_279 = ~_EVAL_310;
  assign _EVAL_84 = _EVAL_106 | _EVAL_233;
  assign _EVAL_161 = ~_EVAL_243;
  assign _EVAL_214 = ~_EVAL_41;
  assign _EVAL_209 = _EVAL_20 | _EVAL_3;
  assign _EVAL_256 = _EVAL_164 | _EVAL_222;
  assign _EVAL_202 = _EVAL & _EVAL_6;
  assign _EVAL_55 = _EVAL_303 + 32'h1;
  assign _EVAL_187 = ~_EVAL_245;
  assign _EVAL_27 = _EVAL_308 | _EVAL_3;
  assign _EVAL_125 = _EVAL_12[2:1];
  assign _EVAL_103 = _EVAL_142 & _EVAL_126;
  assign _EVAL_250 = ~_EVAL_100;
  assign _EVAL_81 = $signed(_EVAL_178) == 31'sh0;
  assign _EVAL_205 = _EVAL_11 == 2'h0;
  assign _EVAL_323 = _EVAL_212 == 6'h0;
  assign _EVAL_86 = ~_EVAL_176;
  assign _EVAL_123 = _EVAL_0 == 3'h2;
  assign _EVAL_22 = ~_EVAL_174;
  assign _EVAL_315 = ~_EVAL_61;
  assign _EVAL_148 = _EVAL_43 | _EVAL_3;
  assign _EVAL_64 = _EVAL_2[0];
  assign _EVAL_35 = _EVAL_231 | _EVAL_3;
  assign _EVAL_128 = _EVAL_115 | _EVAL_3;
  assign _EVAL_325 = _EVAL_5 == _EVAL_79;
  assign _EVAL_63 = _EVAL_266 | _EVAL_290;
  assign _EVAL_144 = 23'hff << _EVAL_2;
  assign _EVAL_36 = _EVAL_238 | _EVAL_3;
  assign _EVAL_193 = _EVAL_216 - 6'h1;
  assign _EVAL_56 = _EVAL_212 - 6'h1;
  assign _EVAL_26 = _EVAL_13 ^ 30'h3000;
  assign _EVAL_302 = _EVAL_90[4:0];
  assign _EVAL_264 = _EVAL_320;
  assign _EVAL_142 = _EVAL_179[0];
  assign _EVAL_99 = _EVAL_125 == 2'h1;
  assign _EVAL_136 = _EVAL_57 | _EVAL_3;
  assign _EVAL_322 = _EVAL_141 | _EVAL_290;
  assign _EVAL_65 = _EVAL_164 | _EVAL_249;
  assign _EVAL_113 = {1'b0,$signed(_EVAL_26)};
  assign _EVAL_28 = _EVAL_11 != 2'h2;
  assign _EVAL_301 = _EVAL_11 == _EVAL_215;
  assign _EVAL_211 = _EVAL_129 | _EVAL_3;
  assign _EVAL_233 = _EVAL_200 == 2'h0;
  assign _EVAL_40 = _EVAL_193[5:0];
  assign _EVAL_169 = ~_EVAL_10;
  assign _EVAL_24 = _EVAL_286 | _EVAL_289;
  assign _EVAL_82 = _EVAL_6 & _EVAL_149;
  assign _EVAL_171 = ~_EVAL_240;
  assign _EVAL_49 = _EVAL_12 == _EVAL_207;
  assign _EVAL_189 = _EVAL_16 & _EVAL_9;
  assign _EVAL_106 = _EVAL_200 == 2'h1;
  assign _EVAL_217 = _EVAL_235 | _EVAL_3;
  assign _EVAL_34 = ~_EVAL_181;
  assign _EVAL_39 = $signed(_EVAL_113) & -31'sh1000;
  assign _EVAL_235 = _EVAL_13 == _EVAL_246;
  assign _EVAL_236 = _EVAL_9 & _EVAL_278;
  assign _EVAL_310 = _EVAL_285 | _EVAL_3;
  assign _EVAL_74 = _EVAL_23 & _EVAL_290;
  assign _EVAL_182 = _EVAL_0 == 3'h0;
  assign _EVAL_203 = _EVAL_8 == _EVAL_232;
  assign _EVAL_153 = _EVAL_304 & _EVAL_170;
  assign _EVAL_190 = _EVAL_76 & _EVAL_257;
  assign _EVAL_114 = _EVAL_9 & _EVAL_52;
  assign _EVAL_327 = _EVAL_14 == _EVAL_168;
  assign _EVAL_172 = _EVAL_9 & _EVAL_258;
  assign _EVAL_291 = _EVAL_305 | _EVAL_3;
  assign _EVAL_240 = _EVAL_228 | _EVAL_3;
  assign _EVAL_44 = ~_EVAL_312;
  assign _EVAL_306 = _EVAL_167 | _EVAL_69;
  assign _EVAL_298 = _EVAL_4 == 3'h6;
  assign _EVAL_139 = _EVAL_10 & _EVAL_101;
  assign _EVAL_265 = _EVAL_325 | _EVAL_3;
  assign _EVAL_196 = _EVAL_9 & _EVAL_182;
  assign _EVAL_206 = _EVAL_262 != 5'h0;
  assign _EVAL_62 = _EVAL_273 & _EVAL_239;
  assign _EVAL_252 = _EVAL_139 == 4'h0;
  assign _EVAL_328 = _EVAL_7 == _EVAL_118;
  assign _EVAL_199 = _EVAL_203 | _EVAL_3;
  assign _EVAL_251 = $signed(_EVAL_32) == 31'sh0;
  assign _EVAL_109 = _EVAL_125 == 2'h0;
  assign _EVAL_88 = _EVAL_4 == 3'h0;
  assign _EVAL_261 = ~_EVAL_67;
  assign _EVAL_173 = _EVAL_2 == _EVAL_47;
  assign _EVAL_54 = {1'b0,$signed(_EVAL_293)};
  assign _EVAL_242 = _EVAL_39;
  assign _EVAL_237 = _EVAL_0 == _EVAL_120;
  assign _EVAL_213 = _EVAL_12 == 3'h4;
  assign _EVAL_269 = ~_EVAL_36;
  assign _EVAL_313 = _EVAL_13[1];
  assign _EVAL_181 = _EVAL_321 | _EVAL_3;
  assign _EVAL_143 = ~_EVAL_146;
  assign _EVAL_271 = ~_EVAL_3;
  assign _EVAL_165 = _EVAL_14 == 3'h4;
  assign _EVAL_112 = _EVAL_13[0];
  assign _EVAL_300 = _EVAL_6 & _EVAL_140;
  assign _EVAL_158 = _EVAL_324[5:0];
  assign _EVAL_311 = ~_EVAL_191;
  assign _EVAL_146 = _EVAL_328 | _EVAL_3;
  assign _EVAL_263 = ~_EVAL_116;
  assign _EVAL_51 = ~_EVAL_298;
  assign _EVAL_50 = ~_EVAL_267;
  assign _EVAL_23 = _EVAL_2 <= 4'h2;
  assign _EVAL_238 = _EVAL_4 == _EVAL_53;
  assign _EVAL_31 = _EVAL_0[2];
  assign _EVAL_116 = _EVAL_327 | _EVAL_3;
  assign _EVAL_25 = _EVAL_142 & _EVAL_160;
  assign _EVAL_226 = _EVAL_239 & _EVAL_29;
  assign _EVAL_314 = _EVAL_276[5:0];
  assign _EVAL_294 = 8'h1 << _EVAL_12;
  assign _EVAL_197 = _EVAL_157 | _EVAL_262;
  assign _EVAL_69 = _EVAL_273 & _EVAL_313;
  assign _EVAL_21 = _EVAL_0 == 3'h7;
  assign _EVAL_260 = 8'h1 << _EVAL_14;
  assign _EVAL_275 = _EVAL_6 & _EVAL_229;
  assign _EVAL_287 = _EVAL_23 & _EVAL_141;
  assign _EVAL_177 = _EVAL_144[7:0];
  assign _EVAL_245 = _EVAL_252 | _EVAL_3;
  assign _EVAL_89 = 2'h1 << _EVAL_64;
  assign _EVAL_131 = ~_EVAL_177;
  assign _EVAL_83 = ~_EVAL_148;
  assign _EVAL_178 = _EVAL_208;
  assign _EVAL_102 = {_EVAL_68,_EVAL_297,_EVAL_65,_EVAL_256};
  assign _EVAL_75 = ~_EVAL_154;
  assign _EVAL_98 = _EVAL_189 | _EVAL_202;
  assign _EVAL_115 = _EVAL_5 != 3'h0;
  assign _EVAL_281 = ~_EVAL_162;
  assign _EVAL_93 = _EVAL_59 == 6'h0;
  assign _EVAL_191 = _EVAL_78 | _EVAL_3;
  assign _EVAL_111 = _EVAL_6 & _EVAL_298;
  assign _EVAL_276 = _EVAL_295 - 6'h1;
  assign _EVAL_122 = _EVAL_23 & _EVAL_63;
  assign _EVAL_43 = _EVAL_18 == _EVAL_219;
  assign _EVAL_135 = _EVAL_4 == 3'h5;
  assign _EVAL_52 = _EVAL_0 == 3'h3;
  assign _EVAL_273 = _EVAL_179[1];
  assign _EVAL_194 = _EVAL_23 & _EVAL_322;
  assign _EVAL_132 = _EVAL_268 | _EVAL_3;
  assign _EVAL_152 = _EVAL_216 == 6'h0;
  assign _EVAL_224 = ~_EVAL_80;
  assign _EVAL_175 = _EVAL_13 ^ 30'h20000000;
  assign _EVAL_32 = _EVAL_66;
  assign _EVAL_149 = _EVAL_4 == 3'h1;
  assign _EVAL_154 = _EVAL_72 | _EVAL_3;
  assign _EVAL_326 = ~_EVAL_211;
  assign _EVAL_162 = _EVAL_157 != 5'h0;
  assign _EVAL_176 = _EVAL_30 | _EVAL_3;
  assign _EVAL_166 = _EVAL_156 | _EVAL_3;
  assign _EVAL_156 = _EVAL_11 <= 2'h2;
  assign _EVAL_159 = _EVAL_262 >> _EVAL_14;
  assign _EVAL_45 = ~_EVAL_166;
  assign _EVAL_192 = ~_EVAL_19;
  assign _EVAL_288 = {1'b0,$signed(_EVAL_175)};
  assign _EVAL_37 = ~_EVAL_35;
  assign _EVAL_304 = _EVAL_2 <= 4'h8;
  assign _EVAL_61 = _EVAL_205 | _EVAL_3;
  assign _EVAL_104 = _EVAL_6 & _EVAL_133;
  assign _EVAL_100 = _EVAL_163 | _EVAL_3;
  assign _EVAL_174 = _EVAL_159[0];
  assign _EVAL_198 = _EVAL_239 & _EVAL_112;
  assign _EVAL_272 = _EVAL_9 & _EVAL_123;
  assign _EVAL_170 = $signed(_EVAL_242) == 31'sh0;
  assign _EVAL_46 = _EVAL_24 | _EVAL_282;
  assign _EVAL_97 = _EVAL_9 & _EVAL_224;
  assign _EVAL_94 = _EVAL_131[7:2];
  assign _EVAL_185 = ~_EVAL_58;
  assign _EVAL_133 = _EVAL_4 == 3'h4;
  assign _EVAL_134 = _EVAL_56[5:0];
  assign _EVAL_138 = _EVAL_49 | _EVAL_3;
  assign _EVAL_316 = ~_EVAL_296;
  assign _EVAL_258 = _EVAL_0 == 3'h6;
  assign _EVAL_255 = _EVAL_84 | _EVAL_165;
  assign _EVAL_259 = _EVAL_237 | _EVAL_3;
  assign _EVAL_151 = ~_EVAL_241;
  assign _EVAL_129 = ~_EVAL_1;
  assign _EVAL_317 = _EVAL_223 | _EVAL_3;
  assign _EVAL_241 = _EVAL_60 | _EVAL_3;
  assign _EVAL_299 = ~_EVAL_128;
  assign _EVAL_231 = _EVAL_4 <= 3'h6;
  assign _EVAL_254 = ~_EVAL_27;
  assign _EVAL_321 = _EVAL_5 <= 3'h4;
  assign _EVAL_42 = _EVAL_5 == 3'h0;
  assign _EVAL_221 = {{22'd0}, _EVAL_131};
  assign _EVAL_277 = ~_EVAL_265;
  assign _EVAL_188 = _EVAL_153 | _EVAL_194;
  assign _EVAL_167 = _EVAL_2 >= 4'h2;
  assign _EVAL_95 = _EVAL_13 & _EVAL_221;
  assign _EVAL_57 = _EVAL_169 == 4'h0;
  assign _EVAL_96 = _EVAL_145 & _EVAL_51;
  assign _EVAL_48 = _EVAL_189 & _EVAL_323;
  assign _EVAL_73 = _EVAL_9 & _EVAL_21;
  assign _EVAL_33 = ~_EVAL_31;
  assign _EVAL_105 = _EVAL_9 & _EVAL_284;
  assign _EVAL_283 = ~_EVAL_227;
  assign _EVAL_186 = _EVAL_157 != _EVAL_302;
  assign _EVAL_20 = _EVAL_78 | _EVAL_1;
  assign _EVAL_130 = _EVAL_197 >> _EVAL_12;
  assign _EVAL_195 = ~_EVAL_220;
  assign _EVAL_155 = _EVAL_48 ? _EVAL_260 : 8'h0;
  assign _EVAL_257 = ~_EVAL_302;
  assign _EVAL_305 = _EVAL_5 <= 3'h3;
  assign _EVAL_266 = _EVAL_307 | _EVAL_81;
  assign _EVAL_319 = _EVAL_42 | _EVAL_3;
  assign _EVAL_284 = _EVAL_0 == 3'h5;
  assign _EVAL_320 = $signed(_EVAL_288) & -31'sh2000;
  assign _EVAL_324 = _EVAL_59 - 6'h1;
  assign _EVAL_67 = _EVAL_210 | _EVAL_3;
  assign _EVAL_68 = _EVAL_306 | _EVAL_25;
  assign _EVAL_164 = _EVAL_167 | _EVAL_62;
  assign _EVAL_234 = ~_EVAL_209;
  assign _EVAL_227 = _EVAL_22 | _EVAL_3;
  assign _EVAL_108 = _EVAL_99 | _EVAL_109;
  assign _EVAL_278 = _EVAL_0 == 3'h4;
  assign _EVAL_307 = _EVAL_170 | _EVAL_251;
  assign _EVAL_70 = ~_EVAL_136;
  assign _EVAL_247 = _EVAL_130[0];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_47 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_53 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_59 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_79 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_118 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_120 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_168 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_207 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_212 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_215 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_216 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_219 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_232 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_246 = _RAND_13[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_262 = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_295 = _RAND_15[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_303 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_17) begin
    if (_EVAL_87) begin
      _EVAL_47 <= _EVAL_2;
    end
    if (_EVAL_150) begin
      _EVAL_53 <= _EVAL_4;
    end
    if (_EVAL_3) begin
      _EVAL_59 <= 6'h0;
    end else if (_EVAL_202) begin
      if (_EVAL_93) begin
        if (_EVAL_91) begin
          _EVAL_59 <= _EVAL_184;
        end else begin
          _EVAL_59 <= 6'h0;
        end
      end else begin
        _EVAL_59 <= _EVAL_158;
      end
    end
    if (_EVAL_87) begin
      _EVAL_79 <= _EVAL_5;
    end
    if (_EVAL_150) begin
      _EVAL_118 <= _EVAL_7;
    end
    if (_EVAL_87) begin
      _EVAL_120 <= _EVAL_0;
    end
    if (_EVAL_87) begin
      _EVAL_168 <= _EVAL_14;
    end
    if (_EVAL_150) begin
      _EVAL_207 <= _EVAL_12;
    end
    if (_EVAL_3) begin
      _EVAL_212 <= 6'h0;
    end else if (_EVAL_189) begin
      if (_EVAL_323) begin
        if (_EVAL_33) begin
          _EVAL_212 <= _EVAL_94;
        end else begin
          _EVAL_212 <= 6'h0;
        end
      end else begin
        _EVAL_212 <= _EVAL_134;
      end
    end
    if (_EVAL_150) begin
      _EVAL_215 <= _EVAL_11;
    end
    if (_EVAL_3) begin
      _EVAL_216 <= 6'h0;
    end else if (_EVAL_202) begin
      if (_EVAL_152) begin
        if (_EVAL_91) begin
          _EVAL_216 <= _EVAL_184;
        end else begin
          _EVAL_216 <= 6'h0;
        end
      end else begin
        _EVAL_216 <= _EVAL_40;
      end
    end
    if (_EVAL_150) begin
      _EVAL_219 <= _EVAL_18;
    end
    if (_EVAL_150) begin
      _EVAL_232 <= _EVAL_8;
    end
    if (_EVAL_87) begin
      _EVAL_246 <= _EVAL_13;
    end
    if (_EVAL_3) begin
      _EVAL_262 <= 5'h0;
    end else begin
      _EVAL_262 <= _EVAL_190;
    end
    if (_EVAL_3) begin
      _EVAL_295 <= 6'h0;
    end else if (_EVAL_189) begin
      if (_EVAL_80) begin
        if (_EVAL_33) begin
          _EVAL_295 <= _EVAL_94;
        end else begin
          _EVAL_295 <= 6'h0;
        end
      end else begin
        _EVAL_295 <= _EVAL_314;
      end
    end
    if (_EVAL_3) begin
      _EVAL_303 <= 32'h0;
    end else if (_EVAL_98) begin
      _EVAL_303 <= 32'h0;
    end else begin
      _EVAL_303 <= _EVAL_110;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fa40640)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_315) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb37614c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7f38a3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(928493d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8283a2b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_316) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4d3bbf0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a735556)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b3e5b7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bd11c33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef72ccf1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24bbc2e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fded497)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(588ee2fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c661c3ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea510d66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8597974)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e044dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b50cd0a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f153b933)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_315) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_316) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76856916)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae542bd9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6a7b77a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2f1b03f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d75f6d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb69f67c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e98919b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8a85551)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(503bd64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78aaf8e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22569d43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dcbc300)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9432dfc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_299) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(832a2f23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_326) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58a01a1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ee41ec8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78e6c073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_311) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(142ac00e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abbdbe1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_315) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a2a8eb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7e138bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f723c44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_326) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88c3a401)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1a4c508)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(781a99a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_326) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f00fc8dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa4ecc49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1be3f668)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84d0092a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2604eba2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(161a701e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d296070e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(288f7fe0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_316) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e54899f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(209fe8e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_315) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5e1b2fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_326) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81d7eb0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62eed0c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31c50a9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_315) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef800dd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e66a53d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28121978)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(809a9c60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61ff4225)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27ffe693)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1df7baef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25cd420f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a307cb1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(616a730b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_315) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a24387cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_315) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8c0d850)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9113b407)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea9e0e51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_326) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d4d2e22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26ba438d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(374a9769)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d97fde5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_315) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df275cb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc494ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_326) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7f53ee8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e797217)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50b3dba2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d70a4bf0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_326) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a88941c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f70d98bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_274) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(531165f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_311) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92cef5d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_299) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_316) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(465b70fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b4dd5c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_326) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9f56510)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(151db744)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48b8e9df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
