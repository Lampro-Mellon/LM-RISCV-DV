//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_67(
  input         _EVAL,
  input  [1:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  output        _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  output        _EVAL_8,
  output        _EVAL_9,
  output [3:0]  _EVAL_10,
  output        _EVAL_11,
  input         _EVAL_12,
  output        _EVAL_13,
  output        _EVAL_14,
  input  [31:0] _EVAL_15,
  input         _EVAL_16,
  input  [2:0]  _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  output        _EVAL_20,
  output [3:0]  _EVAL_21,
  output        _EVAL_22,
  input  [3:0]  _EVAL_23,
  output [2:0]  _EVAL_24,
  output        _EVAL_25,
  output        _EVAL_26,
  output [2:0]  _EVAL_27,
  output        _EVAL_28,
  input  [3:0]  _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  output [3:0]  _EVAL_33,
  output [1:0]  _EVAL_34,
  output [2:0]  _EVAL_35,
  input  [29:0] _EVAL_36,
  input  [3:0]  _EVAL_37,
  output        _EVAL_38,
  output [31:0] _EVAL_39,
  output [29:0] _EVAL_40,
  input  [2:0]  _EVAL_41,
  output [2:0]  _EVAL_42,
  input         _EVAL_43,
  output [31:0] _EVAL_44,
  input         _EVAL_45,
  input  [2:0]  _EVAL_46,
  output [2:0]  _EVAL_47,
  input  [31:0] _EVAL_48
);
  wire  Queue__EVAL;
  wire  Queue__EVAL_0;
  wire  Queue__EVAL_1;
  wire [29:0] Queue__EVAL_2;
  wire [2:0] Queue__EVAL_3;
  wire  Queue__EVAL_4;
  wire [3:0] Queue__EVAL_5;
  wire [2:0] Queue__EVAL_6;
  wire  Queue__EVAL_7;
  wire  Queue__EVAL_8;
  wire  Queue__EVAL_9;
  wire  Queue__EVAL_10;
  wire  Queue__EVAL_11;
  wire  Queue__EVAL_12;
  wire [31:0] Queue__EVAL_13;
  wire  Queue__EVAL_14;
  wire  Queue__EVAL_15;
  wire [3:0] Queue__EVAL_16;
  wire [31:0] Queue__EVAL_17;
  wire [3:0] Queue__EVAL_18;
  wire [2:0] Queue__EVAL_19;
  wire  Queue__EVAL_20;
  wire [29:0] Queue__EVAL_21;
  wire [2:0] Queue__EVAL_22;
  wire [3:0] Queue__EVAL_23;
  wire  Queue__EVAL_24;
  wire  Queue__EVAL_25;
  wire [2:0] Queue__EVAL_26;
  wire [2:0] Queue__EVAL_27;
  wire  Queue__EVAL_28;
  wire  Queue_1__EVAL;
  wire [2:0] Queue_1__EVAL_0;
  wire  Queue_1__EVAL_1;
  wire  Queue_1__EVAL_2;
  wire  Queue_1__EVAL_3;
  wire  Queue_1__EVAL_4;
  wire  Queue_1__EVAL_5;
  wire [3:0] Queue_1__EVAL_6;
  wire  Queue_1__EVAL_7;
  wire [1:0] Queue_1__EVAL_8;
  wire [31:0] Queue_1__EVAL_9;
  wire [1:0] Queue_1__EVAL_10;
  wire [31:0] Queue_1__EVAL_11;
  wire [2:0] Queue_1__EVAL_12;
  wire [3:0] Queue_1__EVAL_13;
  wire  Queue_1__EVAL_14;
  wire  Queue_1__EVAL_15;
  wire [2:0] Queue_1__EVAL_16;
  wire  Queue_1__EVAL_17;
  wire  Queue_1__EVAL_18;
  wire  Queue_1__EVAL_19;
  wire [2:0] Queue_1__EVAL_20;
  _EVAL_65 Queue (
    ._EVAL(Queue__EVAL),
    ._EVAL_0(Queue__EVAL_0),
    ._EVAL_1(Queue__EVAL_1),
    ._EVAL_2(Queue__EVAL_2),
    ._EVAL_3(Queue__EVAL_3),
    ._EVAL_4(Queue__EVAL_4),
    ._EVAL_5(Queue__EVAL_5),
    ._EVAL_6(Queue__EVAL_6),
    ._EVAL_7(Queue__EVAL_7),
    ._EVAL_8(Queue__EVAL_8),
    ._EVAL_9(Queue__EVAL_9),
    ._EVAL_10(Queue__EVAL_10),
    ._EVAL_11(Queue__EVAL_11),
    ._EVAL_12(Queue__EVAL_12),
    ._EVAL_13(Queue__EVAL_13),
    ._EVAL_14(Queue__EVAL_14),
    ._EVAL_15(Queue__EVAL_15),
    ._EVAL_16(Queue__EVAL_16),
    ._EVAL_17(Queue__EVAL_17),
    ._EVAL_18(Queue__EVAL_18),
    ._EVAL_19(Queue__EVAL_19),
    ._EVAL_20(Queue__EVAL_20),
    ._EVAL_21(Queue__EVAL_21),
    ._EVAL_22(Queue__EVAL_22),
    ._EVAL_23(Queue__EVAL_23),
    ._EVAL_24(Queue__EVAL_24),
    ._EVAL_25(Queue__EVAL_25),
    ._EVAL_26(Queue__EVAL_26),
    ._EVAL_27(Queue__EVAL_27),
    ._EVAL_28(Queue__EVAL_28)
  );
  _EVAL_66 Queue_1 (
    ._EVAL(Queue_1__EVAL),
    ._EVAL_0(Queue_1__EVAL_0),
    ._EVAL_1(Queue_1__EVAL_1),
    ._EVAL_2(Queue_1__EVAL_2),
    ._EVAL_3(Queue_1__EVAL_3),
    ._EVAL_4(Queue_1__EVAL_4),
    ._EVAL_5(Queue_1__EVAL_5),
    ._EVAL_6(Queue_1__EVAL_6),
    ._EVAL_7(Queue_1__EVAL_7),
    ._EVAL_8(Queue_1__EVAL_8),
    ._EVAL_9(Queue_1__EVAL_9),
    ._EVAL_10(Queue_1__EVAL_10),
    ._EVAL_11(Queue_1__EVAL_11),
    ._EVAL_12(Queue_1__EVAL_12),
    ._EVAL_13(Queue_1__EVAL_13),
    ._EVAL_14(Queue_1__EVAL_14),
    ._EVAL_15(Queue_1__EVAL_15),
    ._EVAL_16(Queue_1__EVAL_16),
    ._EVAL_17(Queue_1__EVAL_17),
    ._EVAL_18(Queue_1__EVAL_18),
    ._EVAL_19(Queue_1__EVAL_19),
    ._EVAL_20(Queue_1__EVAL_20)
  );
  assign Queue_1__EVAL_7 = _EVAL;
  assign _EVAL_38 = Queue__EVAL_1;
  assign Queue__EVAL_27 = _EVAL_41;
  assign _EVAL_14 = Queue__EVAL_10;
  assign Queue_1__EVAL_19 = _EVAL_18;
  assign Queue_1__EVAL_3 = _EVAL_43;
  assign _EVAL_42 = Queue_1__EVAL_16;
  assign _EVAL_34 = Queue_1__EVAL_8;
  assign Queue__EVAL_4 = _EVAL_30;
  assign _EVAL_28 = Queue_1__EVAL_17;
  assign Queue_1__EVAL_2 = _EVAL_45;
  assign Queue__EVAL_14 = _EVAL_32;
  assign Queue__EVAL_3 = _EVAL_17;
  assign _EVAL_8 = Queue__EVAL;
  assign Queue_1__EVAL_9 = _EVAL_15;
  assign Queue_1__EVAL_20 = _EVAL_46;
  assign Queue__EVAL_21 = _EVAL_36;
  assign Queue__EVAL_25 = _EVAL_6;
  assign Queue__EVAL_7 = _EVAL_43;
  assign Queue__EVAL_23 = _EVAL_37;
  assign Queue__EVAL_24 = _EVAL_4;
  assign Queue_1__EVAL_5 = _EVAL_16;
  assign Queue__EVAL_8 = _EVAL_1;
  assign _EVAL_47 = Queue__EVAL_6;
  assign _EVAL_35 = Queue__EVAL_22;
  assign _EVAL_21 = Queue_1__EVAL_6;
  assign _EVAL_24 = Queue__EVAL_26;
  assign _EVAL_39 = Queue__EVAL_13;
  assign _EVAL_26 = Queue_1__EVAL_14;
  assign Queue_1__EVAL_10 = _EVAL_0;
  assign Queue_1__EVAL_1 = _EVAL_31;
  assign _EVAL_22 = Queue_1__EVAL_4;
  assign Queue_1__EVAL_13 = _EVAL_29;
  assign _EVAL_40 = Queue__EVAL_2;
  assign _EVAL_10 = Queue__EVAL_18;
  assign _EVAL_25 = Queue__EVAL_12;
  assign _EVAL_20 = Queue__EVAL_9;
  assign Queue__EVAL_28 = _EVAL_19;
  assign Queue_1__EVAL_18 = _EVAL_32;
  assign _EVAL_33 = Queue__EVAL_5;
  assign _EVAL_3 = Queue__EVAL_11;
  assign Queue_1__EVAL_0 = _EVAL_7;
  assign Queue__EVAL_20 = _EVAL_12;
  assign Queue__EVAL_19 = _EVAL_5;
  assign Queue__EVAL_17 = _EVAL_48;
  assign _EVAL_13 = Queue_1__EVAL_15;
  assign _EVAL_11 = Queue__EVAL_15;
  assign _EVAL_44 = Queue_1__EVAL_11;
  assign _EVAL_9 = Queue_1__EVAL;
  assign Queue__EVAL_16 = _EVAL_23;
  assign _EVAL_27 = Queue_1__EVAL_12;
  assign Queue__EVAL_0 = _EVAL_2;
endmodule
