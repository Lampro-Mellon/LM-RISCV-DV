//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_6_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [31:0] _EVAL_10,
  input         _EVAL_12,
  input         _EVAL_16,
  input  [1:0]  _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_33,
  input  [3:0]  _EVAL_37,
  input         _EVAL_40,
  input         _EVAL_41,
  input         _EVAL_42,
  input  [3:0]  _EVAL_43,
  input         _EVAL_44,
  input  [2:0]  _EVAL_54,
  input  [2:0]  _EVAL_56,
  input         _EVAL_58,
  input  [2:0]  _EVAL_61,
  input         _EVAL_65,
  input  [3:0]  _EVAL_67,
  input         _EVAL_69,
  input  [2:0]  _EVAL_73,
  input  [31:0] _EVAL_75,
  input         _EVAL_79,
  input  [1:0]  _EVAL_81,
  input         _EVAL_82,
  input         _EVAL_85,
  input  [3:0]  _EVAL_86,
  input         _EVAL_89,
  input  [3:0]  _EVAL_90,
  input         _EVAL_91,
  input         _EVAL_97,
  input  [3:0]  _EVAL_100,
  input         _EVAL_103,
  input         _EVAL_108
);
  wire  TLMonitor__EVAL;
  wire [3:0] TLMonitor__EVAL_0;
  wire  TLMonitor__EVAL_1;
  wire  TLMonitor__EVAL_2;
  wire [2:0] TLMonitor__EVAL_3;
  wire [3:0] TLMonitor__EVAL_4;
  wire  TLMonitor__EVAL_5;
  wire  TLMonitor__EVAL_6;
  wire [3:0] TLMonitor__EVAL_7;
  wire [2:0] TLMonitor__EVAL_8;
  wire  TLMonitor__EVAL_9;
  wire  TLMonitor__EVAL_10;
  wire  TLMonitor__EVAL_11;
  wire  TLMonitor__EVAL_12;
  wire  TLMonitor__EVAL_13;
  wire [1:0] TLMonitor__EVAL_14;
  wire [31:0] TLMonitor__EVAL_15;
  wire  TLMonitor__EVAL_16;
  wire  TLMonitor__EVAL_17;
  wire [2:0] TLMonitor__EVAL_18;
  wire  TLMonitor_1__EVAL;
  wire [3:0] TLMonitor_1__EVAL_0;
  wire  TLMonitor_1__EVAL_1;
  wire  TLMonitor_1__EVAL_2;
  wire [2:0] TLMonitor_1__EVAL_3;
  wire [3:0] TLMonitor_1__EVAL_4;
  wire  TLMonitor_1__EVAL_5;
  wire  TLMonitor_1__EVAL_6;
  wire [3:0] TLMonitor_1__EVAL_7;
  wire [2:0] TLMonitor_1__EVAL_8;
  wire  TLMonitor_1__EVAL_9;
  wire  TLMonitor_1__EVAL_10;
  wire  TLMonitor_1__EVAL_11;
  wire  TLMonitor_1__EVAL_12;
  wire  TLMonitor_1__EVAL_13;
  wire [1:0] TLMonitor_1__EVAL_14;
  wire [31:0] TLMonitor_1__EVAL_15;
  wire  TLMonitor_1__EVAL_16;
  wire  TLMonitor_1__EVAL_17;
  wire [2:0] TLMonitor_1__EVAL_18;
  _EVAL_5_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14),
    ._EVAL_15(TLMonitor__EVAL_15),
    ._EVAL_16(TLMonitor__EVAL_16),
    ._EVAL_17(TLMonitor__EVAL_17),
    ._EVAL_18(TLMonitor__EVAL_18)
  );
  _EVAL_5_assert TLMonitor_1 (
    ._EVAL(TLMonitor_1__EVAL),
    ._EVAL_0(TLMonitor_1__EVAL_0),
    ._EVAL_1(TLMonitor_1__EVAL_1),
    ._EVAL_2(TLMonitor_1__EVAL_2),
    ._EVAL_3(TLMonitor_1__EVAL_3),
    ._EVAL_4(TLMonitor_1__EVAL_4),
    ._EVAL_5(TLMonitor_1__EVAL_5),
    ._EVAL_6(TLMonitor_1__EVAL_6),
    ._EVAL_7(TLMonitor_1__EVAL_7),
    ._EVAL_8(TLMonitor_1__EVAL_8),
    ._EVAL_9(TLMonitor_1__EVAL_9),
    ._EVAL_10(TLMonitor_1__EVAL_10),
    ._EVAL_11(TLMonitor_1__EVAL_11),
    ._EVAL_12(TLMonitor_1__EVAL_12),
    ._EVAL_13(TLMonitor_1__EVAL_13),
    ._EVAL_14(TLMonitor_1__EVAL_14),
    ._EVAL_15(TLMonitor_1__EVAL_15),
    ._EVAL_16(TLMonitor_1__EVAL_16),
    ._EVAL_17(TLMonitor_1__EVAL_17),
    ._EVAL_18(TLMonitor_1__EVAL_18)
  );
  assign TLMonitor_1__EVAL_5 = _EVAL_40;
  assign TLMonitor_1__EVAL_15 = _EVAL_75;
  assign TLMonitor__EVAL_17 = _EVAL_44;
  assign TLMonitor__EVAL_15 = _EVAL_10;
  assign TLMonitor__EVAL_3 = _EVAL_0;
  assign TLMonitor__EVAL_1 = _EVAL_97;
  assign TLMonitor_1__EVAL_3 = _EVAL_1;
  assign TLMonitor__EVAL_13 = _EVAL_91;
  assign TLMonitor_1__EVAL_9 = _EVAL_85;
  assign TLMonitor__EVAL_14 = _EVAL_17;
  assign TLMonitor__EVAL_0 = _EVAL_90;
  assign TLMonitor__EVAL_12 = _EVAL_33;
  assign TLMonitor__EVAL_4 = _EVAL_67;
  assign TLMonitor__EVAL_7 = _EVAL_43;
  assign TLMonitor_1__EVAL_8 = _EVAL_56;
  assign TLMonitor__EVAL_18 = _EVAL_61;
  assign TLMonitor_1__EVAL_12 = _EVAL_33;
  assign TLMonitor_1__EVAL_0 = _EVAL_100;
  assign TLMonitor_1__EVAL_10 = _EVAL_16;
  assign TLMonitor_1__EVAL = _EVAL;
  assign TLMonitor_1__EVAL_14 = _EVAL_81;
  assign TLMonitor__EVAL_11 = _EVAL_30;
  assign TLMonitor_1__EVAL_4 = _EVAL_37;
  assign TLMonitor_1__EVAL_13 = _EVAL_89;
  assign TLMonitor__EVAL_2 = _EVAL_82;
  assign TLMonitor_1__EVAL_11 = _EVAL_12;
  assign TLMonitor__EVAL_9 = _EVAL_69;
  assign TLMonitor__EVAL_5 = _EVAL_40;
  assign TLMonitor_1__EVAL_6 = _EVAL_41;
  assign TLMonitor_1__EVAL_17 = _EVAL_58;
  assign TLMonitor_1__EVAL_1 = _EVAL_65;
  assign TLMonitor__EVAL_6 = _EVAL_103;
  assign TLMonitor_1__EVAL_16 = _EVAL_108;
  assign TLMonitor_1__EVAL_18 = _EVAL_54;
  assign TLMonitor__EVAL_10 = _EVAL_42;
  assign TLMonitor__EVAL = _EVAL_31;
  assign TLMonitor_1__EVAL_7 = _EVAL_86;
  assign TLMonitor__EVAL_8 = _EVAL_73;
  assign TLMonitor_1__EVAL_2 = _EVAL_79;
  assign TLMonitor__EVAL_16 = _EVAL_18;

endmodule
