//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_60_assert(
  input         _EVAL,
  input  [3:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [29:0] _EVAL_10,
  input         _EVAL_11,
  input  [3:0]  _EVAL_12,
  input  [2:0]  _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input  [3:0]  _EVAL_16,
  input  [2:0]  _EVAL_17,
  input  [1:0]  _EVAL_18
);
  wire  _EVAL_19;
  wire  _EVAL_20;
  reg [5:0] _EVAL_22;
  reg [31:0] _RAND_0;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire [29:0] _EVAL_25;
  wire  _EVAL_26;
  wire [3:0] _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  reg [2:0] _EVAL_31;
  reg [31:0] _RAND_1;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire [7:0] _EVAL_41;
  wire  _EVAL_42;
  reg [5:0] _EVAL_43;
  reg [31:0] _RAND_2;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire [6:0] _EVAL_50;
  wire  _EVAL_51;
  wire [5:0] _EVAL_52;
  wire [30:0] _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire [30:0] _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire [1:0] _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_80;
  wire [30:0] _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire [1:0] _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire [4:0] _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  reg [2:0] _EVAL_101;
  reg [31:0] _RAND_3;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_105;
  wire [4:0] _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire [30:0] _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire [31:0] _EVAL_120;
  wire [30:0] _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire [5:0] _EVAL_128;
  wire [5:0] _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire [22:0] _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  reg  _EVAL_139;
  reg [31:0] _RAND_4;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [29:0] _EVAL_143;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire [5:0] _EVAL_147;
  wire [3:0] _EVAL_148;
  reg [5:0] _EVAL_149;
  reg [31:0] _RAND_5;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire [7:0] _EVAL_152;
  wire  _EVAL_153;
  reg [2:0] _EVAL_154;
  reg [31:0] _RAND_6;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire [7:0] _EVAL_161;
  wire [30:0] _EVAL_162;
  wire [4:0] _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  reg [2:0] _EVAL_167;
  reg [31:0] _RAND_7;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  reg [31:0] _EVAL_171;
  reg [31:0] _RAND_8;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [4:0] _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire [4:0] _EVAL_178;
  wire  _EVAL_179;
  wire [32:0] _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  reg [29:0] _EVAL_183;
  reg [31:0] _RAND_9;
  wire  _EVAL_184;
  wire [1:0] _EVAL_185;
  wire  _EVAL_186;
  wire [30:0] _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire [30:0] _EVAL_191;
  wire [3:0] _EVAL_192;
  wire [30:0] _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire [7:0] _EVAL_200;
  wire [31:0] plusarg_reader_out;
  wire [29:0] _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  reg  _EVAL_213;
  reg [31:0] _RAND_10;
  wire [29:0] _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire [1:0] _EVAL_217;
  wire  _EVAL_218;
  reg [3:0] _EVAL_219;
  reg [31:0] _RAND_11;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire [30:0] _EVAL_229;
  wire [7:0] _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire [6:0] _EVAL_234;
  wire  _EVAL_235;
  wire [30:0] _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire [4:0] _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire [30:0] _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  reg [4:0] _EVAL_256;
  reg [31:0] _RAND_12;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  reg [5:0] _EVAL_264;
  reg [31:0] _RAND_13;
  wire  _EVAL_265;
  reg [2:0] _EVAL_266;
  reg [31:0] _RAND_14;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire [6:0] _EVAL_282;
  wire  _EVAL_283;
  reg [3:0] _EVAL_284;
  reg [31:0] _RAND_15;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire [7:0] _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire [29:0] _EVAL_297;
  reg [1:0] _EVAL_298;
  reg [31:0] _RAND_16;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire [5:0] _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire [4:0] _EVAL_310;
  wire [6:0] _EVAL_311;
  wire [7:0] _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire [7:0] _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire  _EVAL_318;
  wire [22:0] _EVAL_319;
  wire  _EVAL_320;
  wire  _EVAL_321;
  wire [3:0] _EVAL_322;
  wire [5:0] _EVAL_323;
  wire  _EVAL_324;
  wire  _EVAL_325;
  wire  _EVAL_326;
  wire  _EVAL_327;
  wire [4:0] _EVAL_328;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_231 = ~_EVAL_247;
  assign _EVAL_224 = _EVAL_116 | _EVAL_7;
  assign _EVAL_321 = ~_EVAL_194;
  assign _EVAL_237 = _EVAL_221 | _EVAL_7;
  assign _EVAL_281 = _EVAL_0 >= 4'h2;
  assign _EVAL_180 = _EVAL_171 + 32'h1;
  assign _EVAL_288 = _EVAL_38 & _EVAL_321;
  assign _EVAL_158 = _EVAL_228 & _EVAL_157;
  assign _EVAL_226 = _EVAL_1 & _EVAL_85;
  assign _EVAL_238 = _EVAL_98[0];
  assign _EVAL_229 = {1'b0,$signed(_EVAL_214)};
  assign _EVAL_145 = ~_EVAL_124;
  assign _EVAL_236 = {1'b0,$signed(_EVAL_25)};
  assign _EVAL_65 = $signed(_EVAL_236) & -31'sh1000000;
  assign _EVAL_170 = _EVAL_264 == 6'h0;
  assign _EVAL_28 = _EVAL_322 == 4'h0;
  assign _EVAL_98 = _EVAL_256 >> _EVAL_13;
  assign _EVAL_143 = _EVAL_10 ^ 30'h20000000;
  assign _EVAL_249 = ~_EVAL_283;
  assign _EVAL_181 = ~_EVAL_289;
  assign _EVAL_122 = _EVAL_181 | _EVAL_119;
  assign _EVAL_114 = _EVAL_65;
  assign _EVAL_293 = _EVAL_328[0];
  assign _EVAL_40 = _EVAL_1 & _EVAL_253;
  assign _EVAL_34 = ~_EVAL_137;
  assign _EVAL_87 = $signed(_EVAL_121) == 31'sh0;
  assign _EVAL_164 = ~_EVAL_210;
  assign _EVAL_279 = _EVAL_94 == 2'h1;
  assign _EVAL_323 = _EVAL_234[5:0];
  assign _EVAL_173 = _EVAL_258 | _EVAL_244;
  assign _EVAL_134 = _EVAL_190 | _EVAL_7;
  assign _EVAL_275 = _EVAL_3 == 3'h2;
  assign _EVAL_83 = _EVAL_206 | _EVAL_7;
  assign _EVAL_196 = _EVAL_67 | _EVAL_7;
  assign _EVAL_97 = _EVAL_12 <= 4'h2;
  assign _EVAL_109 = ~_EVAL_4;
  assign _EVAL_318 = _EVAL_16 == _EVAL_192;
  assign _EVAL_129 = _EVAL_50[5:0];
  assign _EVAL_276 = _EVAL_17 <= 3'h3;
  assign _EVAL_261 = ~_EVAL_265;
  assign _EVAL_127 = _EVAL_222 | _EVAL_243;
  assign _EVAL_128 = _EVAL_312[7:2];
  assign _EVAL_50 = _EVAL_43 - 6'h1;
  assign _EVAL_23 = ~_EVAL_68;
  assign _EVAL_198 = _EVAL_15 & _EVAL_220;
  assign _EVAL_242 = _EVAL_15 & _EVAL_138;
  assign _EVAL_78 = ~_EVAL_45;
  assign _EVAL_192 = {_EVAL_42,_EVAL_62,_EVAL_117,_EVAL_127};
  assign _EVAL_91 = ~_EVAL_83;
  assign _EVAL_244 = ~_EVAL_169;
  assign _EVAL_325 = _EVAL_0 == _EVAL_219;
  assign _EVAL_166 = _EVAL_217 == 2'h0;
  assign _EVAL_115 = ~_EVAL_212;
  assign _EVAL_163 = _EVAL_310 | _EVAL_256;
  assign _EVAL_26 = _EVAL_3 == 3'h0;
  assign _EVAL_70 = _EVAL_17 <= 3'h2;
  assign _EVAL_175 = _EVAL_9 == _EVAL_101;
  assign _EVAL_117 = _EVAL_222 | _EVAL_158;
  assign _EVAL_57 = ~_EVAL_218;
  assign _EVAL_312 = ~_EVAL_161;
  assign _EVAL_286 = ~_EVAL_134;
  assign _EVAL_186 = _EVAL_6 == 3'h4;
  assign _EVAL_306 = _EVAL_33 | _EVAL_7;
  assign _EVAL_202 = _EVAL_10 & _EVAL_297;
  assign _EVAL_270 = _EVAL_15 & _EVAL_186;
  assign _EVAL_136 = _EVAL_179 | _EVAL_7;
  assign _EVAL_69 = _EVAL_257 | _EVAL_7;
  assign _EVAL_19 = _EVAL_216 | _EVAL_7;
  assign _EVAL_294 = _EVAL_326 | _EVAL_7;
  assign _EVAL_245 = _EVAL_152[4:0];
  assign _EVAL_108 = ~_EVAL_153;
  assign _EVAL_95 = _EVAL_88 | _EVAL_166;
  assign _EVAL_322 = _EVAL_16 & _EVAL_148;
  assign _EVAL_314 = _EVAL_103 | _EVAL_7;
  assign _EVAL_52 = _EVAL_292[7:2];
  assign _EVAL_38 = _EVAL_273 & _EVAL_75;
  assign _EVAL_58 = _EVAL_173 | _EVAL_7;
  assign _EVAL_72 = _EVAL_15 & _EVAL_194;
  assign _EVAL_93 = _EVAL_278 | _EVAL_7;
  assign _EVAL_85 = _EVAL_3 == 3'h1;
  assign _EVAL_302 = _EVAL_6 == 3'h1;
  assign _EVAL_320 = _EVAL_97 & _EVAL_111;
  assign _EVAL_310 = _EVAL_41[4:0];
  assign _EVAL_326 = _EVAL_327 | _EVAL_320;
  assign _EVAL_296 = _EVAL_293 | _EVAL_7;
  assign _EVAL_287 = ~_EVAL_296;
  assign _EVAL_24 = _EVAL_73 | _EVAL_273;
  assign _EVAL_243 = _EVAL_228 & _EVAL_295;
  assign _EVAL_274 = _EVAL_1 & _EVAL_300;
  assign _EVAL_209 = ~_EVAL_246;
  assign _EVAL_77 = _EVAL_10[0];
  assign _EVAL_68 = _EVAL_160 | _EVAL_7;
  assign _EVAL_315 = 8'h1 << _EVAL_13;
  assign _EVAL_160 = _EVAL_27 == 4'h0;
  assign _EVAL_60 = ~_EVAL_176;
  assign _EVAL_227 = _EVAL_9 == 3'h4;
  assign _EVAL_297 = {{22'd0}, _EVAL_292};
  assign _EVAL_141 = _EVAL_10[1];
  assign _EVAL_313 = ~_EVAL_141;
  assign _EVAL_125 = _EVAL_3 == 3'h5;
  assign _EVAL_47 = ~_EVAL_208;
  assign _EVAL_153 = _EVAL_290 | _EVAL_7;
  assign _EVAL_126 = ~_EVAL_305;
  assign _EVAL_234 = _EVAL_149 - 6'h1;
  assign _EVAL_215 = _EVAL_6[0];
  assign _EVAL_41 = _EVAL_74 ? _EVAL_315 : 8'h0;
  assign _EVAL_204 = _EVAL_18 == 2'h0;
  assign _EVAL_291 = _EVAL_12 >= 4'h2;
  assign _EVAL_301 = ~_EVAL_77;
  assign _EVAL_247 = _EVAL_195 | _EVAL_7;
  assign _EVAL_208 = _EVAL_82 | _EVAL_7;
  assign _EVAL_280 = _EVAL_12 <= 4'h8;
  assign _EVAL_124 = _EVAL_204 | _EVAL_7;
  assign _EVAL_178 = ~_EVAL_245;
  assign _EVAL_169 = _EVAL_310 != 5'h0;
  assign _EVAL_55 = _EVAL_13 == 3'h4;
  assign _EVAL_123 = ~_EVAL_294;
  assign _EVAL_121 = _EVAL_193;
  assign _EVAL_273 = _EVAL_2 & _EVAL_15;
  assign _EVAL_257 = _EVAL_17 <= 3'h1;
  assign _EVAL_252 = _EVAL_240 | _EVAL_7;
  assign _EVAL_200 = 8'h1 << _EVAL_9;
  assign _EVAL_190 = _EVAL_95 | _EVAL_227;
  assign _EVAL_112 = _EVAL_18 != 2'h2;
  assign _EVAL_107 = ~_EVAL_136;
  assign _EVAL_110 = ~_EVAL_285;
  assign _EVAL_290 = _EVAL_18 == _EVAL_298;
  assign _EVAL_216 = _EVAL_17 == _EVAL_154;
  assign _EVAL_73 = _EVAL & _EVAL_1;
  assign _EVAL_212 = _EVAL_318 | _EVAL_7;
  assign _EVAL_254 = ~_EVAL_252;
  assign _EVAL_222 = _EVAL_291 | _EVAL_54;
  assign _EVAL_197 = ~_EVAL_316;
  assign _EVAL_35 = _EVAL_207 | _EVAL_7;
  assign _EVAL_80 = ~_EVAL_189;
  assign _EVAL_189 = _EVAL_28 | _EVAL_7;
  assign _EVAL_253 = _EVAL_3 == 3'h7;
  assign _EVAL_185 = _EVAL_71 | 2'h1;
  assign _EVAL_39 = _EVAL_1 & _EVAL_63;
  assign _EVAL_327 = _EVAL_280 & _EVAL_113;
  assign _EVAL_84 = _EVAL_122 | _EVAL_92;
  assign _EVAL_142 = _EVAL_1 & _EVAL_60;
  assign _EVAL_25 = _EVAL_10 ^ 30'h2000000;
  assign _EVAL_214 = _EVAL_10 ^ 30'h3000;
  assign _EVAL_96 = _EVAL_277 | _EVAL_7;
  assign _EVAL_61 = _EVAL_141 & _EVAL_301;
  assign _EVAL_260 = _EVAL_97 & _EVAL_87;
  assign _EVAL_67 = _EVAL_202 == 30'h0;
  assign _EVAL_316 = _EVAL_165 | _EVAL_7;
  assign _EVAL_246 = _EVAL_177 | _EVAL_7;
  assign _EVAL_20 = _EVAL_228 & _EVAL_44;
  assign _EVAL_207 = _EVAL_17 != 3'h0;
  assign _EVAL_42 = _EVAL_263 | _EVAL_20;
  assign _EVAL_99 = _EVAL_205 | _EVAL_7;
  assign _EVAL_295 = _EVAL_313 & _EVAL_301;
  assign _EVAL_289 = _EVAL_256 != 5'h0;
  assign _EVAL_206 = _EVAL_327 | _EVAL_260;
  assign _EVAL_305 = _EVAL_291 | _EVAL_7;
  assign _EVAL_255 = _EVAL_12[0];
  assign _EVAL_75 = _EVAL_43 == 6'h0;
  assign _EVAL_86 = ~_EVAL_19;
  assign _EVAL_268 = _EVAL_73 & _EVAL_176;
  assign _EVAL_137 = _EVAL_112 | _EVAL_7;
  assign _EVAL_49 = ~_EVAL_159;
  assign _EVAL_210 = _EVAL_105 | _EVAL_7;
  assign _EVAL_74 = _EVAL_73 & _EVAL_308;
  assign _EVAL_262 = ~_EVAL_7;
  assign _EVAL_303 = _EVAL_311[5:0];
  assign _EVAL_45 = _EVAL_211 | _EVAL_7;
  assign _EVAL_89 = _EVAL_225 | _EVAL_7;
  assign _EVAL_277 = ~_EVAL_5;
  assign _EVAL_120 = _EVAL_180[31:0];
  assign _EVAL_46 = ~_EVAL_233;
  assign _EVAL_272 = ~_EVAL_196;
  assign _EVAL_195 = _EVAL_4 == _EVAL_213;
  assign _EVAL_299 = _EVAL_15 & _EVAL_250;
  assign _EVAL_71 = 2'h1 << _EVAL_255;
  assign _EVAL_168 = ~_EVAL_259;
  assign _EVAL_150 = $signed(_EVAL_114) == 31'sh0;
  assign _EVAL_221 = _EVAL_3 == _EVAL_31;
  assign _EVAL_241 = _EVAL_1 & _EVAL_275;
  assign _EVAL_59 = _EVAL_97 & _EVAL_232;
  assign _EVAL_54 = _EVAL_130 & _EVAL_313;
  assign _EVAL_193 = $signed(_EVAL_187) & -31'sh2000;
  assign _EVAL_162 = _EVAL_248;
  assign _EVAL_56 = ~_EVAL_170;
  assign _EVAL_146 = ~_EVAL_237;
  assign _EVAL_179 = _EVAL_18 <= 2'h2;
  assign _EVAL_33 = _EVAL_6 <= 3'h6;
  assign _EVAL_48 = _EVAL_113 | _EVAL_150;
  assign _EVAL_155 = $signed(_EVAL_53) == 31'sh0;
  assign _EVAL_106 = _EVAL_174 & _EVAL_178;
  assign _EVAL_132 = _EVAL_70 | _EVAL_7;
  assign _EVAL_205 = _EVAL_10 == _EVAL_183;
  assign _EVAL_292 = ~_EVAL_230;
  assign _EVAL_311 = _EVAL_22 - 6'h1;
  assign _EVAL_27 = ~_EVAL_16;
  assign _EVAL_161 = _EVAL_319[7:0];
  assign _EVAL_182 = ~_EVAL_269;
  assign _EVAL_248 = $signed(_EVAL_229) & -31'sh1000;
  assign _EVAL_174 = _EVAL_256 | _EVAL_310;
  assign _EVAL_328 = _EVAL_163 >> _EVAL_9;
  assign _EVAL_36 = ~_EVAL_35;
  assign _EVAL_147 = _EVAL_282[5:0];
  assign _EVAL_105 = _EVAL_17 <= 3'h4;
  assign _EVAL_278 = _EVAL_12 == _EVAL_284;
  assign _EVAL_135 = _EVAL_325 | _EVAL_7;
  assign _EVAL_44 = _EVAL_141 & _EVAL_77;
  assign _EVAL_177 = _EVAL_6 == _EVAL_167;
  assign _EVAL_304 = _EVAL_97 & _EVAL_324;
  assign _EVAL_263 = _EVAL_291 | _EVAL_66;
  assign _EVAL_220 = _EVAL_6 == 3'h2;
  assign _EVAL_131 = ~_EVAL_314;
  assign _EVAL_191 = {1'b0,$signed(_EVAL_10)};
  assign _EVAL_259 = _EVAL_109 | _EVAL_7;
  assign _EVAL_233 = _EVAL_3[2];
  assign _EVAL_228 = _EVAL_185[0];
  assign _EVAL_138 = _EVAL_6 == 3'h5;
  assign _EVAL_165 = _EVAL_11 == _EVAL_139;
  assign _EVAL_62 = _EVAL_263 | _EVAL_235;
  assign _EVAL_156 = ~_EVAL_96;
  assign _EVAL_211 = ~_EVAL_8;
  assign _EVAL_118 = _EVAL_1 & _EVAL_64;
  assign _EVAL_53 = _EVAL_81;
  assign _EVAL_176 = _EVAL_22 == 6'h0;
  assign _EVAL_111 = _EVAL_324 | _EVAL_87;
  assign _EVAL_29 = _EVAL_48 | _EVAL_155;
  assign _EVAL_317 = ~_EVAL_306;
  assign _EVAL_283 = _EVAL_59 | _EVAL_7;
  assign _EVAL_94 = _EVAL_13[2:1];
  assign _EVAL_103 = _EVAL_109 | _EVAL_8;
  assign _EVAL_194 = _EVAL_6 == 3'h6;
  assign _EVAL_151 = _EVAL_327 | _EVAL_304;
  assign _EVAL_225 = ~_EVAL_238;
  assign _EVAL_157 = _EVAL_313 & _EVAL_77;
  assign _EVAL_235 = _EVAL_228 & _EVAL_61;
  assign _EVAL_240 = _EVAL_251 | _EVAL_55;
  assign _EVAL_319 = 23'hff << _EVAL_0;
  assign _EVAL_184 = ~_EVAL_99;
  assign _EVAL_76 = ~_EVAL_89;
  assign _EVAL_37 = ~_EVAL_224;
  assign _EVAL_130 = _EVAL_185[1];
  assign _EVAL_269 = _EVAL_175 | _EVAL_7;
  assign _EVAL_81 = $signed(_EVAL_191) & -31'sh5000;
  assign _EVAL_217 = _EVAL_9[2:1];
  assign _EVAL_285 = _EVAL_84 | _EVAL_7;
  assign _EVAL_282 = _EVAL_264 - 6'h1;
  assign _EVAL_172 = _EVAL_1 & _EVAL_125;
  assign _EVAL_66 = _EVAL_130 & _EVAL_141;
  assign _EVAL_88 = _EVAL_217 == 2'h1;
  assign _EVAL_251 = _EVAL_279 | _EVAL_51;
  assign _EVAL_203 = ~_EVAL_69;
  assign _EVAL_258 = _EVAL_310 != _EVAL_245;
  assign _EVAL_92 = _EVAL_171 < plusarg_reader_out;
  assign _EVAL_230 = _EVAL_133[7:0];
  assign _EVAL_187 = {1'b0,$signed(_EVAL_143)};
  assign _EVAL_152 = _EVAL_288 ? _EVAL_200 : 8'h0;
  assign _EVAL_119 = plusarg_reader_out == 32'h0;
  assign _EVAL_113 = $signed(_EVAL_162) == 31'sh0;
  assign _EVAL_267 = _EVAL_15 & _EVAL_302;
  assign _EVAL_63 = _EVAL_3 == 3'h3;
  assign _EVAL_51 = _EVAL_94 == 2'h0;
  assign _EVAL_133 = 23'hff << _EVAL_12;
  assign _EVAL_250 = _EVAL_6 == 3'h0;
  assign _EVAL_82 = _EVAL_13 == _EVAL_266;
  assign _EVAL_218 = _EVAL_281 | _EVAL_7;
  assign _EVAL_32 = ~_EVAL_58;
  assign _EVAL_100 = ~_EVAL_132;
  assign _EVAL_309 = ~_EVAL_93;
  assign _EVAL_308 = _EVAL_149 == 6'h0;
  assign _EVAL_159 = _EVAL_276 | _EVAL_7;
  assign _EVAL_300 = _EVAL_3 == 3'h4;
  assign _EVAL_102 = _EVAL_273 & _EVAL_170;
  assign _EVAL_116 = _EVAL_17 == 3'h0;
  assign _EVAL_30 = _EVAL_15 & _EVAL_56;
  assign _EVAL_307 = _EVAL_1 & _EVAL_26;
  assign _EVAL_188 = ~_EVAL_135;
  assign _EVAL_148 = ~_EVAL_192;
  assign _EVAL_265 = _EVAL_151 | _EVAL_7;
  assign _EVAL_324 = _EVAL_150 | _EVAL_155;
  assign _EVAL_64 = _EVAL_3 == 3'h6;
  assign _EVAL_232 = _EVAL_29 | _EVAL_87;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_22 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_31 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_43 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_101 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_139 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_149 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_154 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_167 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_171 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_183 = _RAND_9[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_213 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_219 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_256 = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_264 = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_266 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_284 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_298 = _RAND_16[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_14) begin
    if (_EVAL_7) begin
      _EVAL_22 <= 6'h0;
    end else if (_EVAL_73) begin
      if (_EVAL_176) begin
        if (_EVAL_46) begin
          _EVAL_22 <= _EVAL_52;
        end else begin
          _EVAL_22 <= 6'h0;
        end
      end else begin
        _EVAL_22 <= _EVAL_303;
      end
    end
    if (_EVAL_268) begin
      _EVAL_31 <= _EVAL_3;
    end
    if (_EVAL_7) begin
      _EVAL_43 <= 6'h0;
    end else if (_EVAL_273) begin
      if (_EVAL_75) begin
        if (_EVAL_215) begin
          _EVAL_43 <= _EVAL_128;
        end else begin
          _EVAL_43 <= 6'h0;
        end
      end else begin
        _EVAL_43 <= _EVAL_129;
      end
    end
    if (_EVAL_102) begin
      _EVAL_101 <= _EVAL_9;
    end
    if (_EVAL_102) begin
      _EVAL_139 <= _EVAL_11;
    end
    if (_EVAL_7) begin
      _EVAL_149 <= 6'h0;
    end else if (_EVAL_73) begin
      if (_EVAL_308) begin
        if (_EVAL_46) begin
          _EVAL_149 <= _EVAL_52;
        end else begin
          _EVAL_149 <= 6'h0;
        end
      end else begin
        _EVAL_149 <= _EVAL_323;
      end
    end
    if (_EVAL_268) begin
      _EVAL_154 <= _EVAL_17;
    end
    if (_EVAL_102) begin
      _EVAL_167 <= _EVAL_6;
    end
    if (_EVAL_7) begin
      _EVAL_171 <= 32'h0;
    end else if (_EVAL_24) begin
      _EVAL_171 <= 32'h0;
    end else begin
      _EVAL_171 <= _EVAL_120;
    end
    if (_EVAL_268) begin
      _EVAL_183 <= _EVAL_10;
    end
    if (_EVAL_102) begin
      _EVAL_213 <= _EVAL_4;
    end
    if (_EVAL_102) begin
      _EVAL_219 <= _EVAL_0;
    end
    if (_EVAL_7) begin
      _EVAL_256 <= 5'h0;
    end else begin
      _EVAL_256 <= _EVAL_106;
    end
    if (_EVAL_7) begin
      _EVAL_264 <= 6'h0;
    end else if (_EVAL_273) begin
      if (_EVAL_170) begin
        if (_EVAL_215) begin
          _EVAL_264 <= _EVAL_128;
        end else begin
          _EVAL_264 <= 6'h0;
        end
      end else begin
        _EVAL_264 <= _EVAL_147;
      end
    end
    if (_EVAL_268) begin
      _EVAL_266 <= _EVAL_13;
    end
    if (_EVAL_268) begin
      _EVAL_284 <= _EVAL_12;
    end
    if (_EVAL_102) begin
      _EVAL_298 <= _EVAL_18;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11005592)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa1ec43a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3abde3a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dddfc867)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5c490ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6940c86b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a6a7cf8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cf07d04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3fd5d0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(900fca35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(840dc32e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13620057)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(205447f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91e8135c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(766ca263)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6540d3e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27398fe2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8742a04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d55ab57f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbee73ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acd6be12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c30ee17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccf1561b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca7c1036)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(997fd192)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99542aca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1cb998a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f50de34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85b42961)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56818047)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(423fdddb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c8ccfc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c096dfd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(614c2c58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c444832)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fab3db20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8eaf14a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12c23952)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87e983f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(694b3aa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23af42bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcbce7ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86076fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f20b596)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81d432d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3fa20ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3858f8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f77a0b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4843d21a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74ea9711)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd5e1c9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f985fc39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d96f5b73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_287) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fe223f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1971cb10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7cf48d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_309) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7ddbad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_309) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(719ec368)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d31429d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e8999da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4144783a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(428b0ef7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a79ac508)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(655caa4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ae8322f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57bf4dbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c07a360c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd91cd68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(487a0621)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc535e0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ec43300)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f03b136)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed4d2b11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef3e3366)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7bc5bce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16db8ef4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74f24815)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cc28306)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_287) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31668ac4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84ef941b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba1b75e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89b2bbb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5219079a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d63897cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73eeb965)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6e37d56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8cdd93f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a440d73b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13f014c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f5c9cc7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32b4781e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
