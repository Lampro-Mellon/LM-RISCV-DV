//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_163_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [1:0]  _EVAL_4,
  input  [31:0] _EVAL_5,
  input  [3:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [3:0]  _EVAL_12,
  input         _EVAL_13,
  input  [3:0]  _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18
);
  wire [32:0] _EVAL_19;
  wire [1:0] _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire [32:0] _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  reg [3:0] _EVAL_28;
  reg [31:0] _RAND_0;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire [32:0] _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire [32:0] _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire [32:0] _EVAL_55;
  wire [5:0] _EVAL_56;
  wire  _EVAL_57;
  reg [1:0] _EVAL_58;
  reg [31:0] _RAND_1;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  reg  _EVAL_69;
  reg [31:0] _RAND_2;
  wire [1:0] _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire [32:0] _EVAL_74;
  wire [32:0] _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire [31:0] _EVAL_79;
  wire [6:0] _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire [7:0] _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  reg [31:0] _EVAL_90;
  reg [31:0] _RAND_3;
  wire [32:0] _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  reg [3:0] _EVAL_94;
  reg [31:0] _RAND_4;
  wire  _EVAL_96;
  wire [31:0] _EVAL_97;
  wire [31:0] _EVAL_98;
  wire  _EVAL_99;
  wire [31:0] plusarg_reader_out;
  wire [32:0] _EVAL_100;
  wire [6:0] _EVAL_101;
  wire [1:0] _EVAL_102;
  wire [32:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_114;
  wire  _EVAL_116;
  reg [5:0] _EVAL_118;
  reg [31:0] _RAND_5;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  reg [1:0] _EVAL_123;
  reg [31:0] _RAND_6;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire [32:0] _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire [6:0] _EVAL_133;
  wire  _EVAL_134;
  reg  _EVAL_135;
  reg [31:0] _RAND_7;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire [32:0] _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire [1:0] _EVAL_148;
  wire [3:0] _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire [5:0] _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire [5:0] _EVAL_172;
  wire [22:0] _EVAL_173;
  wire  _EVAL_174;
  wire [1:0] _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire [31:0] _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  reg  _EVAL_186;
  reg [31:0] _RAND_8;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire [1:0] _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  reg [2:0] _EVAL_203;
  reg [31:0] _RAND_9;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  reg [5:0] _EVAL_210;
  reg [31:0] _RAND_10;
  wire [32:0] _EVAL_211;
  wire [7:0] _EVAL_212;
  wire  _EVAL_213;
  reg [5:0] _EVAL_214;
  reg [31:0] _RAND_11;
  wire [32:0] _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  reg  _EVAL_228;
  reg [31:0] _RAND_12;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire [3:0] _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire [1:0] _EVAL_234;
  wire  _EVAL_235;
  wire [1:0] _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire [31:0] _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  reg [2:0] _EVAL_243;
  reg [31:0] _RAND_13;
  wire  _EVAL_244;
  wire [5:0] _EVAL_245;
  wire [31:0] _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire [32:0] _EVAL_250;
  reg [5:0] _EVAL_251;
  reg [31:0] _RAND_14;
  wire [31:0] _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_257;
  wire [5:0] _EVAL_258;
  wire  _EVAL_259;
  wire [1:0] _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire [7:0] _EVAL_269;
  wire [6:0] _EVAL_270;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire [3:0] _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire [31:0] _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire [5:0] _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  reg [2:0] _EVAL_287;
  reg [31:0] _RAND_15;
  wire  _EVAL_288;
  wire [1:0] _EVAL_289;
  wire [1:0] _EVAL_290;
  wire [7:0] _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  reg [31:0] _EVAL_295;
  reg [31:0] _RAND_16;
  wire [32:0] _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_299;
  wire [32:0] _EVAL_300;
  wire [32:0] _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire [3:0] _EVAL_309;
  wire [1:0] _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire [22:0] _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire  _EVAL_318;
  wire [32:0] _EVAL_319;
  wire  _EVAL_320;
  wire  _EVAL_322;
  wire  _EVAL_323;
  wire  _EVAL_324;
  wire  _EVAL_325;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_241 = _EVAL_3 == 3'h0;
  assign _EVAL_78 = _EVAL_2 == 3'h2;
  assign _EVAL_183 = _EVAL_240 | _EVAL_11;
  assign _EVAL_97 = _EVAL_5 ^ 32'h3000;
  assign _EVAL_35 = _EVAL_14[0];
  assign _EVAL_250 = _EVAL_75;
  assign _EVAL_188 = _EVAL_288 | _EVAL_156;
  assign _EVAL_134 = _EVAL_9 == _EVAL_228;
  assign _EVAL_264 = _EVAL_109 | _EVAL_11;
  assign _EVAL_209 = _EVAL_17 == _EVAL_186;
  assign _EVAL_249 = ~_EVAL_27;
  assign _EVAL_285 = _EVAL_210 == 6'h0;
  assign _EVAL_279 = _EVAL_100[31:0];
  assign _EVAL_86 = _EVAL_8 & _EVAL_83;
  assign _EVAL_275 = {_EVAL_76,_EVAL_201,_EVAL_194,_EVAL_62};
  assign _EVAL_175 = _EVAL_70 >> _EVAL_9;
  assign _EVAL_231 = ~_EVAL_12;
  assign _EVAL_263 = ~_EVAL_224;
  assign _EVAL_236 = 2'h1 << _EVAL_35;
  assign _EVAL_223 = _EVAL_105 | _EVAL_142;
  assign _EVAL_244 = _EVAL_179 | _EVAL_325;
  assign _EVAL_281 = _EVAL & _EVAL_8;
  assign _EVAL_142 = _EVAL_112 & _EVAL_38;
  assign _EVAL_45 = _EVAL_84 | _EVAL_11;
  assign _EVAL_198 = _EVAL_281 & _EVAL_293;
  assign _EVAL_288 = _EVAL_14 >= 4'h2;
  assign _EVAL_82 = _EVAL_1 & _EVAL_48;
  assign _EVAL_36 = ~_EVAL_72;
  assign _EVAL_258 = _EVAL_270[5:0];
  assign _EVAL_242 = _EVAL_15 <= 3'h4;
  assign _EVAL_127 = _EVAL_1 & _EVAL_299;
  assign _EVAL_229 = ~_EVAL_204;
  assign _EVAL_206 = _EVAL_4 == 2'h0;
  assign _EVAL_213 = _EVAL_4 <= 2'h2;
  assign _EVAL_110 = _EVAL_134 | _EVAL_11;
  assign _EVAL_71 = ~_EVAL_99;
  assign _EVAL_139 = _EVAL_118 == 6'h0;
  assign _EVAL_184 = ~_EVAL_126;
  assign _EVAL_144 = _EVAL_3 == 3'h1;
  assign _EVAL_306 = ~_EVAL_16;
  assign _EVAL_168 = _EVAL_5[1];
  assign _EVAL_212 = ~_EVAL_291;
  assign _EVAL_181 = plusarg_reader_out == 32'h0;
  assign _EVAL_283 = _EVAL_101[5:0];
  assign _EVAL_51 = _EVAL_15 <= 3'h3;
  assign _EVAL_107 = _EVAL_3 == 3'h2;
  assign _EVAL_297 = $signed(_EVAL_25) == 33'sh0;
  assign _EVAL_141 = ~_EVAL_168;
  assign _EVAL_240 = _EVAL_15 == 3'h0;
  assign _EVAL_255 = _EVAL_15 != 3'h0;
  assign _EVAL_316 = _EVAL_51 | _EVAL_11;
  assign _EVAL_146 = ~_EVAL_262;
  assign _EVAL_171 = ~_EVAL_47;
  assign _EVAL_33 = ~_EVAL_268;
  assign _EVAL_220 = _EVAL_3[2];
  assign _EVAL_25 = _EVAL_44;
  assign _EVAL_130 = _EVAL_251 == 6'h0;
  assign _EVAL_178 = _EVAL_5 & _EVAL_98;
  assign _EVAL_132 = _EVAL_1 & _EVAL_78;
  assign _EVAL_309 = ~_EVAL_275;
  assign _EVAL_34 = _EVAL_301;
  assign _EVAL_89 = _EVAL_59 | _EVAL_16;
  assign _EVAL_311 = _EVAL_116 | _EVAL_11;
  assign _EVAL_315 = _EVAL_180 | _EVAL_11;
  assign _EVAL_67 = _EVAL_278 | _EVAL_11;
  assign _EVAL_77 = ~_EVAL_159;
  assign _EVAL_121 = ~_EVAL_124;
  assign _EVAL_138 = _EVAL_310[0];
  assign _EVAL_197 = _EVAL_43 | _EVAL_145;
  assign _EVAL_29 = ~_EVAL_130;
  assign _EVAL_267 = ~_EVAL_324;
  assign _EVAL_152 = _EVAL_138 & _EVAL_266;
  assign _EVAL_119 = _EVAL_59 | _EVAL_11;
  assign _EVAL_176 = ~_EVAL_41;
  assign _EVAL_59 = ~_EVAL_13;
  assign _EVAL_52 = _EVAL_5 == _EVAL_295;
  assign _EVAL_191 = _EVAL_15 == _EVAL_287;
  assign _EVAL_312 = _EVAL_102 != 2'h0;
  assign _EVAL_219 = ~_EVAL_316;
  assign _EVAL_47 = _EVAL_255 | _EVAL_11;
  assign _EVAL_204 = _EVAL_123 != 2'h0;
  assign _EVAL_266 = _EVAL_168 & _EVAL_131;
  assign _EVAL_96 = _EVAL_2 == 3'h6;
  assign _EVAL_46 = _EVAL_3 == 3'h6;
  assign _EVAL_79 = _EVAL_5 ^ 32'h80000000;
  assign _EVAL_38 = $signed(_EVAL_250) == 33'sh0;
  assign _EVAL_208 = _EVAL_102 != _EVAL_234;
  assign _EVAL_238 = _EVAL_196 & _EVAL_197;
  assign _EVAL_325 = _EVAL_90 < plusarg_reader_out;
  assign _EVAL_20 = _EVAL_123 >> _EVAL_17;
  assign _EVAL_154 = ~_EVAL_170;
  assign _EVAL_274 = _EVAL_288 | _EVAL_318;
  assign _EVAL_172 = _EVAL_80[5:0];
  assign _EVAL_153 = _EVAL_294 & _EVAL_182;
  assign _EVAL_91 = $signed(_EVAL_300) & -33'sh1000000;
  assign _EVAL_114 = ~_EVAL_202;
  assign _EVAL_310 = _EVAL_236 | 2'h1;
  assign _EVAL_98 = {{24'd0}, _EVAL_87};
  assign _EVAL_49 = $signed(_EVAL_34) == 33'sh0;
  assign _EVAL_122 = _EVAL_0 & _EVAL_1;
  assign _EVAL_300 = {1'b0,$signed(_EVAL_239)};
  assign _EVAL_124 = _EVAL_288 | _EVAL_11;
  assign _EVAL_221 = ~_EVAL_160;
  assign _EVAL_276 = ~_EVAL_259;
  assign _EVAL_100 = _EVAL_90 + 32'h1;
  assign _EVAL_260 = 2'h1 << _EVAL_9;
  assign _EVAL_161 = _EVAL_8 & _EVAL_57;
  assign _EVAL_239 = _EVAL_5 ^ 32'h2000000;
  assign _EVAL_145 = $signed(_EVAL_103) == 33'sh0;
  assign _EVAL_87 = ~_EVAL_269;
  assign _EVAL_270 = _EVAL_251 - 6'h1;
  assign _EVAL_226 = _EVAL_8 & _EVAL_241;
  assign _EVAL_247 = _EVAL_197 | _EVAL_297;
  assign _EVAL_245 = _EVAL_212[7:2];
  assign _EVAL_173 = 23'hff << _EVAL_6;
  assign _EVAL_31 = ~_EVAL_285;
  assign _EVAL_272 = _EVAL_169 | _EVAL_11;
  assign _EVAL_324 = _EVAL_261 | _EVAL_11;
  assign _EVAL_24 = _EVAL_3 == 3'h7;
  assign _EVAL_55 = {1'b0,$signed(_EVAL_79)};
  assign _EVAL_125 = _EVAL_8 & _EVAL_24;
  assign _EVAL_313 = _EVAL_138 & _EVAL_167;
  assign _EVAL_136 = _EVAL_2 <= 3'h6;
  assign _EVAL_56 = _EVAL_133[5:0];
  assign _EVAL_268 = _EVAL_52 | _EVAL_11;
  assign _EVAL_26 = _EVAL_22 | _EVAL_11;
  assign _EVAL_167 = _EVAL_168 & _EVAL_302;
  assign _EVAL_169 = _EVAL_3 == _EVAL_243;
  assign _EVAL_140 = {1'b0,$signed(_EVAL_97)};
  assign _EVAL_296 = {1'b0,$signed(_EVAL_253)};
  assign _EVAL_44 = $signed(_EVAL_296) & -33'sh2000;
  assign _EVAL_222 = $signed(_EVAL_211) == 33'sh0;
  assign _EVAL_160 = _EVAL_273 | _EVAL_11;
  assign _EVAL_174 = ~_EVAL_11;
  assign _EVAL_180 = _EVAL_231 == 4'h0;
  assign _EVAL_126 = _EVAL_223 | _EVAL_11;
  assign _EVAL_194 = _EVAL_188 | _EVAL_323;
  assign _EVAL_207 = ~_EVAL_110;
  assign _EVAL_215 = _EVAL_19;
  assign _EVAL_104 = ~_EVAL_73;
  assign _EVAL_305 = _EVAL_281 & _EVAL_130;
  assign _EVAL_158 = _EVAL_87[7:2];
  assign _EVAL_62 = _EVAL_188 | _EVAL_166;
  assign _EVAL_224 = _EVAL_65 | _EVAL_11;
  assign _EVAL_131 = _EVAL_5[0];
  assign _EVAL_277 = _EVAL_2 == 3'h4;
  assign _EVAL_217 = _EVAL_306 | _EVAL_11;
  assign _EVAL_234 = _EVAL_92 ? _EVAL_260 : 2'h0;
  assign _EVAL_262 = _EVAL_189 | _EVAL_11;
  assign _EVAL_233 = _EVAL_282 | _EVAL_11;
  assign _EVAL_273 = _EVAL_12 == _EVAL_275;
  assign _EVAL_68 = _EVAL_196 & _EVAL_247;
  assign _EVAL_74 = {1'b0,$signed(_EVAL_5)};
  assign _EVAL_63 = _EVAL_15 <= 3'h1;
  assign _EVAL_66 = _EVAL_196 & _EVAL_297;
  assign _EVAL_314 = 23'hff << _EVAL_14;
  assign _EVAL_42 = ~_EVAL_187;
  assign _EVAL_254 = _EVAL_310[1];
  assign _EVAL_261 = _EVAL_178 == 32'h0;
  assign _EVAL_137 = ~_EVAL_45;
  assign _EVAL_85 = _EVAL_238 | _EVAL_142;
  assign _EVAL_202 = _EVAL_242 | _EVAL_11;
  assign _EVAL_292 = _EVAL_136 | _EVAL_11;
  assign _EVAL_103 = _EVAL_319;
  assign _EVAL_227 = _EVAL_4 != 2'h2;
  assign _EVAL_147 = _EVAL_175[0];
  assign _EVAL_88 = _EVAL_303 | _EVAL_66;
  assign _EVAL_216 = _EVAL_281 | _EVAL_122;
  assign _EVAL_170 = _EVAL_147 | _EVAL_11;
  assign _EVAL_269 = _EVAL_314[7:0];
  assign _EVAL_101 = _EVAL_210 - 6'h1;
  assign _EVAL_317 = ~_EVAL_220;
  assign _EVAL_189 = _EVAL_6 == _EVAL_28;
  assign _EVAL_156 = _EVAL_254 & _EVAL_141;
  assign _EVAL_282 = ~_EVAL_320;
  assign _EVAL_319 = $signed(_EVAL_74) & -33'sh5000;
  assign _EVAL_303 = _EVAL_153 | _EVAL_142;
  assign _EVAL_143 = ~_EVAL_286;
  assign _EVAL_187 = _EVAL_206 | _EVAL_11;
  assign _EVAL_108 = ~_EVAL_96;
  assign _EVAL_22 = _EVAL_14 == _EVAL_94;
  assign _EVAL_166 = _EVAL_138 & _EVAL_265;
  assign _EVAL_257 = ~_EVAL_26;
  assign _EVAL_308 = ~_EVAL_304;
  assign _EVAL_211 = _EVAL_91;
  assign _EVAL_133 = _EVAL_118 - 6'h1;
  assign _EVAL_301 = $signed(_EVAL_55) & -33'shc000;
  assign _EVAL_177 = _EVAL_199 | _EVAL_11;
  assign _EVAL_290 = 2'h1 << _EVAL_17;
  assign _EVAL_265 = _EVAL_141 & _EVAL_302;
  assign _EVAL_294 = _EVAL_14 <= 4'h6;
  assign _EVAL_190 = _EVAL_225 | _EVAL_11;
  assign _EVAL_109 = _EVAL_15 <= 3'h2;
  assign _EVAL_112 = _EVAL_14 <= 4'h8;
  assign _EVAL_280 = _EVAL_1 & _EVAL_185;
  assign _EVAL_155 = _EVAL_122 & _EVAL_285;
  assign _EVAL_70 = _EVAL_102 | _EVAL_123;
  assign _EVAL_57 = _EVAL_3 == 3'h3;
  assign _EVAL_32 = _EVAL_38 | _EVAL_222;
  assign _EVAL_200 = ~_EVAL_234;
  assign _EVAL_116 = _EVAL_149 == 4'h0;
  assign _EVAL_27 = _EVAL_227 | _EVAL_11;
  assign _EVAL_75 = $signed(_EVAL_140) & -33'sh1000;
  assign _EVAL_259 = _EVAL_88 | _EVAL_11;
  assign _EVAL_302 = ~_EVAL_131;
  assign _EVAL_293 = _EVAL_214 == 6'h0;
  assign _EVAL_157 = _EVAL_37 | _EVAL_297;
  assign _EVAL_149 = _EVAL_12 & _EVAL_309;
  assign _EVAL_299 = _EVAL_2 == 3'h5;
  assign _EVAL_72 = _EVAL_63 | _EVAL_11;
  assign _EVAL_225 = _EVAL_208 | _EVAL_284;
  assign _EVAL_54 = _EVAL_3 == 3'h4;
  assign _EVAL_39 = _EVAL_53 | _EVAL_11;
  assign _EVAL_235 = ~_EVAL_233;
  assign _EVAL_148 = _EVAL_123 | _EVAL_102;
  assign _EVAL_304 = _EVAL_244 | _EVAL_11;
  assign _EVAL_76 = _EVAL_274 | _EVAL_152;
  assign _EVAL_83 = _EVAL_3 == 3'h5;
  assign _EVAL_195 = _EVAL_2[0];
  assign _EVAL_205 = ~_EVAL_272;
  assign _EVAL_237 = _EVAL_8 & _EVAL_144;
  assign _EVAL_53 = _EVAL_2 == _EVAL_203;
  assign _EVAL_201 = _EVAL_274 | _EVAL_313;
  assign _EVAL_65 = ~_EVAL_10;
  assign _EVAL_199 = _EVAL_7 == _EVAL_135;
  assign _EVAL_60 = ~_EVAL_190;
  assign _EVAL_84 = _EVAL_13 == _EVAL_69;
  assign _EVAL_278 = _EVAL_6 >= 4'h2;
  assign _EVAL_322 = _EVAL_4 == _EVAL_58;
  assign _EVAL_128 = {1'b0,$signed(_EVAL_246)};
  assign _EVAL_48 = _EVAL_2 == 3'h1;
  assign _EVAL_318 = _EVAL_254 & _EVAL_168;
  assign _EVAL_164 = _EVAL_141 & _EVAL_131;
  assign _EVAL_40 = _EVAL_8 & _EVAL_54;
  assign _EVAL_41 = _EVAL_213 | _EVAL_11;
  assign _EVAL_150 = ~_EVAL_183;
  assign _EVAL_21 = _EVAL_1 & _EVAL_96;
  assign _EVAL_92 = _EVAL_192 & _EVAL_108;
  assign _EVAL_185 = _EVAL_2 == 3'h0;
  assign _EVAL_106 = ~_EVAL_315;
  assign _EVAL_102 = _EVAL_198 ? _EVAL_290 : 2'h0;
  assign _EVAL_182 = $signed(_EVAL_215) == 33'sh0;
  assign _EVAL_323 = _EVAL_138 & _EVAL_164;
  assign _EVAL_111 = ~_EVAL_217;
  assign _EVAL_179 = _EVAL_229 | _EVAL_181;
  assign _EVAL_232 = ~_EVAL_50;
  assign _EVAL_165 = _EVAL_196 & _EVAL_157;
  assign _EVAL_246 = _EVAL_5 ^ 32'h40000000;
  assign _EVAL_192 = _EVAL_122 & _EVAL_139;
  assign _EVAL_23 = ~_EVAL_30;
  assign _EVAL_151 = ~_EVAL_119;
  assign _EVAL_159 = _EVAL_209 | _EVAL_11;
  assign _EVAL_291 = _EVAL_173[7:0];
  assign _EVAL_193 = _EVAL_8 & _EVAL_46;
  assign _EVAL_129 = _EVAL_1 & _EVAL_31;
  assign _EVAL_37 = _EVAL_32 | _EVAL_145;
  assign _EVAL_253 = _EVAL_5 ^ 32'h20000000;
  assign _EVAL_230 = ~_EVAL_292;
  assign _EVAL_289 = _EVAL_148 & _EVAL_200;
  assign _EVAL_80 = _EVAL_214 - 6'h1;
  assign _EVAL_50 = _EVAL_322 | _EVAL_11;
  assign _EVAL_73 = _EVAL_85 | _EVAL_11;
  assign _EVAL_105 = _EVAL_68 | _EVAL_153;
  assign _EVAL_19 = $signed(_EVAL_128) & -33'sh2000;
  assign _EVAL_248 = ~_EVAL_39;
  assign _EVAL_320 = _EVAL_20[0];
  assign _EVAL_43 = _EVAL_49 | _EVAL_222;
  assign _EVAL_120 = ~_EVAL_264;
  assign _EVAL_284 = ~_EVAL_312;
  assign _EVAL_93 = _EVAL_8 & _EVAL_29;
  assign _EVAL_307 = ~_EVAL_311;
  assign _EVAL_64 = _EVAL_1 & _EVAL_277;
  assign _EVAL_81 = _EVAL_8 & _EVAL_107;
  assign _EVAL_196 = _EVAL_14 <= 4'h2;
  assign _EVAL_163 = ~_EVAL_177;
  assign _EVAL_99 = _EVAL_191 | _EVAL_11;
  assign _EVAL_30 = _EVAL_165 | _EVAL_11;
  assign _EVAL_286 = _EVAL_89 | _EVAL_11;
  assign _EVAL_218 = ~_EVAL_67;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_28 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_58 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_69 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_90 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_94 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_118 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_123 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_135 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_186 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_203 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_210 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_214 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_228 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_243 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_251 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_287 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_295 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_18) begin
    if (_EVAL_155) begin
      _EVAL_28 <= _EVAL_6;
    end
    if (_EVAL_155) begin
      _EVAL_58 <= _EVAL_4;
    end
    if (_EVAL_155) begin
      _EVAL_69 <= _EVAL_13;
    end
    if (_EVAL_11) begin
      _EVAL_90 <= 32'h0;
    end else if (_EVAL_216) begin
      _EVAL_90 <= 32'h0;
    end else begin
      _EVAL_90 <= _EVAL_279;
    end
    if (_EVAL_305) begin
      _EVAL_94 <= _EVAL_14;
    end
    if (_EVAL_11) begin
      _EVAL_118 <= 6'h0;
    end else if (_EVAL_122) begin
      if (_EVAL_139) begin
        if (_EVAL_195) begin
          _EVAL_118 <= _EVAL_245;
        end else begin
          _EVAL_118 <= 6'h0;
        end
      end else begin
        _EVAL_118 <= _EVAL_56;
      end
    end
    if (_EVAL_11) begin
      _EVAL_123 <= 2'h0;
    end else begin
      _EVAL_123 <= _EVAL_289;
    end
    if (_EVAL_155) begin
      _EVAL_135 <= _EVAL_7;
    end
    if (_EVAL_305) begin
      _EVAL_186 <= _EVAL_17;
    end
    if (_EVAL_155) begin
      _EVAL_203 <= _EVAL_2;
    end
    if (_EVAL_11) begin
      _EVAL_210 <= 6'h0;
    end else if (_EVAL_122) begin
      if (_EVAL_285) begin
        if (_EVAL_195) begin
          _EVAL_210 <= _EVAL_245;
        end else begin
          _EVAL_210 <= 6'h0;
        end
      end else begin
        _EVAL_210 <= _EVAL_283;
      end
    end
    if (_EVAL_11) begin
      _EVAL_214 <= 6'h0;
    end else if (_EVAL_281) begin
      if (_EVAL_293) begin
        if (_EVAL_317) begin
          _EVAL_214 <= _EVAL_158;
        end else begin
          _EVAL_214 <= 6'h0;
        end
      end else begin
        _EVAL_214 <= _EVAL_172;
      end
    end
    if (_EVAL_155) begin
      _EVAL_228 <= _EVAL_9;
    end
    if (_EVAL_305) begin
      _EVAL_243 <= _EVAL_3;
    end
    if (_EVAL_11) begin
      _EVAL_251 <= 6'h0;
    end else if (_EVAL_281) begin
      if (_EVAL_130) begin
        if (_EVAL_317) begin
          _EVAL_251 <= _EVAL_158;
        end else begin
          _EVAL_251 <= 6'h0;
        end
      end else begin
        _EVAL_251 <= _EVAL_258;
      end
    end
    if (_EVAL_305) begin
      _EVAL_287 <= _EVAL_15;
    end
    if (_EVAL_305) begin
      _EVAL_295 <= _EVAL_5;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbd1de7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3879979d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69219bab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a1f8a09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fea92950)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(673a8de7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(994e5ee3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cab0925e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9baf7eea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0471b4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a57d90a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35d36280)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cef455b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13ddba57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d638ea3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6c5457e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_308) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c25ab55d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e1ab22b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a5d0f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e205a12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f55fa41c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d82f152)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(558d7513)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(485056c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1602382)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec6dbcac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34b9f105)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_307) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bff8b648)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c58e501e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffdd95a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6eb91f67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_307) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_308) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(744627c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c22f48fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8793b5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a16350da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffcd9843)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c382d4e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3af52e82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42741129)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(206d14d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4aebeeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b3b9cc4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b86b16f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f12255b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae9b751a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7047f3fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdd0dddb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebc31213)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(310abcd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5379f74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79af1693)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(249ed36b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(634bc176)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad625f62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4313905)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d08a293)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6e52b22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4ffac33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b52eeb42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4554fd86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d32e7053)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70d33460)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(923737d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9af49a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6329dd2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(830e4bc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ceeb6029)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46d571f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a57d2f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45b949ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d31ef4bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f620f4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d287d6ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44ba9f37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a90f547)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79527ee9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be47aba3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
