//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_158(
  input         _EVAL,
  output        _EVAL_0,
  input  [7:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  output        _EVAL_3,
  output        _EVAL_4,
  output        _EVAL_5,
  output [31:0] _EVAL_6,
  input  [3:0]  _EVAL_7,
  input         _EVAL_8,
  output [2:0]  _EVAL_9,
  output        _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [7:0]  _EVAL_14,
  output        _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  output        _EVAL_18,
  output [3:0]  _EVAL_19,
  input         _EVAL_20,
  output [31:0] _EVAL_21,
  output        _EVAL_22,
  input         _EVAL_23,
  output        _EVAL_24,
  input  [1:0]  _EVAL_25,
  output [2:0]  _EVAL_26,
  output [2:0]  _EVAL_27,
  output        _EVAL_28,
  input         _EVAL_29,
  output        _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  output        _EVAL_33,
  output        _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36,
  output        _EVAL_37,
  output        _EVAL_38,
  output        _EVAL_39,
  input         _EVAL_40,
  output        _EVAL_41,
  output        _EVAL_42,
  output        _EVAL_43,
  output        _EVAL_44,
  output [31:0] _EVAL_45,
  output        _EVAL_46,
  input         _EVAL_47,
  input  [3:0]  _EVAL_48,
  output [2:0]  _EVAL_49,
  output        _EVAL_50,
  input  [31:0] _EVAL_51,
  output        _EVAL_52,
  input  [31:0] _EVAL_53,
  output        _EVAL_54,
  input         _EVAL_55,
  output [31:0] _EVAL_56,
  input         _EVAL_57,
  output [3:0]  _EVAL_58,
  output [3:0]  _EVAL_59,
  input  [31:0] _EVAL_60,
  input  [1:0]  _EVAL_61,
  output [3:0]  _EVAL_62,
  output        _EVAL_63,
  input         _EVAL_64,
  output        _EVAL_65,
  output        _EVAL_66,
  input         _EVAL_67,
  input  [2:0]  _EVAL_68
);
  wire [2:0] _EVAL_92;
  wire [32:0] _EVAL_98;
  wire [2:0] _EVAL_127;
  wire [2:0] _EVAL_151;
  wire  _EVAL_221;
  wire [31:0] _EVAL_236;
  wire  _EVAL_241;
  wire [31:0] _EVAL_272;
  wire  _EVAL_284;
  wire  _EVAL_319;
  wire  _EVAL_403;
  wire  _EVAL_409;
  wire  _EVAL_413;
  wire [3:0] _EVAL_423;
  wire [32:0] _EVAL_427;
  wire [9:0] _EVAL_434;
  wire  _EVAL_437;
  wire  _EVAL_464;
  wire  _EVAL_477;
  wire  _EVAL_500;
  wire  _EVAL_528;
  wire [1:0] _EVAL_551;
  wire  _EVAL_573;
  wire  _EVAL_586;
  wire  _EVAL_588;
  wire  _EVAL_636;
  wire  _EVAL_637;
  wire  _EVAL_639;
  wire [31:0] _EVAL_641;
  wire [31:0] _EVAL_642;
  wire  _EVAL_703;
  wire  _EVAL_706;
  wire [31:0] _EVAL_779;
  wire [31:0] _EVAL_805;
  wire  _EVAL_814;
  wire  _EVAL_840;
  wire  _EVAL_849;
  wire [2:0] _EVAL_857;
  wire  _EVAL_869;
  wire  _EVAL_874;
  wire [31:0] _EVAL_880;
  wire  _EVAL_884;
  wire  _EVAL_897;
  wire  _EVAL_909;
  wire  _EVAL_919;
  wire  _EVAL_935;
  wire  _EVAL_948;
  wire  _EVAL_952;
  wire  _EVAL_968;
  wire  _EVAL_974;
  wire  _EVAL_982;
  wire [31:0] _EVAL_1027;
  wire  _EVAL_1067;
  wire  _EVAL_1087;
  wire [4:0] _EVAL_1128;
  wire  fetch_pmp_checker__EVAL;
  wire  fetch_pmp_checker__EVAL_0;
  wire [31:0] fetch_pmp_checker__EVAL_1;
  wire [1:0] fetch_pmp_checker__EVAL_2;
  wire  fetch_pmp_checker__EVAL_3;
  wire  fetch_pmp_checker__EVAL_4;
  wire  fetch_pmp_checker__EVAL_5;
  wire  fetch_pmp_checker__EVAL_6;
  wire  fetch_pmp_checker__EVAL_7;
  wire  fetch_pmp_checker__EVAL_8;
  wire  fetch_pmp_checker__EVAL_9;
  wire [29:0] fetch_pmp_checker__EVAL_10;
  wire [1:0] fetch_pmp_checker__EVAL_11;
  wire [31:0] fetch_pmp_checker__EVAL_12;
  wire  fetch_pmp_checker__EVAL_13;
  wire [29:0] fetch_pmp_checker__EVAL_14;
  wire  fetch_pmp_checker__EVAL_15;
  wire  fetch_pmp_checker__EVAL_16;
  wire [29:0] fetch_pmp_checker__EVAL_17;
  wire  fetch_pmp_checker__EVAL_18;
  wire [31:0] fetch_pmp_checker__EVAL_19;
  wire [1:0] fetch_pmp_checker__EVAL_20;
  wire  fetch_pmp_checker__EVAL_21;
  wire  fetch_pmp_checker__EVAL_22;
  wire [1:0] fetch_pmp_checker__EVAL_23;
  wire  fetch_pmp_checker__EVAL_24;
  wire [29:0] fetch_pmp_checker__EVAL_25;
  wire [31:0] fetch_pmp_checker__EVAL_26;
  wire  fetch_pmp_checker__EVAL_27;
  wire  fetch_pmp_checker__EVAL_28;
  wire  fetch_pmp_checker__EVAL_29;
  wire [1:0] fetch_pmp_checker__EVAL_30;
  wire  fetch_pmp_checker__EVAL_31;
  wire [31:0] fetch_pmp_checker__EVAL_32;
  wire  fetch_pmp_checker__EVAL_33;
  wire [32:0] _EVAL_1185;
  wire  _EVAL_1267;
  wire  _EVAL_1297;
  wire [31:0] _EVAL_1311;
  wire  _EVAL_1324;
  wire  _EVAL_1336;
  wire  _EVAL_1372;
  wire  _EVAL_1385;
  wire  _EVAL_1389;
  wire  _EVAL_1397;
  wire  _EVAL_1404;
  wire  _EVAL_1437;
  wire [4:0] _EVAL_1451;
  wire  _EVAL_1478;
  wire [3:0] _EVAL_1503;
  wire [31:0] _EVAL_1530;
  wire  _EVAL_1546;
  wire [31:0] _EVAL_1606;
  wire  _EVAL_1627;
  wire  _EVAL_1636;
  wire  _EVAL_1638;
  wire  _EVAL_1640;
  wire  _EVAL_1738;
  wire  _EVAL_1739;
  wire [1:0] _EVAL_1745;
  wire  _EVAL_1801;
  wire [23:0] _EVAL_1811;
  wire  _EVAL_1860;
  wire [33:0] _EVAL_1888;
  wire  _EVAL_1962;
  wire  _EVAL_1969;
  wire  _EVAL_1983;
  wire [31:0] _EVAL_1988;
  wire  _EVAL_1995;
  wire  _EVAL_2021;
  wire  _EVAL_2058;
  wire  _EVAL_2080;
  wire  _EVAL_2084;
  wire [31:0] _EVAL_2086;
  reg [3:0] _EVAL_2097;
  reg [31:0] _RAND_0;
  wire [23:0] _EVAL_2100;
  wire  _EVAL_2109;
  wire [31:0] _EVAL_2113;
  wire  _EVAL_2125;
  wire  _EVAL_2139;
  wire  _EVAL_2198;
  reg [2:0] _EVAL_2215;
  reg [31:0] _RAND_1;
  wire  _EVAL_2225;
  wire  _EVAL_2238;
  wire  _EVAL_2258;
  wire [2:0] _EVAL_2265;
  wire  _EVAL_2277;
  wire  _EVAL_2293;
  wire  _EVAL_2322;
  wire  _EVAL_2373;
  wire  _EVAL_2446;
  wire  _EVAL_2447;
  wire  _EVAL_2458;
  wire  _EVAL_2483;
  wire  _EVAL_2488;
  wire  _EVAL_2492;
  wire  _EVAL_2508;
  wire  _EVAL_2558;
  wire  _EVAL_2593;
  wire [2:0] _EVAL_2604;
  wire  _EVAL_2629;
  wire  _EVAL_2638;
  wire  _EVAL_2644;
  wire [1:0] _EVAL_2653;
  wire  _EVAL_2654;
  reg [1:0] _EVAL_2667;
  reg [31:0] _RAND_2;
  wire [31:0] _EVAL_2703;
  wire [31:0] _EVAL_2706;
  wire [32:0] _EVAL_2727;
  wire [31:0] _EVAL_2740;
  wire  _EVAL_2743;
  reg [4:0] _EVAL_2751;
  reg [31:0] _RAND_3;
  wire  _EVAL_2761;
  wire  _EVAL_2764;
  wire [31:0] _EVAL_2793;
  wire [31:0] _EVAL_2832;
  wire  _EVAL_2835;
  wire [31:0] _EVAL_2845;
  wire  _EVAL_2871;
  wire  _EVAL_2872;
  wire  _EVAL_2895;
  wire [1:0] _EVAL_2900;
  wire [32:0] _EVAL_2941;
  wire  _EVAL_2945;
  wire  _EVAL_2953;
  wire [31:0] _EVAL_3045;
  reg [31:0] _EVAL_3051;
  reg [31:0] _RAND_4;
  wire [31:0] _EVAL_3102;
  wire [2:0] _EVAL_3104;
  wire  _EVAL_3117;
  wire  _EVAL_3121;
  reg  _EVAL_3130;
  reg [31:0] _RAND_5;
  wire  _EVAL_3139;
  wire  _EVAL_3157;
  wire  _EVAL_3170;
  wire  _EVAL_3248;
  wire [2:0] _EVAL_3302;
  wire  _EVAL_3320;
  wire [31:0] _EVAL_3322;
  wire [31:0] _EVAL_3330;
  wire  _EVAL_3352;
  wire  _EVAL_3442;
  wire  _EVAL_3444;
  wire  _EVAL_3448;
  wire  _EVAL_3491;
  wire  _EVAL_3495;
  wire  _EVAL_3497;
  wire  _EVAL_3500;
  wire [32:0] _EVAL_3544;
  wire  _EVAL_3556;
  wire  _EVAL_3585;
  wire  _EVAL_3593;
  wire  _EVAL_3601;
  wire  _EVAL_3607;
  wire  _EVAL_3611;
  wire  _EVAL_3623;
  wire [23:0] _EVAL_3630;
  wire  _EVAL_3707;
  wire  _EVAL_3741;
  wire [31:0] _EVAL_3775;
  wire  _EVAL_3816;
  wire  _EVAL_3820;
  wire [32:0] _EVAL_3837;
  wire  _EVAL_3841;
  wire  _EVAL_3852;
  wire  _EVAL_3858;
  wire  _EVAL_3875;
  wire  _EVAL_3878;
  wire [31:0] _EVAL_3888;
  wire [1:0] _EVAL_3902;
  wire  _EVAL_3930;
  wire [2:0] _EVAL_3973;
  wire [32:0] _EVAL_3993;
  wire  _EVAL_4027;
  wire [31:0] _EVAL_4030;
  wire [32:0] _EVAL_4042;
  wire [31:0] _EVAL_4045;
  wire  _EVAL_4070;
  wire  _EVAL_4090;
  wire [31:0] _EVAL_4157;
  wire  _EVAL_4184;
  wire  _EVAL_4189;
  wire [32:0] _EVAL_4191;
  wire  _EVAL_4213;
  wire  _EVAL_4216;
  wire  _EVAL_4218;
  wire  _EVAL_4257;
  wire  _EVAL_4266;
  wire [23:0] _EVAL_4267;
  wire  _EVAL_4292;
  wire  _EVAL_4295;
  reg [4:0] _EVAL_4297;
  reg [31:0] _RAND_6;
  wire  _EVAL_4323;
  wire  _EVAL_4361;
  wire  _EVAL_4376;
  reg [2:0] _EVAL_4377;
  reg [31:0] _RAND_7;
  wire  _EVAL_4380;
  wire  _EVAL_4381;
  wire  _EVAL_4446;
  wire [31:0] _EVAL_4450;
  wire [3:0] _EVAL_4453;
  wire  _EVAL_4467;
  wire  _EVAL_4469;
  wire  _EVAL_4475;
  wire [2:0] _EVAL_4495;
  wire  _EVAL_4521;
  wire  _EVAL_4545;
  wire  _EVAL_4564;
  wire  _EVAL_4619;
  wire  _EVAL_4626;
  wire [32:0] _EVAL_4646;
  wire  _EVAL_4647;
  wire  _EVAL_4660;
  wire [31:0] _EVAL_4663;
  wire  _EVAL_4673;
  wire  _EVAL_4680;
  wire  _EVAL_4688;
  wire [32:0] _EVAL_4709;
  wire  _EVAL_4753;
  wire [32:0] _EVAL_4798;
  wire  _EVAL_4830;
  wire [10:0] _EVAL_4834;
  wire  _EVAL_4872;
  wire  _EVAL_4888;
  wire [31:0] _EVAL_4897;
  wire  _EVAL_4937;
  wire  _EVAL_4961;
  wire [31:0] _EVAL_4973;
  wire [2:0] _EVAL_5001;
  wire [7:0] _EVAL_5009;
  wire  _EVAL_5049;
  wire  _EVAL_5066;
  wire  _EVAL_5117;
  wire [31:0] _EVAL_5138;
  wire  _EVAL_5146;
  wire  _EVAL_5162;
  wire  _EVAL_5164;
  wire [7:0] _EVAL_5171;
  wire  _EVAL_5227;
  wire  _EVAL_5236;
  wire  _EVAL_5252;
  reg  _EVAL_5301;
  reg [31:0] _RAND_8;
  wire [31:0] _EVAL_5325;
  wire  _EVAL_5332;
  wire [31:0] _EVAL_5341;
  wire  _EVAL_5346;
  wire  _EVAL_5381;
  wire  _EVAL_5387;
  wire  _EVAL_5412;
  wire  _EVAL_5512;
  reg  _EVAL_5564;
  reg [31:0] _RAND_9;
  wire  _EVAL_5566;
  wire [4:0] _EVAL_5579;
  wire  _EVAL_5589;
  wire [2:0] _EVAL_5590;
  wire [31:0] _EVAL_5612;
  wire [32:0] _EVAL_5613;
  wire [31:0] _EVAL_5622;
  wire  _EVAL_5625;
  wire  _EVAL_5648;
  wire [4:0] _EVAL_5671;
  wire  _EVAL_5684;
  wire  _EVAL_5726;
  wire  _EVAL_5728;
  wire  _EVAL_5737;
  wire [32:0] _EVAL_5784;
  wire  _EVAL_5883;
  reg [2:0] _EVAL_5900;
  reg [31:0] _RAND_10;
  wire  _EVAL_5906;
  wire  _EVAL_5907;
  wire [32:0] _EVAL_5908;
  wire [1:0] _EVAL_5933;
  wire  _EVAL_5949;
  wire [10:0] _EVAL_5960;
  wire  _EVAL_5962;
  wire [2:0] _EVAL_6053;
  wire  _EVAL_6057;
  wire  _EVAL_6064;
  wire [31:0] _EVAL_6101;
  wire  _EVAL_6146;
  wire  _EVAL_6156;
  reg [31:0] _EVAL_6190;
  reg [31:0] _RAND_11;
  wire  _EVAL_6196;
  wire [32:0] _EVAL_6214;
  wire  _EVAL_6248;
  wire  _EVAL_6252;
  wire [7:0] _EVAL_6261;
  wire  _EVAL_6265;
  wire  _EVAL_6270;
  wire  _EVAL_6286;
  wire  _EVAL_6328;
  wire  _EVAL_6336;
  wire [31:0] _EVAL_6400;
  wire  _EVAL_6422;
  wire  _EVAL_6449;
  wire  _EVAL_6454;
  wire  _EVAL_6481;
  wire  _EVAL_6492;
  wire [31:0] _EVAL_6530;
  wire  _EVAL_6533;
  reg [4:0] _EVAL_6538;
  reg [31:0] _RAND_12;
  wire  _EVAL_6548;
  wire  _EVAL_6556;
  wire  _EVAL_6571;
  wire  _EVAL_6584;
  wire [31:0] _EVAL_6586;
  wire [31:0] _EVAL_6629;
  reg  _EVAL_6647;
  reg [31:0] _RAND_13;
  wire  _EVAL_6706;
  wire  _EVAL_6719;
  wire [2:0] _EVAL_6735;
  wire  _EVAL_6741;
  wire [32:0] _EVAL_6756;
  wire [31:0] _EVAL_6765;
  wire  _EVAL_6767;
  wire  _EVAL_6770;
  wire  _EVAL_6789;
  reg [3:0] _EVAL_6792;
  reg [31:0] _RAND_14;
  wire  _EVAL_6830;
  wire  _EVAL_6840;
  wire  _EVAL_6884;
  wire [31:0] _EVAL_6918;
  wire  _EVAL_6941;
  wire [31:0] _EVAL_6945;
  wire  _EVAL_6951;
  wire  _EVAL_6999;
  wire  _EVAL_7009;
  wire  _EVAL_7046;
  wire  _EVAL_7053;
  wire  _EVAL_7086;
  wire  _EVAL_7137;
  wire  _EVAL_7142;
  wire  _EVAL_7156;
  wire  _EVAL_7194;
  wire  _EVAL_7201;
  wire [31:0] _EVAL_7342;
  wire  _EVAL_7366;
  wire [32:0] _EVAL_7378;
  wire  _EVAL_7387;
  wire  _EVAL_7407;
  wire [31:0] _EVAL_7414;
  wire [32:0] _EVAL_7483;
  wire  _EVAL_7487;
  wire  _EVAL_7502;
  wire  _EVAL_7611;
  wire [31:0] _EVAL_7614;
  wire [31:0] _EVAL_7616;
  wire  _EVAL_7638;
  wire [32:0] _EVAL_7679;
  wire [31:0] _EVAL_7689;
  reg [1:0] _EVAL_7693;
  reg [31:0] _RAND_15;
  wire [31:0] _EVAL_7717;
  wire  _EVAL_7743;
  wire  _EVAL_7800;
  wire  _EVAL_7809;
  wire  _EVAL_7840;
  wire  _EVAL_7862;
  wire [31:0] _EVAL_7868;
  wire [31:0] _EVAL_7879;
  wire [32:0] _EVAL_7880;
  wire [31:0] _EVAL_7894;
  wire  _EVAL_7895;
  wire  _EVAL_7897;
  wire  _EVAL_7934;
  wire  _EVAL_7993;
  wire  _EVAL_7994;
  wire  _EVAL_8013;
  wire [2:0] _EVAL_8051;
  wire  _EVAL_8070;
  wire  _EVAL_8110;
  wire  _EVAL_8112;
  wire  _EVAL_8116;
  wire [31:0] _EVAL_8128;
  wire  _EVAL_8137;
  wire  _EVAL_8148;
  wire  _EVAL_8163;
  wire  _EVAL_8178;
  wire [32:0] _EVAL_8187;
  wire  _EVAL_8195;
  wire  _EVAL_8200;
  wire [31:0] _EVAL_8228;
  wire [31:0] _EVAL_8292;
  wire [1:0] _EVAL_8299;
  wire  _EVAL_8312;
  wire  _EVAL_8336;
  wire  _EVAL_8339;
  reg  _EVAL_8342;
  reg [31:0] _RAND_16;
  wire  _EVAL_8400;
  wire  _EVAL_8412;
  wire  _EVAL_8452;
  wire  _EVAL_8462;
  wire  bpu__EVAL;
  wire [1:0] bpu__EVAL_0;
  wire  bpu__EVAL_1;
  wire [31:0] bpu__EVAL_2;
  wire  bpu__EVAL_3;
  wire  bpu__EVAL_4;
  wire  bpu__EVAL_5;
  wire  bpu__EVAL_6;
  wire  bpu__EVAL_7;
  wire [31:0] bpu__EVAL_8;
  wire [1:0] bpu__EVAL_9;
  wire  bpu__EVAL_10;
  wire  bpu__EVAL_11;
  wire [31:0] bpu__EVAL_12;
  wire [31:0] bpu__EVAL_13;
  wire [31:0] bpu__EVAL_14;
  wire [1:0] bpu__EVAL_15;
  wire [31:0] bpu__EVAL_16;
  wire  bpu__EVAL_17;
  wire  bpu__EVAL_18;
  wire  bpu__EVAL_19;
  wire  bpu__EVAL_20;
  wire  bpu__EVAL_21;
  wire  bpu__EVAL_22;
  wire  bpu__EVAL_23;
  wire  bpu__EVAL_24;
  wire  bpu__EVAL_25;
  wire [1:0] bpu__EVAL_26;
  wire  bpu__EVAL_27;
  wire  bpu__EVAL_28;
  wire  bpu__EVAL_29;
  wire  bpu__EVAL_30;
  wire  bpu__EVAL_31;
  wire  bpu__EVAL_32;
  wire  bpu__EVAL_33;
  wire  bpu__EVAL_34;
  wire  bpu__EVAL_35;
  wire  bpu__EVAL_36;
  wire  bpu__EVAL_37;
  wire  bpu__EVAL_38;
  wire [1:0] bpu__EVAL_39;
  wire  bpu__EVAL_40;
  wire  bpu__EVAL_41;
  wire  bpu__EVAL_42;
  wire  bpu__EVAL_43;
  wire [32:0] _EVAL_8522;
  wire  _EVAL_8534;
  reg [4:0] _EVAL_8580;
  reg [31:0] _RAND_17;
  wire  _EVAL_8584;
  wire [31:0] _EVAL_8601;
  wire  _EVAL_8607;
  wire  _EVAL_8610;
  wire  _EVAL_8621;
  wire  _EVAL_8627;
  reg [31:0] _EVAL_8631;
  reg [31:0] _RAND_18;
  wire [31:0] _EVAL_8646;
  wire [32:0] _EVAL_8649;
  wire  _EVAL_8672;
  wire  _EVAL_8698;
  wire  _EVAL_8702;
  wire  _EVAL_8706;
  wire [3:0] _EVAL_8759;
  wire  _EVAL_8864;
  wire  _EVAL_8865;
  wire [23:0] _EVAL_8869;
  wire  _EVAL_8872;
  wire  _EVAL_8873;
  reg  _EVAL_8874;
  reg [31:0] _RAND_19;
  wire  _EVAL_8892;
  wire  _EVAL_8899;
  wire [32:0] _EVAL_8912;
  wire  _EVAL_8917;
  wire  _EVAL_8923;
  wire  _EVAL_8949;
  wire  _EVAL_8958;
  wire  _EVAL_8990;
  reg  _EVAL_8999;
  reg [31:0] _RAND_20;
  wire [31:0] _EVAL_9039;
  wire  _EVAL_9061;
  wire  _EVAL_9066;
  wire [15:0] _EVAL_9075;
  wire  _EVAL_9086;
  reg  _EVAL_9119;
  reg [31:0] _RAND_21;
  wire [31:0] _EVAL_9169;
  wire  _EVAL_9183;
  wire  _EVAL_9187;
  wire [31:0] _EVAL_9241;
  wire  _EVAL_9277;
  wire  _EVAL_9300;
  wire [32:0] _EVAL_9314;
  wire  _EVAL_9364;
  wire  _EVAL_9376;
  wire  _EVAL_9378;
  wire  _EVAL_9383;
  wire  _EVAL_9411;
  reg  _EVAL_9429;
  reg [31:0] _RAND_22;
  reg  _EVAL_9449;
  reg [31:0] _RAND_23;
  wire  _EVAL_9451;
  wire  _EVAL_9464;
  wire  _EVAL_9472;
  wire  _EVAL_9491;
  wire  _EVAL_9496;
  reg  _EVAL_9510;
  reg [31:0] _RAND_24;
  wire  _EVAL_9514;
  wire  _EVAL_9545;
  wire [31:0] _EVAL_9548;
  wire  _EVAL_9556;
  wire  _EVAL_9565;
  wire  _EVAL_9583;
  wire  _EVAL_9589;
  wire  _EVAL_9594;
  wire  _EVAL_9658;
  wire  _EVAL_9667;
  wire  _EVAL_9689;
  wire [10:0] _EVAL_9697;
  wire  _EVAL_9700;
  wire  _EVAL_9734;
  wire [31:0] _EVAL_9768;
  wire [31:0] _EVAL_9792;
  wire [31:0] _EVAL_9820;
  wire [31:0] _EVAL_9822;
  wire [31:0] _EVAL_9843;
  wire  _EVAL_9882;
  wire  _EVAL_9896;
  wire  _EVAL_9941;
  wire  _EVAL_9965;
  wire  _EVAL_10012;
  wire [32:0] _EVAL_10019;
  wire  _EVAL_10051;
  wire  _EVAL_10091;
  wire [3:0] _EVAL_10107;
  wire  _EVAL_10111;
  wire  _EVAL_10114;
  wire [31:0] _EVAL_10127;
  wire  _EVAL_10140;
  wire  _EVAL_10147;
  wire [31:0] _EVAL_10148;
  wire  _EVAL_10156;
  wire  _EVAL_10181;
  wire  _EVAL_10207;
  wire  _EVAL_10233;
  wire  _EVAL_10239;
  wire  _EVAL_10284;
  wire  _EVAL_10289;
  wire  _EVAL_10302;
  wire [31:0] _EVAL_10331;
  reg [31:0] _EVAL_10347;
  reg [31:0] _RAND_25;
  reg [4:0] _EVAL_10353;
  reg [31:0] _RAND_26;
  wire  _EVAL_10368;
  wire  _EVAL_10371;
  wire [4:0] _EVAL_10383;
  wire  _EVAL_10444;
  reg  _EVAL_10468;
  reg [31:0] _RAND_27;
  wire [31:0] _EVAL_10480;
  wire [15:0] _EVAL_10491;
  wire [2:0] _EVAL_10553;
  wire [31:0] rf__EVAL;
  wire [31:0] rf__EVAL_0;
  wire [4:0] rf__EVAL_1;
  wire [31:0] rf__EVAL_2;
  wire [4:0] rf__EVAL_3;
  wire  rf__EVAL_4;
  wire [4:0] rf__EVAL_5;
  wire  rf__EVAL_6;
  wire  _EVAL_10566;
  wire [31:0] _EVAL_10588;
  reg  _EVAL_10593;
  reg [31:0] _RAND_28;
  wire  _EVAL_10622;
  wire [31:0] _EVAL_10627;
  wire [32:0] _EVAL_10668;
  wire  _EVAL_10679;
  wire [2:0] _EVAL_10692;
  wire  _EVAL_10735;
  wire [7:0] _EVAL_10764;
  wire  _EVAL_10778;
  wire  _EVAL_10782;
  wire [32:0] _EVAL_10803;
  wire  _EVAL_10825;
  wire  _EVAL_10831;
  wire  _EVAL_10856;
  wire  _EVAL_10858;
  reg [31:0] _EVAL_10894;
  reg [31:0] _RAND_29;
  wire  _EVAL_10896;
  wire  _EVAL_10919;
  wire  _EVAL_10928;
  wire  _EVAL_10948;
  wire  _EVAL_10975;
  wire  _EVAL_11005;
  wire  _EVAL_11046;
  wire [4:0] alu__EVAL;
  wire [31:0] alu__EVAL_0;
  wire [31:0] alu__EVAL_1;
  wire [31:0] alu__EVAL_2;
  wire [31:0] alu__EVAL_3;
  wire [31:0] _EVAL_11129;
  wire  _EVAL_11154;
  reg  _EVAL_11162;
  reg [31:0] _RAND_30;
  wire  _EVAL_11178;
  wire [31:0] _EVAL_11189;
  wire  _EVAL_11215;
  wire  _EVAL_11218;
  wire [15:0] _EVAL_11230;
  wire  _EVAL_11251;
  wire [15:0] _EVAL_11252;
  wire  _EVAL_11278;
  wire  _EVAL_11286;
  wire  _EVAL_11311;
  wire  _EVAL_11321;
  wire  _EVAL_11327;
  wire [15:0] _EVAL_11356;
  wire [7:0] _EVAL_11436;
  wire [31:0] _EVAL_11443;
  wire  fetch__EVAL;
  wire [31:0] fetch__EVAL_0;
  wire  fetch__EVAL_1;
  wire [4:0] fetch__EVAL_2;
  wire [4:0] fetch__EVAL_3;
  wire  fetch__EVAL_4;
  wire  fetch__EVAL_5;
  wire  fetch__EVAL_6;
  wire [4:0] fetch__EVAL_7;
  wire  fetch__EVAL_8;
  wire  fetch__EVAL_9;
  wire  fetch__EVAL_10;
  wire [31:0] fetch__EVAL_11;
  wire  fetch__EVAL_12;
  wire [31:0] fetch__EVAL_13;
  wire  fetch__EVAL_14;
  wire [31:0] fetch__EVAL_15;
  wire  fetch__EVAL_16;
  wire [4:0] fetch__EVAL_17;
  wire  fetch__EVAL_18;
  wire  fetch__EVAL_19;
  wire  fetch__EVAL_20;
  wire [31:0] fetch__EVAL_21;
  wire  fetch__EVAL_22;
  wire  fetch__EVAL_23;
  wire  _EVAL_11458;
  wire [31:0] _EVAL_11480;
  wire [32:0] _EVAL_11503;
  wire  _EVAL_11504;
  wire  _EVAL_11521;
  wire  _EVAL_11531;
  wire [2:0] _EVAL_11533;
  wire [1:0] _EVAL_11557;
  wire [4:0] _EVAL_11561;
  wire  _EVAL_11578;
  wire  _EVAL_11596;
  wire [31:0] _EVAL_11607;
  wire  _EVAL_11609;
  wire [23:0] _EVAL_11610;
  wire  _EVAL_11613;
  wire  _EVAL_11654;
  wire  _EVAL_11701;
  wire [2:0] _EVAL_11712;
  wire  _EVAL_11716;
  wire  _EVAL_11801;
  wire  _EVAL_11807;
  wire  _EVAL_11823;
  wire  _EVAL_11838;
  wire  _EVAL_11858;
  wire [32:0] _EVAL_11868;
  wire  _EVAL_11875;
  wire  _EVAL_11894;
  wire [32:0] _EVAL_11900;
  wire  _EVAL_11919;
  wire  _EVAL_12009;
  wire  _EVAL_12010;
  wire  _EVAL_12018;
  wire  _EVAL_12043;
  wire [31:0] _EVAL_12058;
  wire [31:0] _EVAL_12083;
  wire  _EVAL_12096;
  wire [4:0] _EVAL_12112;
  wire [1:0] _EVAL_12173;
  wire  _EVAL_12191;
  wire  _EVAL_12216;
  wire [2:0] _EVAL_12232;
  wire [3:0] _EVAL_12244;
  wire  _EVAL_12247;
  wire [31:0] _EVAL_12251;
  wire  _EVAL_12263;
  wire [2:0] _EVAL_12268;
  wire  _EVAL_12282;
  wire  _EVAL_12302;
  wire [32:0] _EVAL_12339;
  wire [31:0] _EVAL_12352;
  wire  _EVAL_12356;
  wire [31:0] _EVAL_12360;
  reg  _EVAL_12371;
  reg [31:0] _RAND_31;
  wire [1:0] _EVAL_12376;
  reg  _EVAL_12379;
  reg [31:0] _RAND_32;
  wire  _EVAL_12395;
  wire [31:0] _EVAL_12411;
  wire [31:0] _EVAL_12413;
  wire [2:0] _EVAL_12424;
  wire  _EVAL_12427;
  wire [1:0] _EVAL_12438;
  wire  _EVAL_12439;
  wire [32:0] _EVAL_12444;
  wire  _EVAL_12468;
  wire  _EVAL_12476;
  wire  _EVAL_12477;
  reg  _EVAL_12498;
  reg [31:0] _RAND_33;
  wire  _EVAL_12502;
  wire [2:0] _EVAL_12503;
  reg  _EVAL_12508;
  reg [31:0] _RAND_34;
  wire  _EVAL_12521;
  wire [2:0] _EVAL_12525;
  wire  _EVAL_12529;
  wire  _EVAL_12545;
  wire  _EVAL_12548;
  wire  _EVAL_12566;
  wire  _EVAL_12568;
  wire  _EVAL_12589;
  wire  _EVAL_12601;
  wire  _EVAL_12603;
  wire  _EVAL_12608;
  wire [32:0] _EVAL_12611;
  wire  _EVAL_12623;
  wire [31:0] _EVAL_12651;
  wire  _EVAL_12682;
  reg [31:0] _EVAL_12724;
  reg [31:0] _RAND_35;
  wire  _EVAL_12732;
  wire  _EVAL_12751;
  wire [7:0] _EVAL_12793;
  wire  _EVAL_12794;
  wire [31:0] _EVAL_12823;
  wire [3:0] _EVAL_12829;
  wire  _EVAL_12850;
  wire  _EVAL_12887;
  wire [3:0] _EVAL_12929;
  wire  _EVAL_12957;
  wire  _EVAL_12967;
  wire  _EVAL_12968;
  wire  _EVAL_12981;
  wire [32:0] _EVAL_13002;
  wire [31:0] _EVAL_13006;
  wire [32:0] _EVAL_13007;
  wire [15:0] _EVAL_13022;
  wire [31:0] _EVAL_13045;
  wire  _EVAL_13047;
  wire [31:0] _EVAL_13052;
  wire  _EVAL_13053;
  wire [31:0] _EVAL_13072;
  wire  _EVAL_13093;
  wire  _EVAL_13097;
  wire  _EVAL_13099;
  wire  _EVAL_13129;
  wire  _EVAL_13130;
  wire [3:0] _EVAL_13133;
  wire  _EVAL_13139;
  wire  _EVAL_13144;
  wire  _EVAL_13157;
  wire  _EVAL_13158;
  wire [31:0] _EVAL_13170;
  wire  _EVAL_13198;
  wire  _EVAL_13210;
  wire  _EVAL_13225;
  wire  _EVAL_13253;
  wire [2:0] _EVAL_13287;
  wire  _EVAL_13298;
  wire  _EVAL_13304;
  wire  _EVAL_13311;
  reg  _EVAL_13327;
  reg [31:0] _RAND_36;
  wire  _EVAL_13371;
  wire [32:0] _EVAL_13389;
  wire  _EVAL_13586;
  wire  _EVAL_13609;
  wire [31:0] _EVAL_13687;
  wire [32:0] _EVAL_13694;
  wire  _EVAL_13703;
  wire  _EVAL_13706;
  wire  _EVAL_13723;
  wire [5:0] _EVAL_13735;
  wire [2:0] _EVAL_13756;
  wire [31:0] _EVAL_13761;
  wire  _EVAL_13772;
  wire [3:0] _EVAL_13825;
  wire  _EVAL_13835;
  wire  _EVAL_13874;
  wire  _EVAL_13906;
  wire  _EVAL_13977;
  wire  _EVAL_14001;
  wire [3:0] _EVAL_14010;
  wire  _EVAL_14011;
  wire  _EVAL_14051;
  wire  _EVAL_14053;
  wire  _EVAL_14092;
  wire  _EVAL_14107;
  wire [32:0] _EVAL_14115;
  wire  _EVAL_14142;
  wire [31:0] _EVAL_14156;
  wire  _EVAL_14159;
  reg  _EVAL_14160;
  reg [31:0] _RAND_37;
  wire  _EVAL_14169;
  wire [31:0] _EVAL_14183;
  reg [31:0] _EVAL_14184;
  reg [31:0] _RAND_38;
  wire [7:0] _EVAL_14196;
  wire  _EVAL_14231;
  wire [31:0] _EVAL_14251;
  wire [31:0] _EVAL_14257;
  wire [32:0] _EVAL_14263;
  wire  _EVAL_14322;
  wire  _EVAL_14355;
  wire  _EVAL_14356;
  wire  _EVAL_14418;
  wire  _EVAL_14448;
  reg  _EVAL_14478;
  reg [31:0] _RAND_39;
  wire [31:0] _EVAL_14573;
  wire [3:0] _EVAL_14650;
  wire  _EVAL_14680;
  wire  _EVAL_14682;
  wire [31:0] _EVAL_14722;
  wire  _EVAL_14726;
  wire  _EVAL_14763;
  wire [31:0] _EVAL_14765;
  wire [32:0] _EVAL_14767;
  wire [31:0] _EVAL_14777;
  wire [2:0] _EVAL_14804;
  wire  _EVAL_14808;
  wire  _EVAL_14809;
  wire [32:0] _EVAL_14814;
  wire  _EVAL_14832;
  wire  _EVAL_14855;
  wire  _EVAL_14879;
  wire  _EVAL_14892;
  reg [4:0] _EVAL_14896;
  reg [31:0] _RAND_40;
  wire [4:0] _EVAL_14920;
  wire [32:0] _EVAL_14959;
  wire  _EVAL_14969;
  wire  _EVAL_15003;
  wire  _EVAL_15039;
  wire [31:0] _EVAL_15053;
  wire [1:0] _EVAL_15097;
  wire  _EVAL_15106;
  wire  _EVAL_15112;
  wire [4:0] _EVAL_15130;
  wire [31:0] _EVAL_15131;
  wire  _EVAL_15156;
  wire  _EVAL_15184;
  wire [4:0] _EVAL_15219;
  wire [32:0] _EVAL_15238;
  wire  _EVAL_15242;
  wire  _EVAL_15272;
  wire  _EVAL_15312;
  wire  _EVAL_15340;
  wire  _EVAL_15349;
  wire  _EVAL_15382;
  wire [2:0] _EVAL_15396;
  wire [31:0] _EVAL_15398;
  wire  _EVAL_15409;
  wire  _EVAL_15411;
  wire [10:0] _EVAL_15418;
  wire  _EVAL_15427;
  wire  _EVAL_15431;
  wire  _EVAL_15453;
  wire  _EVAL_15461;
  wire  _EVAL_15467;
  wire  _EVAL_15479;
  wire  _EVAL_15497;
  wire [31:0] _EVAL_15504;
  wire  _EVAL_15511;
  wire  _EVAL_15526;
  reg [4:0] _EVAL_15545;
  reg [31:0] _RAND_41;
  wire  _EVAL_15553;
  wire  _EVAL_15561;
  wire [4:0] _EVAL_15591;
  wire  _EVAL_15596;
  wire [31:0] _EVAL_15617;
  wire  _EVAL_15648;
  wire  _EVAL_15656;
  wire [31:0] _EVAL_15690;
  wire [2:0] _EVAL_15723;
  wire [32:0] _EVAL_15755;
  reg  _EVAL_15759;
  reg [31:0] _RAND_42;
  wire [31:0] _EVAL_15765;
  wire  _EVAL_15768;
  wire [31:0] _EVAL_15785;
  wire  _EVAL_15801;
  wire  _EVAL_15829;
  wire  pmp_checker__EVAL;
  wire  pmp_checker__EVAL_0;
  wire [31:0] pmp_checker__EVAL_1;
  wire [1:0] pmp_checker__EVAL_2;
  wire  pmp_checker__EVAL_3;
  wire  pmp_checker__EVAL_4;
  wire  pmp_checker__EVAL_5;
  wire  pmp_checker__EVAL_6;
  wire  pmp_checker__EVAL_7;
  wire  pmp_checker__EVAL_8;
  wire  pmp_checker__EVAL_9;
  wire [29:0] pmp_checker__EVAL_10;
  wire [1:0] pmp_checker__EVAL_11;
  wire [31:0] pmp_checker__EVAL_12;
  wire  pmp_checker__EVAL_13;
  wire [29:0] pmp_checker__EVAL_14;
  wire  pmp_checker__EVAL_15;
  wire  pmp_checker__EVAL_16;
  wire [29:0] pmp_checker__EVAL_17;
  wire  pmp_checker__EVAL_18;
  wire [31:0] pmp_checker__EVAL_19;
  wire [1:0] pmp_checker__EVAL_20;
  wire  pmp_checker__EVAL_21;
  wire  pmp_checker__EVAL_22;
  wire [1:0] pmp_checker__EVAL_23;
  wire  pmp_checker__EVAL_24;
  wire [29:0] pmp_checker__EVAL_25;
  wire [31:0] pmp_checker__EVAL_26;
  wire  pmp_checker__EVAL_27;
  wire  pmp_checker__EVAL_28;
  wire  pmp_checker__EVAL_29;
  wire [1:0] pmp_checker__EVAL_30;
  wire  pmp_checker__EVAL_31;
  wire [31:0] pmp_checker__EVAL_32;
  wire  pmp_checker__EVAL_33;
  wire  _EVAL_15856;
  wire  _EVAL_15870;
  wire  _EVAL_15890;
  wire  _EVAL_15910;
  wire [31:0] _EVAL_15947;
  wire [7:0] _EVAL_15968;
  wire  _EVAL_15974;
  wire  _EVAL_15976;
  wire  _EVAL_15981;
  wire  _EVAL_16024;
  reg  _EVAL_16030;
  reg [31:0] _RAND_43;
  wire  _EVAL_16034;
  wire [31:0] _EVAL_16060;
  wire  _EVAL_16067;
  wire  _EVAL_16094;
  reg  _EVAL_16096;
  reg [31:0] _RAND_44;
  wire  _EVAL_16155;
  wire  _EVAL_16164;
  wire  _EVAL_16173;
  wire  _EVAL_16200;
  wire  _EVAL_16201;
  wire  _EVAL_16202;
  reg [31:0] _EVAL_16207;
  reg [31:0] _RAND_45;
  wire [2:0] _EVAL_16227;
  wire  _EVAL_16256;
  wire [31:0] _EVAL_16288;
  wire  _EVAL_16306;
  wire  _EVAL_16323;
  wire  _EVAL_16351;
  wire [31:0] _EVAL_16377;
  wire  _EVAL_16380;
  wire  _EVAL_16389;
  wire  _EVAL_16392;
  wire [3:0] _EVAL_16395;
  wire  _EVAL_16398;
  wire  _EVAL_16407;
  wire  _EVAL_16447;
  wire  _EVAL_16448;
  wire [1:0] _EVAL_16483;
  reg  _EVAL_16543;
  reg [31:0] _RAND_46;
  wire [1:0] _EVAL_16547;
  wire  _EVAL_16592;
  wire [31:0] _EVAL_16593;
  wire [31:0] _EVAL_16620;
  reg [31:0] _EVAL_16644;
  reg [31:0] _RAND_47;
  wire  _EVAL_16647;
  wire  _EVAL_16649;
  wire  _EVAL_16668;
  wire [31:0] _EVAL_16692;
  wire  _EVAL_16722;
  reg  _EVAL_16733;
  reg [31:0] _RAND_48;
  wire  _EVAL_16739;
  wire [7:0] _EVAL_16751;
  reg [31:0] _EVAL_16768;
  reg [31:0] _RAND_49;
  wire  _EVAL_16772;
  wire  _EVAL_16796;
  wire  _EVAL_16804;
  wire  _EVAL_16854;
  wire  _EVAL_16866;
  wire [31:0] _EVAL_16867;
  wire [31:0] _EVAL_16869;
  wire [31:0] _EVAL_16872;
  wire  _EVAL_16877;
  wire [23:0] _EVAL_16898;
  wire [3:0] _EVAL_16949;
  wire  csr__EVAL;
  wire  csr__EVAL_0;
  wire [1:0] csr__EVAL_1;
  wire  csr__EVAL_2;
  wire [1:0] csr__EVAL_3;
  wire [31:0] csr__EVAL_4;
  wire [31:0] csr__EVAL_5;
  wire [31:0] csr__EVAL_6;
  wire  csr__EVAL_7;
  wire  csr__EVAL_8;
  wire  csr__EVAL_9;
  wire  csr__EVAL_10;
  wire  csr__EVAL_11;
  wire  csr__EVAL_12;
  wire  csr__EVAL_13;
  wire  csr__EVAL_14;
  wire [7:0] csr__EVAL_15;
  wire  csr__EVAL_16;
  wire [31:0] csr__EVAL_17;
  wire [31:0] csr__EVAL_18;
  wire [31:0] csr__EVAL_19;
  wire  csr__EVAL_20;
  wire  csr__EVAL_21;
  wire  csr__EVAL_22;
  wire  csr__EVAL_23;
  wire  csr__EVAL_24;
  wire [29:0] csr__EVAL_25;
  wire [31:0] csr__EVAL_26;
  wire  csr__EVAL_27;
  wire  csr__EVAL_28;
  wire [31:0] csr__EVAL_29;
  wire [31:0] csr__EVAL_30;
  wire  csr__EVAL_31;
  wire  csr__EVAL_32;
  wire  csr__EVAL_33;
  wire [31:0] csr__EVAL_34;
  wire  csr__EVAL_35;
  wire [1:0] csr__EVAL_36;
  wire [31:0] csr__EVAL_37;
  wire [1:0] csr__EVAL_38;
  wire  csr__EVAL_39;
  wire  csr__EVAL_40;
  wire [1:0] csr__EVAL_41;
  wire  csr__EVAL_42;
  wire  csr__EVAL_43;
  wire  csr__EVAL_44;
  wire  csr__EVAL_45;
  wire [29:0] csr__EVAL_46;
  wire [31:0] csr__EVAL_47;
  wire  csr__EVAL_48;
  wire  csr__EVAL_49;
  wire  csr__EVAL_50;
  wire [31:0] csr__EVAL_51;
  wire  csr__EVAL_52;
  wire  csr__EVAL_53;
  wire  csr__EVAL_54;
  wire [7:0] csr__EVAL_55;
  wire [1:0] csr__EVAL_56;
  wire  csr__EVAL_57;
  wire  csr__EVAL_58;
  wire  csr__EVAL_59;
  wire  csr__EVAL_60;
  wire  csr__EVAL_61;
  wire [1:0] csr__EVAL_62;
  wire  csr__EVAL_63;
  wire [31:0] csr__EVAL_64;
  wire [1:0] csr__EVAL_65;
  wire  csr__EVAL_66;
  wire  csr__EVAL_67;
  wire [29:0] csr__EVAL_68;
  wire  csr__EVAL_69;
  wire  csr__EVAL_70;
  wire  csr__EVAL_71;
  wire  csr__EVAL_72;
  wire [31:0] csr__EVAL_73;
  wire  csr__EVAL_74;
  wire  csr__EVAL_75;
  wire [11:0] csr__EVAL_76;
  wire  csr__EVAL_77;
  wire  csr__EVAL_78;
  wire [31:0] csr__EVAL_79;
  wire  csr__EVAL_80;
  wire [31:0] csr__EVAL_81;
  wire  csr__EVAL_82;
  wire [31:0] csr__EVAL_83;
  wire  csr__EVAL_84;
  wire [31:0] csr__EVAL_85;
  wire [29:0] csr__EVAL_86;
  wire  csr__EVAL_87;
  wire  csr__EVAL_88;
  wire [1:0] csr__EVAL_89;
  wire [31:0] csr__EVAL_90;
  wire [31:0] csr__EVAL_91;
  wire  csr__EVAL_92;
  wire  csr__EVAL_93;
  wire  csr__EVAL_94;
  wire [2:0] csr__EVAL_95;
  wire  csr__EVAL_96;
  wire  csr__EVAL_97;
  wire [2:0] csr__EVAL_98;
  wire  csr__EVAL_99;
  wire  csr__EVAL_100;
  wire [11:0] csr__EVAL_101;
  wire  csr__EVAL_102;
  wire  csr__EVAL_103;
  wire [1:0] csr__EVAL_104;
  wire  csr__EVAL_105;
  wire  csr__EVAL_106;
  wire [31:0] csr__EVAL_107;
  wire [7:0] csr__EVAL_108;
  wire [31:0] csr__EVAL_109;
  wire  csr__EVAL_110;
  wire  csr__EVAL_111;
  wire  csr__EVAL_112;
  wire  csr__EVAL_113;
  wire  csr__EVAL_114;
  wire  csr__EVAL_115;
  wire [1:0] csr__EVAL_116;
  wire  csr__EVAL_117;
  wire  csr__EVAL_118;
  wire  csr__EVAL_119;
  wire  csr__EVAL_120;
  wire  csr__EVAL_121;
  wire  csr__EVAL_122;
  wire  csr__EVAL_123;
  wire  csr__EVAL_124;
  wire [26:0] csr__EVAL_125;
  wire  csr__EVAL_126;
  wire [1:0] csr__EVAL_127;
  wire [1:0] csr__EVAL_128;
  wire [1:0] csr__EVAL_129;
  wire [1:0] csr__EVAL_130;
  wire  csr__EVAL_131;
  wire  csr__EVAL_132;
  wire [31:0] csr__EVAL_133;
  wire  csr__EVAL_134;
  wire [1:0] csr__EVAL_135;
  wire  csr__EVAL_136;
  wire [1:0] csr__EVAL_137;
  wire  csr__EVAL_138;
  wire  csr__EVAL_139;
  wire  csr__EVAL_140;
  wire [1:0] csr__EVAL_141;
  wire [31:0] _EVAL_17033;
  wire  _EVAL_17054;
  wire  _EVAL_17074;
  wire [15:0] _EVAL_17093;
  wire  _EVAL_17118;
  wire  _EVAL_17140;
  wire  _EVAL_17194;
  wire  _EVAL_17211;
  wire  _EVAL_17213;
  wire  _EVAL_17240;
  wire  _EVAL_17254;
  wire  _EVAL_17283;
  wire [32:0] _EVAL_17285;
  wire  _EVAL_17352;
  wire  _EVAL_17356;
  wire  _EVAL_17358;
  reg  _EVAL_17371;
  reg [31:0] _RAND_50;
  wire  _EVAL_17383;
  wire [31:0] _EVAL_17384;
  wire [31:0] _EVAL_17404;
  wire  _EVAL_17447;
  wire [31:0] _EVAL_17451;
  wire [2:0] _EVAL_17519;
  wire  _EVAL_17543;
  wire [23:0] _EVAL_17544;
  wire [1:0] _EVAL_17546;
  wire [31:0] _EVAL_17560;
  wire  _EVAL_17570;
  wire  _EVAL_17583;
  wire  _EVAL_17584;
  wire  _EVAL_17589;
  wire  _EVAL_17605;
  wire  _EVAL_17608;
  wire  _EVAL_17625;
  wire  _EVAL_17640;
  wire  _EVAL_17674;
  wire  _EVAL_17688;
  wire  _EVAL_17705;
  wire  _EVAL_17716;
  wire [1:0] _EVAL_17717;
  wire [31:0] _EVAL_17736;
  wire  _EVAL_17740;
  wire [31:0] _EVAL_17779;
  reg  _EVAL_17801;
  reg [31:0] _RAND_51;
  wire [2:0] _EVAL_17805;
  wire  _EVAL_17821;
  wire  _EVAL_17827;
  wire  _EVAL_17840;
  wire  _EVAL_17854;
  wire  _EVAL_17886;
  wire  _EVAL_17887;
  wire [31:0] _EVAL_17909;
  wire  _EVAL_17934;
  wire  _EVAL_17953;
  wire  _EVAL_17963;
  wire  _EVAL_17967;
  wire  _EVAL_17986;
  wire  _EVAL_17995;
  wire [3:0] _EVAL_17997;
  wire  _EVAL_18030;
  wire [10:0] _EVAL_18078;
  wire  _EVAL_18119;
  wire [31:0] _EVAL_18125;
  wire  _EVAL_18141;
  wire  _EVAL_18202;
  wire [31:0] _EVAL_18210;
  wire  _EVAL_18216;
  wire  _EVAL_18247;
  wire  _EVAL_18258;
  wire  _EVAL_18289;
  wire  _EVAL_18360;
  wire  _EVAL_18361;
  wire [2:0] _EVAL_18401;
  wire  _EVAL_18410;
  wire  _EVAL_18439;
  wire  _EVAL_18449;
  wire [31:0] _EVAL_18452;
  reg  _EVAL_18514;
  reg [31:0] _RAND_52;
  wire  _EVAL_18565;
  wire [1:0] _EVAL_18613;
  wire  _EVAL_18618;
  wire  _EVAL_18634;
  wire  _EVAL_18642;
  wire [31:0] _EVAL_18671;
  wire  _EVAL_18675;
  wire [32:0] _EVAL_18697;
  wire  _EVAL_18765;
  wire  _EVAL_18773;
  wire [10:0] _EVAL_18791;
  wire  _EVAL_18800;
  wire  _EVAL_18877;
  wire  _EVAL_18905;
  wire  _EVAL_18912;
  wire  _EVAL_18942;
  wire [32:0] _EVAL_18960;
  wire  div__EVAL;
  wire [31:0] div__EVAL_0;
  wire  div__EVAL_1;
  wire  div__EVAL_2;
  wire  div__EVAL_3;
  wire [31:0] div__EVAL_4;
  wire  div__EVAL_5;
  wire  div__EVAL_6;
  wire [31:0] div__EVAL_7;
  wire [3:0] div__EVAL_8;
  wire  _EVAL_18990;
  wire  _EVAL_19013;
  wire  _EVAL_19031;
  wire [31:0] _EVAL_19059;
  wire [2:0] _EVAL_19090;
  wire  _EVAL_19144;
  wire  _EVAL_19208;
  wire [31:0] _EVAL_19212;
  wire [7:0] _EVAL_19273;
  wire [3:0] _EVAL_19285;
  wire  _EVAL_19297;
  wire  _EVAL_19336;
  wire [32:0] _EVAL_19337;
  wire  _EVAL_19340;
  wire  _EVAL_19347;
  wire [1:0] _EVAL_19357;
  wire  _EVAL_19368;
  wire [2:0] _EVAL_19408;
  wire  _EVAL_19413;
  wire  _EVAL_19430;
  wire  _EVAL_19458;
  wire  _EVAL_19509;
  wire  _EVAL_19529;
  wire [31:0] _EVAL_19544;
  reg [2:0] _EVAL_19551;
  reg [31:0] _RAND_53;
  wire  _EVAL_19578;
  wire  _EVAL_19597;
  wire [7:0] _EVAL_19607;
  wire  _EVAL_19610;
  wire [31:0] _EVAL_19611;
  _EVAL_156 fetch_pmp_checker (
    ._EVAL(fetch_pmp_checker__EVAL),
    ._EVAL_0(fetch_pmp_checker__EVAL_0),
    ._EVAL_1(fetch_pmp_checker__EVAL_1),
    ._EVAL_2(fetch_pmp_checker__EVAL_2),
    ._EVAL_3(fetch_pmp_checker__EVAL_3),
    ._EVAL_4(fetch_pmp_checker__EVAL_4),
    ._EVAL_5(fetch_pmp_checker__EVAL_5),
    ._EVAL_6(fetch_pmp_checker__EVAL_6),
    ._EVAL_7(fetch_pmp_checker__EVAL_7),
    ._EVAL_8(fetch_pmp_checker__EVAL_8),
    ._EVAL_9(fetch_pmp_checker__EVAL_9),
    ._EVAL_10(fetch_pmp_checker__EVAL_10),
    ._EVAL_11(fetch_pmp_checker__EVAL_11),
    ._EVAL_12(fetch_pmp_checker__EVAL_12),
    ._EVAL_13(fetch_pmp_checker__EVAL_13),
    ._EVAL_14(fetch_pmp_checker__EVAL_14),
    ._EVAL_15(fetch_pmp_checker__EVAL_15),
    ._EVAL_16(fetch_pmp_checker__EVAL_16),
    ._EVAL_17(fetch_pmp_checker__EVAL_17),
    ._EVAL_18(fetch_pmp_checker__EVAL_18),
    ._EVAL_19(fetch_pmp_checker__EVAL_19),
    ._EVAL_20(fetch_pmp_checker__EVAL_20),
    ._EVAL_21(fetch_pmp_checker__EVAL_21),
    ._EVAL_22(fetch_pmp_checker__EVAL_22),
    ._EVAL_23(fetch_pmp_checker__EVAL_23),
    ._EVAL_24(fetch_pmp_checker__EVAL_24),
    ._EVAL_25(fetch_pmp_checker__EVAL_25),
    ._EVAL_26(fetch_pmp_checker__EVAL_26),
    ._EVAL_27(fetch_pmp_checker__EVAL_27),
    ._EVAL_28(fetch_pmp_checker__EVAL_28),
    ._EVAL_29(fetch_pmp_checker__EVAL_29),
    ._EVAL_30(fetch_pmp_checker__EVAL_30),
    ._EVAL_31(fetch_pmp_checker__EVAL_31),
    ._EVAL_32(fetch_pmp_checker__EVAL_32),
    ._EVAL_33(fetch_pmp_checker__EVAL_33)
  );
  _EVAL_157 bpu (
    ._EVAL(bpu__EVAL),
    ._EVAL_0(bpu__EVAL_0),
    ._EVAL_1(bpu__EVAL_1),
    ._EVAL_2(bpu__EVAL_2),
    ._EVAL_3(bpu__EVAL_3),
    ._EVAL_4(bpu__EVAL_4),
    ._EVAL_5(bpu__EVAL_5),
    ._EVAL_6(bpu__EVAL_6),
    ._EVAL_7(bpu__EVAL_7),
    ._EVAL_8(bpu__EVAL_8),
    ._EVAL_9(bpu__EVAL_9),
    ._EVAL_10(bpu__EVAL_10),
    ._EVAL_11(bpu__EVAL_11),
    ._EVAL_12(bpu__EVAL_12),
    ._EVAL_13(bpu__EVAL_13),
    ._EVAL_14(bpu__EVAL_14),
    ._EVAL_15(bpu__EVAL_15),
    ._EVAL_16(bpu__EVAL_16),
    ._EVAL_17(bpu__EVAL_17),
    ._EVAL_18(bpu__EVAL_18),
    ._EVAL_19(bpu__EVAL_19),
    ._EVAL_20(bpu__EVAL_20),
    ._EVAL_21(bpu__EVAL_21),
    ._EVAL_22(bpu__EVAL_22),
    ._EVAL_23(bpu__EVAL_23),
    ._EVAL_24(bpu__EVAL_24),
    ._EVAL_25(bpu__EVAL_25),
    ._EVAL_26(bpu__EVAL_26),
    ._EVAL_27(bpu__EVAL_27),
    ._EVAL_28(bpu__EVAL_28),
    ._EVAL_29(bpu__EVAL_29),
    ._EVAL_30(bpu__EVAL_30),
    ._EVAL_31(bpu__EVAL_31),
    ._EVAL_32(bpu__EVAL_32),
    ._EVAL_33(bpu__EVAL_33),
    ._EVAL_34(bpu__EVAL_34),
    ._EVAL_35(bpu__EVAL_35),
    ._EVAL_36(bpu__EVAL_36),
    ._EVAL_37(bpu__EVAL_37),
    ._EVAL_38(bpu__EVAL_38),
    ._EVAL_39(bpu__EVAL_39),
    ._EVAL_40(bpu__EVAL_40),
    ._EVAL_41(bpu__EVAL_41),
    ._EVAL_42(bpu__EVAL_42),
    ._EVAL_43(bpu__EVAL_43)
  );
  _EVAL_155 rf (
    ._EVAL(rf__EVAL),
    ._EVAL_0(rf__EVAL_0),
    ._EVAL_1(rf__EVAL_1),
    ._EVAL_2(rf__EVAL_2),
    ._EVAL_3(rf__EVAL_3),
    ._EVAL_4(rf__EVAL_4),
    ._EVAL_5(rf__EVAL_5),
    ._EVAL_6(rf__EVAL_6)
  );
  _EVAL_153 alu (
    ._EVAL(alu__EVAL),
    ._EVAL_0(alu__EVAL_0),
    ._EVAL_1(alu__EVAL_1),
    ._EVAL_2(alu__EVAL_2),
    ._EVAL_3(alu__EVAL_3)
  );
  _EVAL_151 fetch (
    ._EVAL(fetch__EVAL),
    ._EVAL_0(fetch__EVAL_0),
    ._EVAL_1(fetch__EVAL_1),
    ._EVAL_2(fetch__EVAL_2),
    ._EVAL_3(fetch__EVAL_3),
    ._EVAL_4(fetch__EVAL_4),
    ._EVAL_5(fetch__EVAL_5),
    ._EVAL_6(fetch__EVAL_6),
    ._EVAL_7(fetch__EVAL_7),
    ._EVAL_8(fetch__EVAL_8),
    ._EVAL_9(fetch__EVAL_9),
    ._EVAL_10(fetch__EVAL_10),
    ._EVAL_11(fetch__EVAL_11),
    ._EVAL_12(fetch__EVAL_12),
    ._EVAL_13(fetch__EVAL_13),
    ._EVAL_14(fetch__EVAL_14),
    ._EVAL_15(fetch__EVAL_15),
    ._EVAL_16(fetch__EVAL_16),
    ._EVAL_17(fetch__EVAL_17),
    ._EVAL_18(fetch__EVAL_18),
    ._EVAL_19(fetch__EVAL_19),
    ._EVAL_20(fetch__EVAL_20),
    ._EVAL_21(fetch__EVAL_21),
    ._EVAL_22(fetch__EVAL_22),
    ._EVAL_23(fetch__EVAL_23)
  );
  _EVAL_156 pmp_checker (
    ._EVAL(pmp_checker__EVAL),
    ._EVAL_0(pmp_checker__EVAL_0),
    ._EVAL_1(pmp_checker__EVAL_1),
    ._EVAL_2(pmp_checker__EVAL_2),
    ._EVAL_3(pmp_checker__EVAL_3),
    ._EVAL_4(pmp_checker__EVAL_4),
    ._EVAL_5(pmp_checker__EVAL_5),
    ._EVAL_6(pmp_checker__EVAL_6),
    ._EVAL_7(pmp_checker__EVAL_7),
    ._EVAL_8(pmp_checker__EVAL_8),
    ._EVAL_9(pmp_checker__EVAL_9),
    ._EVAL_10(pmp_checker__EVAL_10),
    ._EVAL_11(pmp_checker__EVAL_11),
    ._EVAL_12(pmp_checker__EVAL_12),
    ._EVAL_13(pmp_checker__EVAL_13),
    ._EVAL_14(pmp_checker__EVAL_14),
    ._EVAL_15(pmp_checker__EVAL_15),
    ._EVAL_16(pmp_checker__EVAL_16),
    ._EVAL_17(pmp_checker__EVAL_17),
    ._EVAL_18(pmp_checker__EVAL_18),
    ._EVAL_19(pmp_checker__EVAL_19),
    ._EVAL_20(pmp_checker__EVAL_20),
    ._EVAL_21(pmp_checker__EVAL_21),
    ._EVAL_22(pmp_checker__EVAL_22),
    ._EVAL_23(pmp_checker__EVAL_23),
    ._EVAL_24(pmp_checker__EVAL_24),
    ._EVAL_25(pmp_checker__EVAL_25),
    ._EVAL_26(pmp_checker__EVAL_26),
    ._EVAL_27(pmp_checker__EVAL_27),
    ._EVAL_28(pmp_checker__EVAL_28),
    ._EVAL_29(pmp_checker__EVAL_29),
    ._EVAL_30(pmp_checker__EVAL_30),
    ._EVAL_31(pmp_checker__EVAL_31),
    ._EVAL_32(pmp_checker__EVAL_32),
    ._EVAL_33(pmp_checker__EVAL_33)
  );
  _EVAL_154 csr (
    ._EVAL(csr__EVAL),
    ._EVAL_0(csr__EVAL_0),
    ._EVAL_1(csr__EVAL_1),
    ._EVAL_2(csr__EVAL_2),
    ._EVAL_3(csr__EVAL_3),
    ._EVAL_4(csr__EVAL_4),
    ._EVAL_5(csr__EVAL_5),
    ._EVAL_6(csr__EVAL_6),
    ._EVAL_7(csr__EVAL_7),
    ._EVAL_8(csr__EVAL_8),
    ._EVAL_9(csr__EVAL_9),
    ._EVAL_10(csr__EVAL_10),
    ._EVAL_11(csr__EVAL_11),
    ._EVAL_12(csr__EVAL_12),
    ._EVAL_13(csr__EVAL_13),
    ._EVAL_14(csr__EVAL_14),
    ._EVAL_15(csr__EVAL_15),
    ._EVAL_16(csr__EVAL_16),
    ._EVAL_17(csr__EVAL_17),
    ._EVAL_18(csr__EVAL_18),
    ._EVAL_19(csr__EVAL_19),
    ._EVAL_20(csr__EVAL_20),
    ._EVAL_21(csr__EVAL_21),
    ._EVAL_22(csr__EVAL_22),
    ._EVAL_23(csr__EVAL_23),
    ._EVAL_24(csr__EVAL_24),
    ._EVAL_25(csr__EVAL_25),
    ._EVAL_26(csr__EVAL_26),
    ._EVAL_27(csr__EVAL_27),
    ._EVAL_28(csr__EVAL_28),
    ._EVAL_29(csr__EVAL_29),
    ._EVAL_30(csr__EVAL_30),
    ._EVAL_31(csr__EVAL_31),
    ._EVAL_32(csr__EVAL_32),
    ._EVAL_33(csr__EVAL_33),
    ._EVAL_34(csr__EVAL_34),
    ._EVAL_35(csr__EVAL_35),
    ._EVAL_36(csr__EVAL_36),
    ._EVAL_37(csr__EVAL_37),
    ._EVAL_38(csr__EVAL_38),
    ._EVAL_39(csr__EVAL_39),
    ._EVAL_40(csr__EVAL_40),
    ._EVAL_41(csr__EVAL_41),
    ._EVAL_42(csr__EVAL_42),
    ._EVAL_43(csr__EVAL_43),
    ._EVAL_44(csr__EVAL_44),
    ._EVAL_45(csr__EVAL_45),
    ._EVAL_46(csr__EVAL_46),
    ._EVAL_47(csr__EVAL_47),
    ._EVAL_48(csr__EVAL_48),
    ._EVAL_49(csr__EVAL_49),
    ._EVAL_50(csr__EVAL_50),
    ._EVAL_51(csr__EVAL_51),
    ._EVAL_52(csr__EVAL_52),
    ._EVAL_53(csr__EVAL_53),
    ._EVAL_54(csr__EVAL_54),
    ._EVAL_55(csr__EVAL_55),
    ._EVAL_56(csr__EVAL_56),
    ._EVAL_57(csr__EVAL_57),
    ._EVAL_58(csr__EVAL_58),
    ._EVAL_59(csr__EVAL_59),
    ._EVAL_60(csr__EVAL_60),
    ._EVAL_61(csr__EVAL_61),
    ._EVAL_62(csr__EVAL_62),
    ._EVAL_63(csr__EVAL_63),
    ._EVAL_64(csr__EVAL_64),
    ._EVAL_65(csr__EVAL_65),
    ._EVAL_66(csr__EVAL_66),
    ._EVAL_67(csr__EVAL_67),
    ._EVAL_68(csr__EVAL_68),
    ._EVAL_69(csr__EVAL_69),
    ._EVAL_70(csr__EVAL_70),
    ._EVAL_71(csr__EVAL_71),
    ._EVAL_72(csr__EVAL_72),
    ._EVAL_73(csr__EVAL_73),
    ._EVAL_74(csr__EVAL_74),
    ._EVAL_75(csr__EVAL_75),
    ._EVAL_76(csr__EVAL_76),
    ._EVAL_77(csr__EVAL_77),
    ._EVAL_78(csr__EVAL_78),
    ._EVAL_79(csr__EVAL_79),
    ._EVAL_80(csr__EVAL_80),
    ._EVAL_81(csr__EVAL_81),
    ._EVAL_82(csr__EVAL_82),
    ._EVAL_83(csr__EVAL_83),
    ._EVAL_84(csr__EVAL_84),
    ._EVAL_85(csr__EVAL_85),
    ._EVAL_86(csr__EVAL_86),
    ._EVAL_87(csr__EVAL_87),
    ._EVAL_88(csr__EVAL_88),
    ._EVAL_89(csr__EVAL_89),
    ._EVAL_90(csr__EVAL_90),
    ._EVAL_91(csr__EVAL_91),
    ._EVAL_92(csr__EVAL_92),
    ._EVAL_93(csr__EVAL_93),
    ._EVAL_94(csr__EVAL_94),
    ._EVAL_95(csr__EVAL_95),
    ._EVAL_96(csr__EVAL_96),
    ._EVAL_97(csr__EVAL_97),
    ._EVAL_98(csr__EVAL_98),
    ._EVAL_99(csr__EVAL_99),
    ._EVAL_100(csr__EVAL_100),
    ._EVAL_101(csr__EVAL_101),
    ._EVAL_102(csr__EVAL_102),
    ._EVAL_103(csr__EVAL_103),
    ._EVAL_104(csr__EVAL_104),
    ._EVAL_105(csr__EVAL_105),
    ._EVAL_106(csr__EVAL_106),
    ._EVAL_107(csr__EVAL_107),
    ._EVAL_108(csr__EVAL_108),
    ._EVAL_109(csr__EVAL_109),
    ._EVAL_110(csr__EVAL_110),
    ._EVAL_111(csr__EVAL_111),
    ._EVAL_112(csr__EVAL_112),
    ._EVAL_113(csr__EVAL_113),
    ._EVAL_114(csr__EVAL_114),
    ._EVAL_115(csr__EVAL_115),
    ._EVAL_116(csr__EVAL_116),
    ._EVAL_117(csr__EVAL_117),
    ._EVAL_118(csr__EVAL_118),
    ._EVAL_119(csr__EVAL_119),
    ._EVAL_120(csr__EVAL_120),
    ._EVAL_121(csr__EVAL_121),
    ._EVAL_122(csr__EVAL_122),
    ._EVAL_123(csr__EVAL_123),
    ._EVAL_124(csr__EVAL_124),
    ._EVAL_125(csr__EVAL_125),
    ._EVAL_126(csr__EVAL_126),
    ._EVAL_127(csr__EVAL_127),
    ._EVAL_128(csr__EVAL_128),
    ._EVAL_129(csr__EVAL_129),
    ._EVAL_130(csr__EVAL_130),
    ._EVAL_131(csr__EVAL_131),
    ._EVAL_132(csr__EVAL_132),
    ._EVAL_133(csr__EVAL_133),
    ._EVAL_134(csr__EVAL_134),
    ._EVAL_135(csr__EVAL_135),
    ._EVAL_136(csr__EVAL_136),
    ._EVAL_137(csr__EVAL_137),
    ._EVAL_138(csr__EVAL_138),
    ._EVAL_139(csr__EVAL_139),
    ._EVAL_140(csr__EVAL_140),
    ._EVAL_141(csr__EVAL_141)
  );
  _EVAL_152 div (
    ._EVAL(div__EVAL),
    ._EVAL_0(div__EVAL_0),
    ._EVAL_1(div__EVAL_1),
    ._EVAL_2(div__EVAL_2),
    ._EVAL_3(div__EVAL_3),
    ._EVAL_4(div__EVAL_4),
    ._EVAL_5(div__EVAL_5),
    ._EVAL_6(div__EVAL_6),
    ._EVAL_7(div__EVAL_7),
    ._EVAL_8(div__EVAL_8)
  );
  assign _EVAL_17543 = _EVAL_8865 | _EVAL_974;
  assign _EVAL_8013 = 32'h1073 == _EVAL_1530;
  assign _EVAL_805 = _EVAL_11480 & 32'h40003014;
  assign _EVAL_4323 = _EVAL_29;
  assign _EVAL_636 = fetch__EVAL & _EVAL_2953;
  assign _EVAL_1606 = _EVAL_15759 ? _EVAL_3051 : _EVAL_8128;
  assign _EVAL_10114 = _EVAL_10368 | _EVAL_11801;
  assign _EVAL_1988 = _EVAL_11480 & 32'h18;
  assign _EVAL_10588 = _EVAL_11480 & 32'h2050;
  assign _EVAL_6556 = _EVAL_10919 | _EVAL_9896;
  assign _EVAL_8339 = _EVAL_3611 & _EVAL_18675;
  assign _EVAL_4897 = _EVAL_12724;
  assign _EVAL_18675 = _EVAL_9491 | csr__EVAL_49;
  assign _EVAL_16200 = 32'h37 == _EVAL_6918;
  assign div__EVAL_5 = _EVAL_64;
  assign _EVAL_11613 = $signed(_EVAL_11503) == 33'sh0;
  assign _EVAL_6265 = _EVAL_11480[26];
  assign _EVAL_5648 = _EVAL_6884 & _EVAL_3741;
  assign _EVAL_15596 = 32'h1023 == _EVAL_1530;
  assign _EVAL_5883 = _EVAL_10782 | _EVAL_12623;
  assign _EVAL_13198 = _EVAL_6422 & _EVAL_16024;
  assign _EVAL_1027 = _EVAL_12043 ? _EVAL_9768 : _EVAL_14765;
  assign _EVAL_9061 = _EVAL_8706 & _EVAL_13130;
  assign _EVAL_11919 = _EVAL_9300 | _EVAL_17383;
  assign _EVAL_6945 = _EVAL_15785 ^ 32'h3000;
  assign _EVAL_13053 = 1'h0;
  assign _EVAL_15219 = ~_EVAL_1128;
  assign fetch_pmp_checker__EVAL_13 = csr__EVAL_110;
  assign _EVAL_5589 = _EVAL_14011 | _EVAL_11613;
  assign _EVAL_10566 = 32'hc000202f == _EVAL_12083;
  assign _EVAL_14804 = _EVAL_9187 ? 3'h0 : _EVAL_10692;
  assign _EVAL_19347 = _EVAL_12263 | _EVAL_2458;
  assign _EVAL_15156 = _EVAL_16096 | _EVAL_17570;
  assign fetch_pmp_checker__EVAL_20 = csr__EVAL_127;
  assign pmp_checker__EVAL_10 = csr__EVAL_25;
  assign fetch_pmp_checker__EVAL_7 = csr__EVAL_60;
  assign _EVAL_9545 = _EVAL_10588 == 32'h2000;
  assign _EVAL_14142 = _EVAL_2109 & pmp_checker__EVAL_4;
  assign _EVAL_13006 = {{31'd0}, _EVAL_13};
  assign _EVAL_12823 = _EVAL_9843 ^ 32'h3000;
  assign _EVAL_3930 = fetch__EVAL & _EVAL_7638;
  assign _EVAL_1627 = 32'h40005013 == _EVAL_12413;
  assign _EVAL_14573 = _EVAL_16872 | _EVAL_12352;
  assign _EVAL_6706 = _EVAL_2871 | _EVAL_15511;
  assign _EVAL_17967 = _EVAL_2277 & _EVAL_12356;
  assign _EVAL_11701 = _EVAL_16096 & _EVAL_10735;
  assign _EVAL_11868 = $signed(_EVAL_14115) & -33'sh2000;
  assign _EVAL_15398 = _EVAL_7616 | _EVAL_17384;
  assign _EVAL_2373 = _EVAL_12957;
  assign _EVAL_9667 = _EVAL_3248 | _EVAL_437;
  assign _EVAL_5412 = _EVAL_6789 ? 1'h0 : _EVAL_5564;
  assign _EVAL_58 = _EVAL_17997;
  assign _EVAL_11654 = _EVAL_13703 & _EVAL_8336;
  assign _EVAL_17033 = _EVAL_15785 ^ 32'h40000000;
  assign _EVAL_18765 = _EVAL_4888;
  assign _EVAL_12967 = _EVAL_13099 & _EVAL_15106;
  assign fetch_pmp_checker__EVAL_18 = csr__EVAL_114;
  assign _EVAL_22 = _EVAL_3607;
  assign _EVAL_9843 = _EVAL_6756[31:0];
  assign _EVAL_6770 = 32'h202f == _EVAL_12083;
  assign csr__EVAL_113 = _EVAL_8;
  assign _EVAL_17688 = _EVAL_18765;
  assign _EVAL_16668 = _EVAL_11162 & _EVAL_12379;
  assign _EVAL_18361 = ~_EVAL_3130;
  assign _EVAL_11503 = _EVAL_7378;
  assign _EVAL_19458 = ~_EVAL_9449;
  assign _EVAL_16323 = _EVAL_6548 | _EVAL_19509;
  assign _EVAL_6767 = 32'h8000202f == _EVAL_12083;
  assign _EVAL_13735 = _EVAL_11480[30:25];
  assign _EVAL_17640 = _EVAL_6156 | _EVAL_16202;
  assign rf__EVAL_4 = _EVAL_3139 ? 1'h0 : _EVAL_15156;
  assign _EVAL_6336 = 32'h7063 == _EVAL_1530;
  assign _EVAL_15974 = _EVAL_16201 & _EVAL_1478;
  assign _EVAL_9583 = ~_EVAL_9364;
  assign _EVAL_19611 = _EVAL_11480 & 32'h2010;
  assign _EVAL_11712 = 3'h0;
  assign _EVAL_10207 = 32'hf == _EVAL_1530;
  assign _EVAL_11716 = fetch__EVAL & _EVAL_17854;
  assign _EVAL_15976 = _EVAL_9496 | _EVAL_11046;
  assign _EVAL_17352 = $signed(_EVAL_4646) == 33'sh0;
  assign _EVAL_13761 = _EVAL_15785 ^ 32'h20000000;
  assign _EVAL_8112 = _EVAL_4380 | _EVAL_15801;
  assign _EVAL_15106 = _EVAL_11480[25];
  assign _EVAL_3302 = {1'h1,_EVAL_5907,_EVAL_14763};
  assign _EVAL_12829 = {_EVAL_11557,_EVAL_18613};
  assign _EVAL_8873 = _EVAL_11858 | _EVAL_6533;
  assign bpu__EVAL_27 = csr__EVAL_24;
  assign _EVAL_12568 = _EVAL_3816 & _EVAL_5146;
  assign _EVAL_10553 = _EVAL_11716 ? 3'h0 : 3'h4;
  assign _EVAL_9066 = _EVAL_2508 | _EVAL_16392;
  assign pmp_checker__EVAL_29 = csr__EVAL_54;
  assign _EVAL_16202 = _EVAL_14257 == 32'h40000030;
  assign _EVAL_11005 = 32'h6f == _EVAL_6918;
  assign bpu__EVAL_32 = csr__EVAL_80;
  assign div__EVAL_7 = _EVAL_2743 ? _EVAL_16768 : _EVAL_17404;
  assign _EVAL_16593 = _EVAL_8631;
  assign _EVAL_15648 = _EVAL_4267 != 24'h0;
  assign _EVAL_11531 = _EVAL_7414 == 32'h0;
  assign _EVAL_18990 = _EVAL_16096 & _EVAL_18361;
  assign _EVAL_17887 = _EVAL_15759 | _EVAL_17934;
  assign _EVAL_15427 = _EVAL_15097 == 2'h0;
  assign _EVAL_13133 = _EVAL_7880[3:0];
  assign pmp_checker__EVAL_18 = csr__EVAL_114;
  assign _EVAL_9086 = fetch__EVAL & _EVAL_18360;
  assign _EVAL_17074 = ~_EVAL_15890;
  assign _EVAL_49 = _EVAL_15396;
  assign _EVAL_56 = _EVAL_13072;
  assign bpu__EVAL_37 = csr__EVAL_119;
  assign fetch_pmp_checker__EVAL_21 = csr__EVAL_57;
  assign fetch_pmp_checker__EVAL_28 = _EVAL_64;
  assign fetch_pmp_checker__EVAL_26 = csr__EVAL_29;
  assign _EVAL_11218 = _EVAL_15759 ? _EVAL_16733 : _EVAL_17801;
  assign _EVAL_12682 = _EVAL_10181 | _EVAL_2629;
  assign _EVAL_9514 = ~_EVAL_14478;
  assign _EVAL_19285 = _EVAL_11480[11:8];
  assign _EVAL_15242 = _EVAL_10825 & _EVAL_8178;
  assign _EVAL_2293 = 32'h6013 == _EVAL_1530;
  assign _EVAL_4545 = 32'h67 == _EVAL_1530;
  assign csr__EVAL_98 = _EVAL_92 & _EVAL_19408;
  assign _EVAL_7616 = _EVAL_3775 | _EVAL_3102;
  assign _EVAL_5332 = _EVAL_19208 | _EVAL_2080;
  assign _EVAL_16448 = _EVAL_2558 | _EVAL_1546;
  assign _EVAL_6252 = _EVAL_10778 & _EVAL_10735;
  assign _EVAL_4042 = {1'b0,$signed(_EVAL_9820)};
  assign bpu__EVAL_43 = csr__EVAL_140;
  assign _EVAL_1962 = _EVAL_13609 | _EVAL_2644;
  assign _EVAL_4646 = _EVAL_9314;
  assign _EVAL_12477 = _EVAL_10831 & _EVAL_7638;
  assign _EVAL_11533 = _EVAL_1437 ? 3'h0 : 3'h4;
  assign pmp_checker__EVAL_19 = csr__EVAL_5;
  assign alu__EVAL_0 = _EVAL_15398 | _EVAL_4045;
  assign _EVAL_6918 = _EVAL_11480 & 32'h7f;
  assign _EVAL_12247 = _EVAL_14478 | _EVAL_15003;
  assign _EVAL_11838 = ~_EVAL_15759;
  assign bpu__EVAL_11 = csr__EVAL_13;
  assign _EVAL_10831 = _EVAL_1636 & _EVAL_2139;
  assign _EVAL_5341 = ~_EVAL_9843;
  assign _EVAL_8958 = _EVAL_14722 == 32'h1008;
  assign _EVAL_1995 = _EVAL_1801 ? _EVAL_6647 : _EVAL_12379;
  assign _EVAL_5009 = _EVAL_5171;
  assign _EVAL_15131 = _EVAL_11480 & 32'h48;
  assign _EVAL_18642 = _EVAL_4027 | _EVAL_6286;
  assign _EVAL_10147 = ~div__EVAL_3;
  assign _EVAL_17584 = _EVAL_14478 ? _EVAL_12498 : fetch__EVAL_20;
  assign csr__EVAL = _EVAL_10831 & _EVAL_7638;
  assign _EVAL_151 = csr__EVAL_101[7:5];
  assign _EVAL_4660 = _EVAL_8958 | _EVAL_12967;
  assign _EVAL_12216 = 32'h4000202f == _EVAL_12083;
  assign _EVAL_17194 = _EVAL_8999 & _EVAL_14160;
  assign _EVAL_4469 = _EVAL_6706 | _EVAL_1860;
  assign _EVAL_10692 = _EVAL_5726 ? 3'h2 : 3'h1;
  assign _EVAL_5138 = {_EVAL_2373,_EVAL_5960,_EVAL_5009,_EVAL_2373,_EVAL_13735,_EVAL_16395,_EVAL_4888};
  assign _EVAL_8522 = _EVAL_11900;
  assign _EVAL_11230 = _EVAL_14765[15:0];
  assign _EVAL_7638 = ~_EVAL_7993;
  assign _EVAL_2258 = _EVAL_8999 & _EVAL_6647;
  assign _EVAL_11504 = _EVAL_11480[12];
  assign _EVAL_2845 = {21'h0,6'h0,_EVAL_1503,_EVAL_6492};
  assign fetch_pmp_checker__EVAL_30 = csr__EVAL_89;
  assign _EVAL_44 = _EVAL_16649;
  assign _EVAL_16395 = _EVAL_11480[24:21];
  assign _EVAL_8116 = 32'h7b200073 == _EVAL_11480;
  assign _EVAL_13772 = ~_EVAL_10181;
  assign fetch__EVAL_19 = _EVAL_10831 & _EVAL_12589;
  assign _EVAL_5962 = _EVAL_1636 & _EVAL_12247;
  assign _EVAL_12360 = _EVAL_6101;
  assign _EVAL_3121 = 1'h1;
  assign _EVAL_19408 = ~_EVAL_11533;
  assign _EVAL_17953 = _EVAL_5684 | _EVAL_16592;
  assign _EVAL_17740 = _EVAL_11189 == 32'h2008;
  assign _EVAL_14680 = _EVAL_573 ? 1'h0 : _EVAL_14478;
  assign pmp_checker__EVAL_7 = csr__EVAL_60;
  assign _EVAL_272 = _EVAL_11480 & 32'hc;
  assign _EVAL_11521 = 32'h10500073 == _EVAL_11480;
  assign _EVAL_8228 = _EVAL_11480 & 32'h34;
  assign _EVAL_2593 = 1'h0;
  assign _EVAL_16201 = _EVAL_1801 ? _EVAL_12371 : _EVAL_9510;
  assign _EVAL_11458 = _EVAL_272 == 32'h4;
  assign _EVAL_14969 = _EVAL_36;
  assign pmp_checker__EVAL_26 = csr__EVAL_29;
  assign _EVAL_41 = _EVAL_3858;
  assign _EVAL_4830 = _EVAL_14356;
  assign csr__EVAL_3 = _EVAL_2653;
  assign _EVAL_19297 = _EVAL;
  assign _EVAL_4361 = _EVAL_10331 == 32'h4;
  assign rf__EVAL_1 = _EVAL_3139 ? 5'h0 : _EVAL_15219;
  assign _EVAL_9169 = {{27'd0}, fetch__EVAL_17};
  assign _EVAL_7809 = _EVAL_13327 & _EVAL_2125;
  assign _EVAL_12545 = _EVAL_151 == 3'h5;
  assign _EVAL_14814 = $signed(_EVAL_8912) & -33'sh1000;
  assign _EVAL_6449 = _EVAL_17963 | _EVAL_6336;
  assign _EVAL_3500 = _EVAL_1801 ? _EVAL_8874 : _EVAL_12508;
  assign _EVAL_8584 = _EVAL_2832 != 32'h0;
  assign _EVAL_14107 = _EVAL_14356;
  assign pmp_checker__EVAL_23 = csr__EVAL_49 ? csr__EVAL_1 : csr__EVAL_129;
  assign _EVAL_13371 = _EVAL_55;
  assign _EVAL_12282 = _EVAL_14448 ? _EVAL_15910 : _EVAL_12521;
  assign _EVAL_17140 = _EVAL_5907 & _EVAL_15479;
  assign fetch_pmp_checker__EVAL_14 = csr__EVAL_46;
  assign _EVAL_13210 = _EVAL_3495 | bpu__EVAL_34;
  assign _EVAL_7993 = _EVAL_17821;
  assign _EVAL_5387 = _EVAL_4937 | _EVAL_19297;
  assign _EVAL_19059 = _EVAL_6530;
  assign csr__EVAL_108 = _EVAL_19273;
  assign _EVAL_10239 = _EVAL_3930 & _EVAL_8627;
  assign _EVAL_18216 = _EVAL_14896 == _EVAL_15591;
  assign _EVAL_4450 = _EVAL_13703 ? 32'h3 : 32'h0;
  assign _EVAL_15910 = $signed(_EVAL_12611) < $signed(_EVAL_19337);
  assign _EVAL_4191 = {1'b0,$signed(_EVAL_12823)};
  assign bpu__EVAL_5 = csr__EVAL_9;
  assign _EVAL_14832 = _EVAL_10114 | _EVAL_17447;
  assign bpu__EVAL_9 = csr__EVAL_141;
  assign div__EVAL_0 = _EVAL_6270 ? _EVAL_16768 : _EVAL_7879;
  assign _EVAL_14448 = _EVAL_11480[14];
  assign _EVAL_19413 = _EVAL_10284 | _EVAL_14159;
  assign _EVAL_1530 = _EVAL_11480 & 32'h707f;
  assign _EVAL_5512 = _EVAL_4216 & _EVAL_19458;
  assign _EVAL_2238 = _EVAL_9066 | _EVAL_11311;
  assign _EVAL_2483 = _EVAL_7743 | _EVAL_4521;
  assign _EVAL_5066 = 32'h6033 == _EVAL_12413;
  assign _EVAL_18912 = $signed(_EVAL_18960) == 33'sh0;
  assign _EVAL_16024 = _EVAL_11504 ^ _EVAL_12282;
  assign _EVAL_16483 = _EVAL_61;
  assign _EVAL_2727 = _EVAL_5908;
  assign bpu__EVAL_17 = csr__EVAL_123;
  assign _EVAL_9941 = _EVAL_13371 & _EVAL_15981;
  assign _EVAL_16392 = 32'h63 == _EVAL_1530;
  assign bpu__EVAL_4 = csr__EVAL_45;
  assign fetch__EVAL_10 = ~_EVAL_18258;
  assign _EVAL_1640 = 32'h800202f == _EVAL_12083;
  assign fetch__EVAL_13 = _EVAL_6756[31:0];
  assign _EVAL_8412 = _EVAL_2895 & _EVAL_14142;
  assign _EVAL_5001 = _EVAL_9556 ? _EVAL_16227 : 3'h0;
  assign _EVAL_17447 = 32'h2013 == _EVAL_1530;
  assign _EVAL_8051 = _EVAL_5726 ? 3'h1 : 3'h0;
  assign _EVAL_642 = _EVAL_11480 & 32'h70;
  assign _EVAL_46 = _EVAL_16649;
  assign _EVAL_5726 = _EVAL_11480[29];
  assign _EVAL_1745 = {_EVAL_7201,_EVAL_5728};
  assign _EVAL_779 = 32'h0;
  assign _EVAL_13045 = _EVAL_3495 ? csr__EVAL_37 : {{28'd0}, _EVAL_13825};
  assign _EVAL_15968 = _EVAL_2058 ? _EVAL_6261 : _EVAL_11436;
  assign _EVAL_10289 = _EVAL_19347 | _EVAL_8116;
  assign _EVAL_9689 = _EVAL_4218 | _EVAL_4189;
  assign _EVAL_18202 = _EVAL_2761 & csr__EVAL_72;
  assign bpu__EVAL_25 = csr__EVAL_136;
  assign _EVAL_15409 = _EVAL_14092 | _EVAL_2638;
  assign _EVAL_8187 = _EVAL_3993;
  assign _EVAL_284 = 32'h30500073 == _EVAL_11480;
  assign _EVAL_16722 = 1'h0;
  assign bpu__EVAL_39 = csr__EVAL_116;
  assign _EVAL_4292 = _EVAL_2751 == _EVAL_10383;
  assign _EVAL_2900 = _EVAL_11251 ? 2'h2 : 2'h0;
  assign _EVAL_4257 = _EVAL_17953 | _EVAL_19610;
  assign _EVAL_2492 = _EVAL_4297 == _EVAL_10383;
  assign _EVAL_10284 = _EVAL_17909 == 32'h4;
  assign _EVAL_9378 = _EVAL_17570 & _EVAL_16096;
  assign _EVAL_1128 = _EVAL_17570 ? _EVAL_5671 : _EVAL_14896;
  assign fetch_pmp_checker__EVAL_33 = csr__EVAL_14;
  assign _EVAL_16649 = 1'h0;
  assign _EVAL_5049 = _EVAL_8865 & csr__EVAL_70;
  assign _EVAL_39 = _EVAL_15768;
  assign _EVAL_8864 = _EVAL_2258 & _EVAL_4292;
  assign _EVAL_9300 = _EVAL_18449 | _EVAL_18119;
  assign _EVAL_10181 = _EVAL_11480[31];
  assign _EVAL_8312 = _EVAL_7993 ? _EVAL_897 : _EVAL_5227;
  assign _EVAL_3442 = _EVAL_5564 & _EVAL_9364;
  assign _EVAL_9472 = _EVAL_15765 == 32'h10;
  assign _EVAL_15340 = $signed(_EVAL_427) == 33'sh0;
  assign _EVAL_3852 = _EVAL_13170 == 32'h2010;
  assign _EVAL_10825 = _EVAL_11596 & _EVAL_8627;
  assign _EVAL_6196 = _EVAL_12682 ? _EVAL_16323 : _EVAL_16323;
  assign _EVAL_12476 = _EVAL_15097 >= 2'h1;
  assign _EVAL_2740 = _EVAL_9464 ? _EVAL_12411 : 32'h0;
  assign _EVAL_4798 = _EVAL_13007;
  assign _EVAL_2058 = _EVAL_13287[0];
  assign csr__EVAL_6 = _EVAL_10148;
  assign _EVAL_319 = ~_EVAL_11531;
  assign _EVAL_8163 = _EVAL_8137 & _EVAL_2483;
  assign _EVAL_12043 = _EVAL_15097 == 2'h1;
  assign _EVAL_2953 = _EVAL_8872 | _EVAL_4361;
  assign _EVAL_14231 = _EVAL_15242 & fetch__EVAL_22;
  assign _EVAL_5381 = _EVAL_9378 & _EVAL_4213;
  assign csr__EVAL_61 = _EVAL_18514;
  assign _EVAL_12887 = _EVAL_19597 & _EVAL_13129;
  assign _EVAL_3775 = _EVAL_14573 | _EVAL_4030;
  assign _EVAL_17546 = _EVAL_5162 ? _EVAL_1745 : 2'h0;
  assign _EVAL_2265 = 3'h0;
  assign _EVAL_11356 = _EVAL_10148[31:16];
  assign bpu__EVAL_3 = csr__EVAL_32;
  assign _EVAL_12651 = {_EVAL_2373,_EVAL_9697,_EVAL_12793,1'h0,11'h0};
  assign _EVAL_857 = 3'h4;
  assign _EVAL_9039 = _EVAL_3444 ? alu__EVAL_3 : 32'h0;
  assign fetch_pmp_checker__EVAL_11 = csr__EVAL_41;
  assign _EVAL_11557 = _EVAL_17546 | _EVAL_12376;
  assign _EVAL_10896 = _EVAL_47;
  assign pmp_checker__EVAL_5 = csr__EVAL_77;
  assign _EVAL_12427 = _EVAL_8607 | _EVAL_6770;
  assign _EVAL_13253 = _EVAL_10831 & _EVAL_6422;
  assign _EVAL_18960 = _EVAL_7679;
  assign _EVAL_11436 = _EVAL_5612[7:0];
  assign _EVAL_2895 = csr__EVAL_49 & _EVAL_14355;
  assign _EVAL_13835 = _EVAL_15759 ? _EVAL_10468 : _EVAL_5346;
  assign _EVAL_8621 = _EVAL_17356 | _EVAL_11278;
  assign _EVAL_7487 = _EVAL_4376 | _EVAL_12096;
  assign _EVAL_3320 = _EVAL_16620 == 32'h1010;
  assign _EVAL_17093 = _EVAL_14051 ? _EVAL_10491 : _EVAL_11356;
  assign _EVAL_6261 = _EVAL_5612[15:8];
  assign _EVAL_15504 = _EVAL_11480 & 32'h2048;
  assign _EVAL_15418 = {11{_EVAL_12957}};
  assign _EVAL_7897 = _EVAL_17;
  assign _EVAL_14251 = _EVAL_16377;
  assign fetch__EVAL_14 = _EVAL_4323;
  assign _EVAL_10233 = ~_EVAL_11654;
  assign _EVAL_4381 = _EVAL_4753 | _EVAL_9411;
  assign _EVAL_17736 = _EVAL_16768;
  assign pmp_checker__EVAL_3 = csr__EVAL_115;
  assign _EVAL_9314 = $signed(_EVAL_12339) & -33'sh1000;
  assign _EVAL_12850 = _EVAL_1389 | _EVAL_8070;
  assign _EVAL_12525 = _EVAL_15890 ? 3'h3 : _EVAL_14804;
  assign _EVAL_13287 = _EVAL_1801 ? _EVAL_19551 : _EVAL_5900;
  assign _EVAL_703 = _EVAL_11607 == 32'h2000030;
  assign _EVAL_11561 = _EVAL_6538;
  assign _EVAL_10735 = _EVAL_10383 != 5'h0;
  assign _EVAL_12244 = 4'hf;
  assign _EVAL_3820 = _EVAL_19144 | _EVAL_5301;
  assign _EVAL_10012 = _EVAL_15526 | _EVAL_4446;
  assign _EVAL_5908 = $signed(_EVAL_13694) & -33'sh1000000;
  assign _EVAL_8912 = {1'b0,$signed(_EVAL_9843)};
  assign _EVAL_12112 = _EVAL_8580;
  assign _EVAL_17909 = _EVAL_11480 & 32'h2c;
  assign _EVAL_9896 = _EVAL_703 & _EVAL_13139;
  assign _EVAL_18119 = 32'h33 == _EVAL_12413;
  assign _EVAL_12438 = _EVAL_12682 ? 2'h2 : 2'h3;
  assign _EVAL_18360 = ~_EVAL_18258;
  assign _EVAL_4376 = _EVAL_8621 | _EVAL_16034;
  assign _EVAL_16592 = _EVAL_8646 == 32'h20;
  assign _EVAL_14263 = {1'b0,$signed(_EVAL_4663)};
  assign _EVAL_14196 = _EVAL_14;
  assign _EVAL_17589 = _EVAL_7809;
  assign _EVAL_1389 = _EVAL_3623 | _EVAL_10207;
  assign _EVAL_4446 = 32'h6000202f == _EVAL_12083;
  assign _EVAL_10622 = _EVAL_2793 == 32'h0;
  assign _EVAL_3 = _EVAL_10371;
  assign _EVAL_15382 = _EVAL_11838 & _EVAL_14355;
  assign _EVAL_573 = _EVAL_6951 & _EVAL_3858;
  assign _EVAL_16796 = _EVAL_1636 & _EVAL_9514;
  assign _EVAL_9187 = ~_EVAL_8899;
  assign _EVAL_12981 = _EVAL_4469 | _EVAL_11178;
  assign _EVAL_17854 = _EVAL_3045 == 32'h20;
  assign _EVAL_1983 = $signed(_EVAL_8522) == 33'sh0;
  assign _EVAL_16877 = _EVAL_16407 & _EVAL_12545;
  assign _EVAL_16288 = _EVAL_11480 & 32'h4004;
  assign _EVAL_6 = _EVAL_6400;
  assign _EVAL_17560 = _EVAL_16164 ? _EVAL_15785 : _EVAL_9843;
  assign _EVAL_4619 = 32'h2023 == _EVAL_1530;
  assign _EVAL_4380 = _EVAL_5332 | _EVAL_4295;
  assign _EVAL_9965 = _EVAL_13099 & _EVAL_6265;
  assign pmp_checker__EVAL_21 = csr__EVAL_57;
  assign _EVAL_18078 = _EVAL_4834;
  assign _EVAL_10019 = _EVAL_14814;
  assign _EVAL_6214 = $signed(_EVAL_14263) & -33'sh1000;
  assign _EVAL_1478 = _EVAL_15968[7];
  assign _EVAL_7743 = _EVAL_16668 & _EVAL_2446;
  assign _EVAL_8892 = _EVAL_15591 == 5'h0;
  assign _EVAL_2225 = _EVAL_10831 & _EVAL_8312;
  assign _EVAL_6719 = _EVAL_703 & _EVAL_15184;
  assign _EVAL_15272 = _EVAL_17995 | _EVAL_8112;
  assign _EVAL_1546 = 32'h7033 == _EVAL_12413;
  assign _EVAL_8990 = fetch__EVAL & _EVAL_5566;
  assign _EVAL_7366 = _EVAL_14765[31];
  assign _EVAL_6328 = _EVAL_6586 == 32'h10;
  assign _EVAL_11252 = fetch__EVAL_11[15:0];
  assign _EVAL_5671 = _EVAL_1801 ? _EVAL_2751 : _EVAL_4297;
  assign csr__EVAL_0 = _EVAL_20;
  assign _EVAL_16898 = csr__EVAL_4[31:8];
  assign _EVAL_6101 = _EVAL_12651;
  assign _EVAL_3330 = _EVAL_11480 & 32'h1050;
  assign _EVAL_12601 = _EVAL_12477 & _EVAL_13977;
  assign _EVAL_12263 = _EVAL_2198 | _EVAL_13586;
  assign _EVAL_14355 = ~_EVAL_11178;
  assign bpu__EVAL_8 = csr__EVAL_90;
  assign _EVAL_17283 = _EVAL_13371 & _EVAL_3500;
  assign _EVAL_935 = _EVAL_9700 & _EVAL_4213;
  assign _EVAL_17986 = _EVAL_1067 | _EVAL_2488;
  assign _EVAL_4 = _EVAL_16649;
  assign _EVAL_8195 = 32'h5033 == _EVAL_12413;
  assign _EVAL_1969 = _EVAL_6556 | _EVAL_9364;
  assign _EVAL_14726 = 1'h0;
  assign _EVAL_12376 = _EVAL_19430 ? 2'h3 : 2'h0;
  assign _EVAL_1297 = _EVAL_11919 | _EVAL_8702;
  assign _EVAL_11801 = 32'h13 == _EVAL_1530;
  assign _EVAL_3878 = _EVAL_17583 | _EVAL_9472;
  assign _EVAL_409 = 32'h2002033 == _EVAL_12413;
  assign _EVAL_10919 = _EVAL_706 | _EVAL_6328;
  assign _EVAL_16380 = _EVAL_14809 | _EVAL_16256;
  assign _EVAL_6057 = 1'h1;
  assign _EVAL_413 = _EVAL_6765 == 32'h0;
  assign _EVAL_10948 = _EVAL_15553 | _EVAL_869;
  assign _EVAL_15526 = _EVAL_11875 | _EVAL_1640;
  assign _EVAL_6053 = _EVAL_13772 ? 3'h4 : _EVAL_17519;
  assign _EVAL_13298 = _EVAL_13687 == 32'h8;
  assign bpu__EVAL_24 = csr__EVAL_88;
  assign _EVAL_909 = _EVAL_3878 | _EVAL_8872;
  assign _EVAL_54 = _EVAL_16543;
  assign _EVAL_5346 = csr__EVAL_129 == 2'h3;
  assign _EVAL_952 = _EVAL_6840 | _EVAL_3448;
  assign _EVAL_12010 = _EVAL_15112 & _EVAL_5566;
  assign _EVAL_13047 = _EVAL_12601 & _EVAL_13304;
  assign _EVAL_2653 = 2'h3;
  assign csr__EVAL_93 = _EVAL_10831 & _EVAL_7993;
  assign _EVAL_974 = _EVAL_2761 & _EVAL_16877;
  assign pmp_checker__EVAL_12 = csr__EVAL_133;
  assign _EVAL_8646 = _EVAL_11480 & 32'h64;
  assign _EVAL_13139 = ~_EVAL_14448;
  assign _EVAL_4709 = _EVAL_12411 + _EVAL_16060;
  assign bpu__EVAL_28 = csr__EVAL_100;
  assign _EVAL_19578 = alu__EVAL_2[0];
  assign _EVAL_19430 = _EVAL_15097 >= 2'h2;
  assign _EVAL_7053 = _EVAL_16096 & _EVAL_7194;
  assign _EVAL_8148 = _EVAL_5907 & bpu__EVAL_36;
  assign _EVAL_9464 = _EVAL_19413 | _EVAL_8872;
  assign _EVAL_18289 = _EVAL_14183 == 32'h2000030;
  assign _EVAL_10 = _EVAL_16649;
  assign _EVAL_13170 = _EVAL_11480 & 32'h2006014;
  assign _EVAL_13158 = _EVAL_9277;
  assign _EVAL_17254 = _EVAL_17352 | _EVAL_7502;
  assign bpu__EVAL_10 = csr__EVAL_138;
  assign pmp_checker__EVAL_28 = _EVAL_64;
  assign _EVAL_3593 = 32'h2000202f == _EVAL_12083;
  assign _EVAL_26 = _EVAL_19090;
  assign fetch_pmp_checker__EVAL = _EVAL_36;
  assign _EVAL_7387 = _EVAL_4070 | _EVAL_4189;
  assign _EVAL_2638 = _EVAL_2258 & _EVAL_5117;
  assign _EVAL_17451 = _EVAL_11480 & 32'h2000034;
  assign _EVAL_9451 = _EVAL_18634 | _EVAL_528;
  assign _EVAL_19357 = _EVAL_11480[30:29];
  assign _EVAL_4673 = _EVAL_13158;
  assign _EVAL_15039 = _EVAL_17054 & _EVAL_4213;
  assign csr__EVAL_42 = _EVAL_10302;
  assign _EVAL_18800 = _EVAL_1397 & _EVAL_4961;
  assign _EVAL_14777 = div__EVAL_3 ? div__EVAL_4 : 32'h0;
  assign _EVAL_12232 = 3'h4 >> fetch__EVAL_8;
  assign _EVAL_1503 = _EVAL_11480[19:16];
  assign _EVAL_10858 = _EVAL_13977 & bpu__EVAL_33;
  assign fetch_pmp_checker__EVAL_3 = csr__EVAL_115;
  assign pmp_checker__EVAL_32 = csr__EVAL_49 ? csr__EVAL_30 : _EVAL_11443;
  assign _EVAL_19208 = _EVAL_13977 & bpu__EVAL_1;
  assign bpu__EVAL_41 = csr__EVAL_22;
  assign _EVAL_814 = _EVAL_2751 == _EVAL_15591;
  assign _EVAL_15003 = _EVAL_8452 & _EVAL_11823;
  assign _EVAL_10782 = _EVAL_9589 | _EVAL_13706;
  assign _EVAL_8706 = _EVAL_12568 & _EVAL_4213;
  assign _EVAL_98 = {1'b0,$signed(_EVAL_15785)};
  assign _EVAL_15431 = _EVAL_4467 | _EVAL_8958;
  assign _EVAL_869 = 32'h5013 == _EVAL_12413;
  assign _EVAL_16398 = fetch__EVAL & _EVAL_11251;
  assign _EVAL_2945 = _EVAL_7993 & _EVAL_8336;
  assign _EVAL_4834 = _EVAL_11480[30:20];
  assign csr__EVAL_17 = fetch__EVAL_8 ? {{16'd0}, _EVAL_11252} : fetch__EVAL_11;
  assign fetch_pmp_checker__EVAL_27 = csr__EVAL_92;
  assign _EVAL_9697 = _EVAL_18078;
  assign _EVAL_16751 = _EVAL_11480[19:12];
  assign _EVAL_1267 = _EVAL_16448 | _EVAL_5066;
  assign _EVAL_528 = 32'h2073 == _EVAL_1530;
  assign _EVAL_1404 = _EVAL_703 & _EVAL_14448;
  assign _EVAL_1067 = _EVAL_12850 | _EVAL_14001;
  assign bpu__EVAL_6 = csr__EVAL_48;
  assign _EVAL_7934 = 32'h2007033 == _EVAL_12413;
  assign _EVAL_3993 = $signed(_EVAL_18697) & -33'sh2000;
  assign _EVAL_12411 = _EVAL_10347 & 32'hfffffffe;
  assign _EVAL_1385 = $signed(_EVAL_14959) == 33'sh0;
  assign _EVAL_8178 = _EVAL_7387 & pmp_checker__EVAL_0;
  assign _EVAL_4184 = ~_EVAL_16398;
  assign _EVAL_27 = _EVAL_12503;
  assign _EVAL_10368 = _EVAL_15453 | _EVAL_16200;
  assign _EVAL_13022 = _EVAL_10148[15:0];
  assign _EVAL_15467 = _EVAL_16030 ? 1'h0 : _EVAL_16030;
  assign _EVAL_15801 = _EVAL_7895 | _EVAL_13225;
  assign _EVAL_15184 = ~_EVAL_18289;
  assign _EVAL_11858 = _EVAL_11480[13];
  assign _EVAL_13756 = _EVAL_5726 ? 3'h3 : 3'h2;
  assign _EVAL_12623 = _EVAL_3707 & csr__EVAL_123;
  assign _EVAL_3585 = _EVAL_9183 & _EVAL_4184;
  assign fetch__EVAL_5 = _EVAL_15497;
  assign _EVAL_3611 = _EVAL_12794 & _EVAL_11838;
  assign _EVAL_3170 = _EVAL_9061 | _EVAL_9429;
  assign _EVAL_17519 = _EVAL_8899 ? _EVAL_13756 : _EVAL_8051;
  assign _EVAL_6884 = _EVAL_16380 & _EVAL_11858;
  assign csr__EVAL_76 = _EVAL_11480[31:20];
  assign _EVAL_8610 = _EVAL_2706 == 32'h2010;
  assign csr__EVAL_40 = _EVAL_40;
  assign _EVAL_17358 = 32'h23 == _EVAL_1530;
  assign _EVAL_3352 = _EVAL_13093 | _EVAL_464;
  assign _EVAL_9822 = {_EVAL_2373,_EVAL_5960,_EVAL_5009,_EVAL_4673,_EVAL_13735,_EVAL_19285,1'h0};
  assign _EVAL_15561 = csr__EVAL_116 == 2'h3;
  assign _EVAL_16067 = 32'h5003 == _EVAL_1530;
  assign _EVAL_18439 = _EVAL_12302 | _EVAL_3875;
  assign _EVAL_12529 = 32'h3 == _EVAL_1530;
  assign _EVAL_1324 = _EVAL_10831 & _EVAL_15479;
  assign _EVAL_8070 = 32'h100f == _EVAL_1530;
  assign _EVAL_8128 = _EVAL_15427 ? _EVAL_880 : _EVAL_1027;
  assign _EVAL_8462 = _EVAL_17640 | _EVAL_17705;
  assign _EVAL_2706 = _EVAL_11480 & 32'h6034;
  assign _EVAL_12058 = _EVAL_16644;
  assign _EVAL_2793 = _EVAL_11480 & 32'h44;
  assign _EVAL_11609 = ~_EVAL_3495;
  assign _EVAL_4216 = _EVAL_18800 & _EVAL_15479;
  assign _EVAL_12083 = _EVAL_11480 & 32'hf800707f;
  assign _EVAL_849 = _EVAL_935 & _EVAL_13130;
  assign _EVAL_5960 = _EVAL_15418;
  assign fetch_pmp_checker__EVAL_29 = csr__EVAL_54;
  assign _EVAL_12603 = _EVAL_12751 | _EVAL_4361;
  assign _EVAL_9277 = _EVAL_11480[7];
  assign _EVAL_12251 = _EVAL_14478 ? _EVAL_14184 : _EVAL_6629;
  assign _EVAL_19273 = _EVAL_1;
  assign _EVAL_7194 = _EVAL_15591 != 5'h0;
  assign _EVAL_19144 = _EVAL_3495 & csr__EVAL_49;
  assign _EVAL_3888 = _EVAL_11480 & 32'h3050;
  assign _EVAL_12339 = {1'b0,$signed(_EVAL_6945)};
  assign _EVAL_10627 = _EVAL_9843 ^ 32'h20000000;
  assign _EVAL_14808 = _EVAL_15765 == 32'h0;
  assign _EVAL_8452 = _EVAL_14231 | _EVAL_17827;
  assign _EVAL_19597 = fetch__EVAL | _EVAL_14322;
  assign _EVAL_3841 = 32'h4063 == _EVAL_1530;
  assign _EVAL_8702 = 32'h2033 == _EVAL_12413;
  assign _EVAL_13977 = _EVAL_11531 | _EVAL_13099;
  assign _EVAL_17605 = _EVAL_11327 | _EVAL_15596;
  assign _EVAL_5613 = _EVAL_11868;
  assign pmp_checker__EVAL = _EVAL_36;
  assign _EVAL_15053 = _EVAL_12251;
  assign _EVAL_13389 = $signed(_EVAL_15238) & -33'sh4000;
  assign _EVAL_4027 = _EVAL_10156 | _EVAL_11154;
  assign _EVAL_18125 = _EVAL_19059;
  assign _EVAL_4521 = _EVAL_2258 & _EVAL_814;
  assign _EVAL_92 = {_EVAL_6454,_EVAL_15097};
  assign _EVAL_3902 = _EVAL_25;
  assign _EVAL_2109 = _EVAL_9689 | _EVAL_19509;
  assign _EVAL_9383 = _EVAL_2322 | _EVAL_284;
  assign _EVAL_50 = 1'h0;
  assign _EVAL_16351 = _EVAL_3585 & fetch__EVAL_1;
  assign _EVAL_1437 = _EVAL_12502 & _EVAL_5949;
  assign _EVAL_15723 = _EVAL_9556 ? {{1'd0}, _EVAL_12438} : _EVAL_10553;
  assign _EVAL_5162 = alu__EVAL_2[1];
  assign _EVAL_4688 = _EVAL_13144 | _EVAL_16739;
  assign _EVAL_17384 = _EVAL_17854 ? _EVAL_18125 : 32'h0;
  assign fetch__EVAL_23 = _EVAL_64;
  assign _EVAL_5612 = {_EVAL_17093,_EVAL_9075};
  assign div__EVAL_2 = _EVAL_12010 & _EVAL_1404;
  assign _EVAL_10331 = _EVAL_11480 & 32'h1c;
  assign _EVAL_11251 = _EVAL_7046 | _EVAL_5049;
  assign _EVAL_423 = _EVAL_15130[3:0];
  assign pmp_checker__EVAL_16 = csr__EVAL_7;
  assign _EVAL_12548 = _EVAL_7897 & _EVAL_12794;
  assign fetch_pmp_checker__EVAL_6 = csr__EVAL_44;
  assign pmp_checker__EVAL_9 = csr__EVAL_102;
  assign bpu__EVAL_22 = csr__EVAL_134;
  assign _EVAL_11327 = _EVAL_15349 | _EVAL_17358;
  assign csr__EVAL_55 = _EVAL_14196;
  assign _EVAL_2644 = _EVAL_10147 & _EVAL_1404;
  assign _EVAL_14183 = _EVAL_11480 & 32'h2004074;
  assign fetch_pmp_checker__EVAL_31 = csr__EVAL_66;
  assign _EVAL_15856 = _EVAL_19357 == 2'h0;
  assign _EVAL_15097 = _EVAL_11480[13:12];
  assign _EVAL_6530 = {_EVAL_2373,_EVAL_5960,_EVAL_5009,_EVAL_2373,_EVAL_13735,_EVAL_19285,_EVAL_9277};
  assign _EVAL_19337 = _EVAL_15755;
  assign _EVAL_10148 = _EVAL_53;
  assign _EVAL_7840 = _EVAL_5325 == 32'h2010;
  assign _EVAL_12794 = _EVAL_884;
  assign csr__EVAL_63 = _EVAL_64;
  assign _EVAL_897 = _EVAL_16898[0];
  assign _EVAL_11480 = fetch__EVAL_15;
  assign _EVAL_13007 = $signed(_EVAL_98) & -33'sh1000;
  assign _EVAL_4495 = _EVAL_11480[14:12];
  assign _EVAL_2125 = ~_EVAL_9119;
  assign pmp_checker__EVAL_15 = csr__EVAL_27;
  assign _EVAL_15829 = 1'h0;
  assign _EVAL_17383 = 32'h40000033 == _EVAL_12413;
  assign _EVAL_5117 = _EVAL_2751 == _EVAL_14920;
  assign _EVAL_9589 = _EVAL_15870 | _EVAL_15340;
  assign _EVAL_14892 = _EVAL_16668 & _EVAL_2492;
  assign _EVAL_948 = _EVAL_17986 | _EVAL_11894;
  assign fetch_pmp_checker__EVAL_19 = csr__EVAL_5;
  assign _EVAL_4872 = _EVAL_9378 & _EVAL_9583;
  assign _EVAL_24 = _EVAL_6830;
  assign _EVAL_5906 = 1'h0;
  assign _EVAL_3444 = fetch__EVAL & _EVAL_1969;
  assign pmp_checker__EVAL_13 = csr__EVAL_110;
  assign _EVAL_5949 = _EVAL_8865 | _EVAL_16380;
  assign fetch__EVAL_6 = _EVAL_9376 & _EVAL_9514;
  assign _EVAL_3248 = _EVAL_17213 | _EVAL_2021;
  assign _EVAL_2743 = _EVAL_7053 & _EVAL_18216;
  assign _EVAL_19544 = _EVAL_15785 ^ 32'h80000000;
  assign _EVAL_34 = csr__EVAL_103 & _EVAL_14107;
  assign _EVAL_17886 = csr__EVAL_4[0];
  assign _EVAL_7342 = _EVAL_13052;
  assign _EVAL_16389 = 1'h0;
  assign bpu__EVAL_31 = csr__EVAL_67;
  assign _EVAL_12018 = 32'h4033 == _EVAL_12413;
  assign _EVAL_2872 = _EVAL_16173 | _EVAL_5412;
  assign _EVAL_437 = 32'h2005033 == _EVAL_12413;
  assign _EVAL_6951 = _EVAL_35;
  assign _EVAL_7009 = 1'h0;
  assign _EVAL_1372 = _EVAL_16201 & _EVAL_9594;
  assign _EVAL_14765 = _EVAL_2743 ? _EVAL_16768 : _EVAL_17404;
  assign _EVAL_12502 = _EVAL_6064 & _EVAL_1739;
  assign _EVAL_21 = _EVAL_15053;
  assign _EVAL_10111 = csr__EVAL_49;
  assign _EVAL_10803 = $signed(_EVAL_4191) & -33'sh1000;
  assign _EVAL_10107 = _EVAL_48;
  assign _EVAL_588 = 32'h2006033 == _EVAL_12413;
  assign _EVAL_10371 = _EVAL_17584;
  assign _EVAL_7994 = _EVAL_16288 == 32'h0;
  assign _EVAL_14920 = fetch__EVAL_2;
  assign _EVAL_12395 = _EVAL_16796 & _EVAL_13097;
  assign _EVAL_1636 = ~_EVAL_16030;
  assign _EVAL_17625 = _EVAL_9241 == 32'h4;
  assign _EVAL_3495 = _EVAL_15312 & _EVAL_19458;
  assign fetch_pmp_checker__EVAL_25 = csr__EVAL_68;
  assign fetch__EVAL_18 = _EVAL_10896;
  assign _EVAL_14010 = 4'h1 << _EVAL_15097;
  assign fetch_pmp_checker__EVAL_10 = csr__EVAL_25;
  assign pmp_checker__EVAL_22 = csr__EVAL_74;
  assign fetch__EVAL_16 = _EVAL_12395 & _EVAL_11823;
  assign _EVAL_16872 = _EVAL_13311 ? _EVAL_14765 : 32'h0;
  assign _EVAL_13093 = _EVAL_8200 | _EVAL_982;
  assign _EVAL_8869 = {{14'd0}, _EVAL_434};
  assign _EVAL_8672 = ~_EVAL_6951;
  assign rf__EVAL_5 = ~_EVAL_15591;
  assign alu__EVAL_1 = _EVAL_1311 | _EVAL_2740;
  assign _EVAL_12302 = _EVAL_2238 | _EVAL_3841;
  assign _EVAL_14722 = _EVAL_11480 & 32'h1048;
  assign _EVAL_880 = {_EVAL_10764,_EVAL_10764,_EVAL_10764,_EVAL_10764};
  assign _EVAL_6064 = _EVAL_8990 & _EVAL_6146;
  assign _EVAL_3157 = _EVAL_67;
  assign _EVAL_11178 = _EVAL_16447 & _EVAL_10856;
  assign _EVAL_18697 = {1'b0,$signed(_EVAL_13761)};
  assign _EVAL_3102 = _EVAL_13723 ? _EVAL_7894 : 32'h0;
  assign _EVAL_11154 = 32'h2001033 == _EVAL_12413;
  assign _EVAL_1311 = _EVAL_14169 ? _EVAL_4157 : 32'h0;
  assign _EVAL_4090 = _EVAL_4680 | _EVAL_586;
  assign _EVAL_7378 = $signed(_EVAL_12444) & -33'sh2000;
  assign _EVAL_10302 = _EVAL_57;
  assign csr__EVAL_107 = _EVAL_2084 ? 32'h5 : _EVAL_10127;
  assign _EVAL_7502 = $signed(_EVAL_2727) == 33'sh0;
  assign _EVAL_3139 = _EVAL_1128 == 5'h0;
  assign _EVAL_9 = _EVAL_2265;
  assign _EVAL_2139 = _EVAL_12887 | _EVAL_3495;
  assign _EVAL_14682 = _EVAL_1962 | _EVAL_5252;
  assign _EVAL_11215 = csr__EVAL_101[10];
  assign _EVAL_15870 = _EVAL_1385 | _EVAL_1983;
  assign _EVAL_18671 = {{30'd0}, _EVAL_5933};
  assign fetch__EVAL_12 = _EVAL_36;
  assign _EVAL_9075 = _EVAL_17840 ? _EVAL_11356 : _EVAL_13022;
  assign _EVAL_9491 = fetch__EVAL & _EVAL_9364;
  assign _EVAL_9548 = {_EVAL_1811,_EVAL_15968};
  assign _EVAL_9556 = fetch__EVAL & _EVAL_13099;
  assign _EVAL_14763 = ~_EVAL_8584;
  assign _EVAL_12611 = _EVAL_14767;
  assign _EVAL_11129 = _EVAL_6190;
  assign _EVAL_16647 = _EVAL_3858 & _EVAL_9514;
  assign pmp_checker__EVAL_6 = csr__EVAL_44;
  assign _EVAL_1860 = _EVAL_8400 & _EVAL_15409;
  assign csr__EVAL_16 = _EVAL_36;
  assign _EVAL_4266 = _EVAL_10239 & _EVAL_9364;
  assign _EVAL_7483 = _EVAL_2941;
  assign _EVAL_4937 = _EVAL_12;
  assign _EVAL_12444 = {1'b0,$signed(_EVAL_17033)};
  assign csr__EVAL_109 = _EVAL_4475 ? alu__EVAL_2 : 32'h0;
  assign _EVAL_18210 = _EVAL_11480 & 32'h1014;
  assign _EVAL_6270 = _EVAL_11701 & _EVAL_5737;
  assign _EVAL_5146 = _EVAL_2953 | _EVAL_13198;
  assign _EVAL_8698 = ~_EVAL_14169;
  assign _EVAL_15617 = _EVAL_5138;
  assign _EVAL_14011 = _EVAL_5236 | _EVAL_18912;
  assign _EVAL_434 = {_EVAL_2644,1'h0,fetch__EVAL_19,_EVAL_2953,_EVAL_6248,_EVAL_11178,_EVAL_18030,1'h0,1'h0,_EVAL_15511};
  assign _EVAL_8110 = _EVAL_15768 | _EVAL_8999;
  assign _EVAL_5907 = _EVAL_17854 | _EVAL_13099;
  assign _EVAL_19610 = _EVAL_8228 == 32'h20;
  assign _EVAL_8627 = ~_EVAL_13609;
  assign _EVAL_18141 = _EVAL_11610 != 24'h0;
  assign _EVAL_11189 = _EVAL_11480 & 32'h2008;
  assign bpu__EVAL_20 = csr__EVAL_99;
  assign _EVAL_4295 = _EVAL_10858 | _EVAL_8148;
  assign _EVAL_17240 = csr__EVAL_59 ? 1'h0 : _EVAL_17371;
  assign _EVAL_6840 = _EVAL_14832 | _EVAL_8949;
  assign _EVAL_9768 = {_EVAL_11230,_EVAL_11230};
  assign _EVAL_59 = _EVAL_14650;
  assign _EVAL_42 = _EVAL_16649;
  assign _EVAL_7895 = _EVAL_17608 | _EVAL_2764;
  assign _EVAL_10491 = _EVAL_1372 ? 16'hffff : 16'h0;
  assign _EVAL_7800 = _EVAL_10012 | _EVAL_12216;
  assign _EVAL_9700 = _EVAL_4872 & _EVAL_19336;
  assign _EVAL_6571 = _EVAL_4647 & csr__EVAL_123;
  assign _EVAL_17963 = _EVAL_18439 | _EVAL_9565;
  assign _EVAL_15981 = _EVAL_1801 ? _EVAL_8999 : _EVAL_11162;
  assign _EVAL_16060 = {{29'd0}, _EVAL_12232};
  assign _EVAL_5684 = _EVAL_642 == 32'h20;
  assign _EVAL_17779 = _EVAL_9843 ^ 32'h80008000;
  assign _EVAL_13706 = $signed(_EVAL_8649) == 33'sh0;
  assign _EVAL_18565 = 32'h3073 == _EVAL_1530;
  assign _EVAL_9183 = _EVAL_12566 & fetch_pmp_checker__EVAL_0;
  assign _EVAL_4564 = ~_EVAL_6196;
  assign _EVAL_3623 = _EVAL_18905 | _EVAL_14879;
  assign _EVAL_11900 = $signed(_EVAL_5784) & -33'sh4000;
  assign _EVAL_15497 = _EVAL_32;
  assign _EVAL_2447 = _EVAL_18990;
  assign _EVAL_13130 = _EVAL_14920 != 5'h0;
  assign _EVAL_2086 = _EVAL_2845;
  assign fetch_pmp_checker__EVAL_22 = csr__EVAL_74;
  assign _EVAL_33 = _EVAL_16649;
  assign bpu__EVAL_15 = csr__EVAL_56;
  assign _EVAL_7156 = _EVAL_500;
  assign _EVAL_43 = _EVAL_16649;
  assign _EVAL_12751 = _EVAL_14808 | _EVAL_10622;
  assign _EVAL_15112 = fetch__EVAL & _EVAL_1739;
  assign _EVAL_2322 = _EVAL_948 | _EVAL_11521;
  assign _EVAL_1801 = _EVAL_11;
  assign _EVAL_12468 = _EVAL_16772 | _EVAL_16155;
  assign _EVAL_4961 = ~_EVAL_13099;
  assign _EVAL_14115 = {1'b0,$signed(_EVAL_10627)};
  assign _EVAL_884 = _EVAL_17887 | _EVAL_8412;
  assign _EVAL_241 = 1'h0;
  assign _EVAL_2488 = 32'h100073 == _EVAL_11480;
  assign _EVAL_15591 = fetch__EVAL_7;
  assign _EVAL_19509 = $signed(_EVAL_13002) == 33'sh0;
  assign _EVAL_11286 = _EVAL_12981 | _EVAL_9429;
  assign pmp_checker__EVAL_11 = csr__EVAL_41;
  assign _EVAL_16227 = _EVAL_12682 ? _EVAL_6053 : _EVAL_12525;
  assign _EVAL_16620 = _EVAL_11480 & 32'h1010;
  assign _EVAL_16377 = _EVAL_7614;
  assign _EVAL_13687 = _EVAL_11480 & 32'h3048;
  assign _EVAL_7414 = _EVAL_11480 & 32'h38;
  assign _EVAL_17716 = _EVAL_4297 == _EVAL_14920;
  assign _EVAL_13586 = 32'ha000202f == _EVAL_12083;
  assign bpu__EVAL_23 = csr__EVAL_20;
  assign _EVAL_13072 = 32'h0;
  assign _EVAL_127 = _EVAL_6400[2:0];
  assign _EVAL_221 = _EVAL_9119;
  assign _EVAL_7086 = _EVAL_5381 & _EVAL_13130;
  assign _EVAL_10928 = ~_EVAL_17801;
  assign _EVAL_2604 = _EVAL_15759 ? _EVAL_2215 : _EVAL_12268;
  assign _EVAL_4070 = _EVAL_7862 | _EVAL_6571;
  assign bpu__EVAL_38 = csr__EVAL_78;
  assign _EVAL_18410 = _EVAL_6449 | _EVAL_11005;
  assign _EVAL_17544 = {{13'd0}, _EVAL_18791};
  assign _EVAL_11807 = ~_EVAL_16866;
  assign _EVAL_3601 = _EVAL_11609 & _EVAL_1739;
  assign bpu__EVAL_29 = csr__EVAL_35;
  assign _EVAL_19529 = _EVAL_7993 | csr__EVAL_33;
  assign _EVAL_6533 = _EVAL_4157[31];
  assign _EVAL_17805 = _EVAL_2;
  assign pmp_checker__EVAL_20 = csr__EVAL_127;
  assign _EVAL_11443 = fetch__EVAL_21 & _EVAL_7689;
  assign _EVAL_6400 = _EVAL_16692;
  assign _EVAL_15461 = _EVAL_9667 | _EVAL_588;
  assign bpu__EVAL_12 = csr__EVAL_64;
  assign div__EVAL_1 = _EVAL_3495;
  assign _EVAL_11894 = 32'h30200073 == _EVAL_11480;
  assign _EVAL_17054 = _EVAL_9086 & _EVAL_1739;
  assign _EVAL_4157 = _EVAL_6270 ? _EVAL_16768 : _EVAL_7879;
  assign _EVAL_16854 = _EVAL_18210 == 32'h1010;
  assign _EVAL_14257 = _EVAL_11480 & 32'h40000034;
  assign _EVAL_10127 = _EVAL_17995 ? _EVAL_13045 : {{28'd0}, _EVAL_8759};
  assign _EVAL_7137 = _EVAL_3491 | _EVAL_14680;
  assign _EVAL_19336 = ~_EVAL_5146;
  assign _EVAL_7046 = _EVAL_15976 | _EVAL_18202;
  assign csr__EVAL_101 = _EVAL_11480[31:20];
  assign _EVAL_10679 = ~_EVAL_5301;
  assign _EVAL_2446 = _EVAL_4297 == _EVAL_15591;
  assign bpu__EVAL_21 = csr__EVAL_97;
  assign _EVAL_19340 = _EVAL_9429 | _EVAL_5512;
  assign _EVAL_12957 = _EVAL_10181;
  assign _EVAL_13097 = _EVAL_1638 | _EVAL_14231;
  assign _EVAL_8400 = _EVAL_4213 & _EVAL_13130;
  assign _EVAL_15690 = _EVAL_11480 & 32'h28;
  assign _EVAL_15947 = _EVAL_15785 ^ 32'h80008000;
  assign _EVAL_840 = _EVAL_15039 & _EVAL_13130;
  assign _EVAL_14879 = 32'h40005033 == _EVAL_12413;
  assign _EVAL_2021 = 32'h2004033 == _EVAL_12413;
  assign _EVAL_874 = _EVAL_15690 == 32'h0;
  assign _EVAL_17285 = _EVAL_1888[32:0];
  assign csr__EVAL_18 = _EVAL_1311 | _EVAL_9792;
  assign _EVAL_3104 = _EVAL_68;
  assign div__EVAL_6 = _EVAL_36;
  assign _EVAL_11311 = 32'h1063 == _EVAL_1530;
  assign _EVAL_6830 = 1'h1;
  assign _EVAL_5164 = 1'h0;
  assign _EVAL_12268 = csr__EVAL_49 ? 3'h4 : _EVAL_15723;
  assign _EVAL_9594 = _EVAL_9075[15];
  assign _EVAL_8299 = {_EVAL_7840,_EVAL_16854};
  assign _EVAL_3045 = _EVAL_11480 & 32'h78;
  assign _EVAL_18452 = _EVAL_11480 & 32'h4014;
  assign _EVAL_16949 = _EVAL_7;
  assign fetch__EVAL_21 = alu__EVAL_2;
  assign _EVAL_30 = _EVAL_15112 & _EVAL_5625;
  assign _EVAL_8865 = _EVAL_3888 == 32'h50;
  assign _EVAL_17356 = _EVAL_403 | _EVAL_12529;
  assign _EVAL_11578 = _EVAL_9451 | _EVAL_18565;
  assign fetch_pmp_checker__EVAL_32 = ~_EVAL_14156;
  assign _EVAL_2761 = _EVAL_16380 & _EVAL_6454;
  assign _EVAL_18 = _EVAL_16649;
  assign _EVAL_1888 = 33'h100000000 - 33'h1;
  assign _EVAL_18618 = 1'h0;
  assign _EVAL_17827 = _EVAL_16351 & _EVAL_10233;
  assign _EVAL_10091 = 32'h4013 == _EVAL_1530;
  assign _EVAL_18030 = ~fetch__EVAL;
  assign _EVAL_9792 = _EVAL_8698 ? _EVAL_236 : 32'h0;
  assign _EVAL_13052 = csr__EVAL_83;
  assign _EVAL_14418 = _EVAL_1988 == 32'h0;
  assign _EVAL_16173 = _EVAL_12477 & _EVAL_18877;
  assign pmp_checker__EVAL_8 = csr__EVAL_82;
  assign _EVAL_18613 = _EVAL_5162 ? 2'h0 : _EVAL_1745;
  assign _EVAL_4680 = _EVAL_12794 & _EVAL_17674;
  assign _EVAL_7614 = {_EVAL_2373,_EVAL_5960,_EVAL_12793,_EVAL_17688,_EVAL_13735,_EVAL_16395,1'h0};
  assign _EVAL_5622 = _EVAL_4709[31:0];
  assign _EVAL_11278 = 32'h1003 == _EVAL_1530;
  assign _EVAL_13723 = _EVAL_413 | _EVAL_4361;
  assign _EVAL_3556 = 32'h3033 == _EVAL_12413;
  assign _EVAL_13157 = _EVAL_7800 | _EVAL_6767;
  assign _EVAL_10444 = _EVAL_952 | _EVAL_2293;
  assign _EVAL_706 = _EVAL_17625 | _EVAL_16094;
  assign _EVAL_9364 = _EVAL_13977 | _EVAL_17854;
  assign _EVAL_17674 = ~_EVAL_7897;
  assign _EVAL_6735 = _EVAL_15759 ? _EVAL_4377 : _EVAL_5590;
  assign _EVAL_427 = _EVAL_3837;
  assign _EVAL_13311 = _EVAL_8228 == 32'h30;
  assign _EVAL_2941 = $signed(_EVAL_3544) & -33'sh4000;
  assign _EVAL_4663 = _EVAL_15785 ^ 32'h4000;
  assign _EVAL_15396 = _EVAL_2604;
  assign _EVAL_3497 = _EVAL_15112 & _EVAL_8627;
  assign _EVAL_14156 = _EVAL_5341 | 32'h3;
  assign _EVAL_14809 = _EVAL_3330 == 32'h1050;
  assign _EVAL_10383 = fetch__EVAL_3;
  assign _EVAL_17995 = _EVAL_11321 | _EVAL_11251;
  assign csr__EVAL_87 = _EVAL_17371;
  assign _EVAL_14051 = _EVAL_17717 == 2'h1;
  assign _EVAL_5252 = _EVAL_9364 & _EVAL_15759;
  assign _EVAL_18905 = _EVAL_12468 | _EVAL_8195;
  assign _EVAL_5728 = _EVAL_19578 ? 1'h0 : 1'h1;
  assign _EVAL_8534 = _EVAL_12439 | _EVAL_17194;
  assign bpu__EVAL_14 = alu__EVAL_2;
  assign _EVAL_3816 = _EVAL_7407 & _EVAL_9378;
  assign csr__EVAL_59 = _EVAL_17283 | _EVAL_17371;
  assign _EVAL_4213 = _EVAL_12608 | _EVAL_19368;
  assign fetch_pmp_checker__EVAL_8 = csr__EVAL_82;
  assign _EVAL_3741 = _EVAL_10383 == 5'h0;
  assign _EVAL_5227 = _EVAL_7638 & _EVAL_18141;
  assign _EVAL_18247 = _EVAL_14053 | _EVAL_11162;
  assign _EVAL_7879 = _EVAL_3741 ? 32'h0 : rf__EVAL_0;
  assign _EVAL_500 = _EVAL_14478 ? _EVAL_10593 : _EVAL_15561;
  assign _EVAL_10668 = csr__EVAL_49 ? _EVAL_17285 : {{29'd0}, _EVAL_12829};
  assign csr__EVAL_39 = _EVAL_15382 | _EVAL_2084;
  assign _EVAL_5579 = _EVAL_15545;
  assign _EVAL_5171 = {8{_EVAL_12957}};
  assign _EVAL_15511 = _EVAL_9882 | _EVAL_8163;
  assign _EVAL_7201 = _EVAL_19578 | _EVAL_12476;
  assign fetch_pmp_checker__EVAL_12 = csr__EVAL_133;
  assign _EVAL_6765 = _EVAL_11480 & 32'h24;
  assign _EVAL_551 = _EVAL_14322 ? 2'h1 : _EVAL_2900;
  assign _EVAL_4453 = _EVAL_15759 ? _EVAL_2097 : {{2'd0}, _EVAL_16547};
  assign _EVAL_4475 = _EVAL_3601 & _EVAL_8112;
  assign _EVAL_19212 = _EVAL_60;
  assign _EVAL_968 = 1'h0;
  assign _EVAL_1185 = {1'b0,$signed(_EVAL_15947)};
  assign _EVAL_17821 = _EVAL_15272 | _EVAL_2084;
  assign _EVAL_6248 = _EVAL_13253 & _EVAL_16024;
  assign _EVAL_66 = _EVAL_16649;
  assign _EVAL_8601 = _EVAL_636 ? _EVAL_5622 : 32'h0;
  assign _EVAL_52 = _EVAL_7156;
  assign _EVAL_17608 = _EVAL_2654 | _EVAL_2835;
  assign _EVAL_19 = _EVAL_12244;
  assign _EVAL_12732 = _EVAL_14892 | _EVAL_8864;
  assign _EVAL_8137 = _EVAL_4257 & _EVAL_7194;
  assign _EVAL_9411 = _EVAL_6941 & _EVAL_4660;
  assign _EVAL_7868 = _EVAL_15785 ^ 32'h2000000;
  assign fetch_pmp_checker__EVAL_15 = csr__EVAL_27;
  assign _EVAL_6156 = _EVAL_3852 | _EVAL_8610;
  assign _EVAL_14322 = fetch__EVAL ? fetch__EVAL_4 : _EVAL_17967;
  assign _EVAL_13874 = _EVAL_17451 == 32'h2000030;
  assign _EVAL_4218 = _EVAL_6481 | _EVAL_6571;
  assign _EVAL_2764 = _EVAL_5907 & _EVAL_11807;
  assign _EVAL_12356 = ~_EVAL_9183;
  assign _EVAL_15479 = ~csr__EVAL_49;
  assign _EVAL_15238 = {1'b0,$signed(_EVAL_16867)};
  assign _EVAL_14855 = 1'h1;
  assign _EVAL_13703 = fetch__EVAL & _EVAL_5146;
  assign _EVAL_37 = _EVAL_6830;
  assign _EVAL_4753 = _EVAL_10140 | _EVAL_9449;
  assign _EVAL_10856 = _EVAL_15768 ? _EVAL_8999 : _EVAL_11162;
  assign _EVAL_8923 = _EVAL_7994 | _EVAL_10622;
  assign pmp_checker__EVAL_33 = csr__EVAL_14;
  assign _EVAL_16547 = csr__EVAL_49 ? 2'h2 : _EVAL_15097;
  assign _EVAL_403 = _EVAL_15411 | _EVAL_1738;
  assign _EVAL_17583 = _EVAL_874 | _EVAL_11458;
  assign _EVAL_12793 = _EVAL_19607;
  assign _EVAL_5236 = $signed(_EVAL_7483) == 33'sh0;
  assign _EVAL_12968 = _EVAL_18452 == 32'h4010;
  assign _EVAL_6756 = _EVAL_12411 + _EVAL_9169;
  assign _EVAL_15656 = _EVAL_2084 | _EVAL_17240;
  assign _EVAL_6481 = _EVAL_7862 | _EVAL_7502;
  assign rf__EVAL_3 = ~_EVAL_10383;
  assign _EVAL_1397 = _EVAL_840 & _EVAL_319;
  assign _EVAL_6999 = _EVAL_16668 | _EVAL_2258;
  assign _EVAL_17118 = _EVAL_17717 == 2'h0;
  assign _EVAL_65 = _EVAL_6830;
  assign _EVAL_45 = _EVAL_641;
  assign _EVAL_6286 = 32'h2003033 == _EVAL_12413;
  assign _EVAL_11321 = _EVAL_6741 | _EVAL_14322;
  assign _EVAL_2458 = 32'he000202f == _EVAL_12083;
  assign _EVAL_17997 = _EVAL_4453;
  assign _EVAL_14159 = _EVAL_2793 == 32'h40;
  assign _EVAL_16306 = _EVAL_3497 & _EVAL_5146;
  assign bpu__EVAL_7 = csr__EVAL_122;
  assign bpu__EVAL_2 = _EVAL_10347 & 32'hfffffffe;
  assign _EVAL_38 = _EVAL_16649;
  assign _EVAL_16804 = _EVAL_64;
  assign _EVAL_2084 = csr__EVAL_49 & _EVAL_18773;
  assign _EVAL_9565 = 32'h5063 == _EVAL_1530;
  assign _EVAL_13694 = {1'b0,$signed(_EVAL_7868)};
  assign _EVAL_14053 = ~_EVAL_15768;
  assign alu__EVAL = {_EVAL_3973,_EVAL_8299};
  assign _EVAL_6789 = ~_EVAL_6941;
  assign _EVAL_8292 = _EVAL_2113 | _EVAL_8601;
  assign _EVAL_3448 = 32'h7013 == _EVAL_1530;
  assign _EVAL_6492 = _EVAL_11480[15];
  assign _EVAL_16772 = _EVAL_1267 | _EVAL_12018;
  assign fetch__EVAL_0 = _EVAL_19212;
  assign _EVAL_2558 = _EVAL_1297 | _EVAL_3556;
  assign _EVAL_6454 = ~_EVAL_5648;
  assign _EVAL_6584 = _EVAL_16380 | _EVAL_8865;
  assign rf__EVAL_6 = _EVAL_36;
  assign _EVAL_639 = _EVAL_1324 & _EVAL_19458;
  assign _EVAL_13609 = _EVAL_4381 | _EVAL_3442;
  assign _EVAL_19368 = _EVAL_19611 == 32'h2010;
  assign _EVAL_9734 = _EVAL_13371 & _EVAL_5387;
  assign _EVAL_12009 = _EVAL_18452 == 32'h10;
  assign _EVAL_13304 = _EVAL_14920 == _EVAL_14896;
  assign _EVAL_4030 = _EVAL_17625 ? _EVAL_12360 : 32'h0;
  assign _EVAL_18401 = _EVAL_4295 ? 3'h3 : _EVAL_3302;
  assign _EVAL_8200 = _EVAL_11578 | _EVAL_637;
  assign _EVAL_2508 = _EVAL_10948 | _EVAL_1627;
  assign _EVAL_16034 = 32'h2003 == _EVAL_1530;
  assign _EVAL_641 = _EVAL_1606;
  assign _EVAL_9496 = ~_EVAL_3352;
  assign _EVAL_1451 = {_EVAL_6584,_EVAL_13099,_EVAL_17854,_EVAL_11531,1'h0};
  assign _EVAL_1336 = _EVAL_31;
  assign _EVAL_11823 = _EVAL_13906 & _EVAL_8917;
  assign _EVAL_12096 = 32'h4003 == _EVAL_1530;
  assign _EVAL_7717 = _EVAL_8292 | _EVAL_9039;
  assign _EVAL_10480 = _EVAL_7717 | _EVAL_14777;
  assign fetch_pmp_checker__EVAL_23 = csr__EVAL_116;
  assign _EVAL_18791 = {_EVAL_6719,_EVAL_18289,_EVAL_4361,_EVAL_8872,_EVAL_6422,_EVAL_19031,_EVAL_1451};
  assign pmp_checker__EVAL_31 = csr__EVAL_66;
  assign _EVAL_28 = csr__EVAL_8 & _EVAL_14107;
  assign _EVAL_3973 = {_EVAL_13874,_EVAL_8462,_EVAL_12968};
  assign _EVAL_8336 = ~_EVAL_15511;
  assign _EVAL_6629 = _EVAL_17560 & 32'hfffffffc;
  assign _EVAL_6422 = _EVAL_4973 == 32'h40;
  assign _EVAL_17404 = _EVAL_8892 ? 32'h0 : rf__EVAL_2;
  assign _EVAL_6548 = _EVAL_477 | _EVAL_4189;
  assign _EVAL_14092 = _EVAL_16668 & _EVAL_17716;
  assign _EVAL_637 = 32'h5073 == _EVAL_1530;
  assign _EVAL_17570 = _EVAL_9941 & _EVAL_1995;
  assign fetch_pmp_checker__EVAL_5 = csr__EVAL_77;
  assign _EVAL_16407 = ~_EVAL_11215;
  assign _EVAL_16155 = 32'h1033 == _EVAL_12413;
  assign _EVAL_1087 = _EVAL_23;
  assign _EVAL_2080 = _EVAL_5907 & bpu__EVAL_30;
  assign _EVAL_3630 = _EVAL_5612[31:8];
  assign _EVAL_9882 = _EVAL_6252 & _EVAL_12732;
  assign _EVAL_10140 = _EVAL_11286 | csr__EVAL_49;
  assign _EVAL_14169 = _EVAL_12603 | _EVAL_12009;
  assign bpu__EVAL_19 = csr__EVAL_139;
  assign _EVAL_3837 = $signed(_EVAL_4042) & -33'sh2000;
  assign csr__EVAL_51 = _EVAL_2084 ? csr__EVAL_30 : _EVAL_12411;
  assign bpu__EVAL_16 = csr__EVAL_19;
  assign bpu__EVAL_26 = csr__EVAL_135;
  assign _EVAL_15890 = _EVAL_11480[27];
  assign _EVAL_8607 = _EVAL_15461 | _EVAL_7934;
  assign _EVAL_2703 = _EVAL_9822;
  assign _EVAL_3875 = 32'h6063 == _EVAL_1530;
  assign _EVAL_8899 = _EVAL_11480[30];
  assign _EVAL_19031 = _EVAL_4213 & _EVAL_10919;
  assign _EVAL_2871 = csr__EVAL_124;
  assign _EVAL_15130 = _EVAL_14010 - 4'h1;
  assign _EVAL_17934 = _EVAL_4266 & _EVAL_19458;
  assign _EVAL_11610 = _EVAL_16898 & _EVAL_17544;
  assign _EVAL_12929 = _EVAL_5332 ? 4'he : {{1'd0}, _EVAL_18401};
  assign bpu__EVAL = csr__EVAL_10;
  assign _EVAL_8949 = 32'h3013 == _EVAL_1530;
  assign _EVAL_1811 = _EVAL_17118 ? _EVAL_2100 : _EVAL_3630;
  assign _EVAL_3117 = _EVAL_13977 & _EVAL_15479;
  assign _EVAL_13144 = csr__EVAL_49 & csr__EVAL_39;
  assign _EVAL_919 = 1'h1;
  assign _EVAL_7880 = _EVAL_15759 ? {{29'd0}, _EVAL_6792} : _EVAL_10668;
  assign csr__EVAL_121 = _EVAL_13;
  assign _EVAL_13129 = _EVAL_18360 | _EVAL_2945;
  assign _EVAL_6586 = _EVAL_11480 & 32'h30;
  assign _EVAL_2654 = _EVAL_9364 & _EVAL_8584;
  assign _EVAL_16447 = _EVAL_9364 | csr__EVAL_49;
  assign _EVAL_19013 = fetch__EVAL & _EVAL_16380;
  assign _EVAL_13906 = _EVAL_15479 & _EVAL_19458;
  assign _EVAL_7679 = $signed(_EVAL_1185) & -33'sh4000;
  assign _EVAL_19090 = _EVAL_6735;
  assign _EVAL_1638 = _EVAL_3585 & _EVAL_10233;
  assign _EVAL_12503 = 3'h4;
  assign _EVAL_13225 = _EVAL_13977 & _EVAL_18773;
  assign _EVAL_7142 = $signed(_EVAL_5613) == 33'sh0;
  assign _EVAL_4626 = 1'h1;
  assign _EVAL_13099 = _EVAL_15504 == 32'h2008;
  assign _EVAL_12424 = csr__EVAL_95;
  assign _EVAL_10764 = _EVAL_14765[7:0];
  assign _EVAL_7611 = _EVAL_909 | _EVAL_3320;
  assign _EVAL_16739 = csr__EVAL_59 ? 1'h0 : _EVAL_9449;
  assign _EVAL_2198 = _EVAL_13157 | _EVAL_10566;
  assign _EVAL_586 = _EVAL_12548 ? 1'h0 : _EVAL_15759;
  assign _EVAL_9241 = _EVAL_11480 & 32'h4c;
  assign _EVAL_16164 = _EVAL_11596 & _EVAL_8336;
  assign _EVAL_16869 = _EVAL_11480 & 32'h2000050;
  assign bpu__EVAL_0 = csr__EVAL_65;
  assign pmp_checker__EVAL_30 = csr__EVAL_89;
  assign _EVAL_15 = _EVAL_6830;
  assign _EVAL_2277 = ~fetch__EVAL_9;
  assign _EVAL_3544 = {1'b0,$signed(_EVAL_19544)};
  assign _EVAL_8649 = _EVAL_10803;
  assign _EVAL_12589 = _EVAL_15431 | _EVAL_7993;
  assign _EVAL_4973 = _EVAL_11480 & 32'h54;
  assign _EVAL_13002 = _EVAL_6214;
  assign _EVAL_7894 = _EVAL_15617;
  assign bpu__EVAL_35 = csr__EVAL_94;
  assign pmp_checker__EVAL_2 = csr__EVAL_62;
  assign _EVAL_3607 = _EVAL_13835;
  assign _EVAL_5784 = {1'b0,$signed(_EVAL_17779)};
  assign _EVAL_9376 = _EVAL_16306 & _EVAL_8178;
  assign fetch_pmp_checker__EVAL_1 = csr__EVAL_73;
  assign pmp_checker__EVAL_17 = csr__EVAL_86;
  assign _EVAL_15765 = _EVAL_11480 & 32'h50;
  assign _EVAL_4267 = _EVAL_16898 & _EVAL_8869;
  assign _EVAL_11046 = _EVAL_16380 & csr__EVAL_111;
  assign _EVAL_17840 = _EVAL_13287[1];
  assign _EVAL_14767 = {_EVAL_8873,_EVAL_4157};
  assign _EVAL_5590 = csr__EVAL_49 ? 3'h0 : _EVAL_5001;
  assign _EVAL_5566 = ~_EVAL_4753;
  assign _EVAL_5737 = _EVAL_14896 == _EVAL_10383;
  assign _EVAL_17213 = _EVAL_18642 | _EVAL_409;
  assign _EVAL_12566 = _EVAL_5883 | _EVAL_7142;
  assign _EVAL_15553 = _EVAL_10289 | _EVAL_9658;
  assign div__EVAL_8 = {{1'd0}, _EVAL_4495};
  assign _EVAL_18942 = _EVAL_9734 | _EVAL_16543;
  assign _EVAL_2835 = _EVAL_13099 & _EVAL_4564;
  assign fetch_pmp_checker__EVAL_2 = csr__EVAL_62;
  assign _EVAL_1738 = 32'h17 == _EVAL_6918;
  assign _EVAL_477 = _EVAL_17254 | _EVAL_6571;
  assign _EVAL_12521 = _EVAL_4157 == _EVAL_14765;
  assign _EVAL_6146 = ~_EVAL_7086;
  assign _EVAL_12173 = bpu__EVAL_42 ? 2'h3 : _EVAL_551;
  assign _EVAL_14959 = _EVAL_13389;
  assign _EVAL_5325 = _EVAL_11480 & 32'h2014;
  assign bpu__EVAL_13 = csr__EVAL_79;
  assign _EVAL_1739 = ~_EVAL_17995;
  assign _EVAL_3858 = _EVAL_5962;
  assign _EVAL_13825 = bpu__EVAL_34 ? 4'he : {{2'd0}, _EVAL_12173};
  assign _EVAL_15349 = _EVAL_7487 | _EVAL_16067;
  assign pmp_checker__EVAL_14 = csr__EVAL_46;
  assign _EVAL_2629 = _EVAL_17074 & _EVAL_15856;
  assign _EVAL_15768 = _EVAL_11218;
  assign _EVAL_464 = 32'h7073 == _EVAL_1530;
  assign _EVAL_236 = _EVAL_2086;
  assign _EVAL_4647 = $signed(_EVAL_4798) == 33'sh0;
  assign _EVAL_10975 = _EVAL_11858 | _EVAL_7366;
  assign pmp_checker__EVAL_27 = csr__EVAL_92;
  assign _EVAL_9820 = _EVAL_9843 ^ 32'h40000000;
  assign _EVAL_5625 = ~_EVAL_1962;
  assign _EVAL_6741 = _EVAL_13210 | bpu__EVAL_42;
  assign _EVAL_63 = _EVAL_12794;
  assign _EVAL_11875 = _EVAL_12427 | _EVAL_3593;
  assign pmp_checker__EVAL_25 = csr__EVAL_68;
  assign _EVAL_4888 = _EVAL_11480[20];
  assign _EVAL_0 = _EVAL_16649;
  assign _EVAL_19607 = _EVAL_16751;
  assign _EVAL_18877 = _EVAL_13298 | _EVAL_9965;
  assign pmp_checker__EVAL_1 = csr__EVAL_73;
  assign _EVAL_3491 = _EVAL_3858 & _EVAL_8672;
  assign _EVAL_5 = _EVAL_6830;
  assign _EVAL_18449 = _EVAL_10444 | _EVAL_10091;
  assign _EVAL_8759 = _EVAL_8112 ? _EVAL_12929 : 4'h0;
  assign _EVAL_3322 = _EVAL_2703;
  assign csr__EVAL_43 = _EVAL_16;
  assign _EVAL_14001 = 32'h73 == _EVAL_11480;
  assign _EVAL_982 = 32'h6073 == _EVAL_1530;
  assign _EVAL_14650 = 4'h2;
  assign _EVAL_16256 = _EVAL_10588 == 32'h2050;
  assign _EVAL_12352 = _EVAL_8872 ? _EVAL_14251 : 32'h0;
  assign _EVAL_10051 = _EVAL_9378 | _EVAL_19340;
  assign _EVAL_14356 = _EVAL_6789 & _EVAL_2277;
  assign _EVAL_16094 = _EVAL_16869 == 32'h10;
  assign _EVAL_12413 = _EVAL_11480 & 32'hfe00707f;
  assign _EVAL_17717 = _EVAL_1801 ? _EVAL_7693 : _EVAL_2667;
  assign _EVAL_4045 = _EVAL_6422 ? _EVAL_3322 : 32'h0;
  assign _EVAL_12608 = _EVAL_7611 | _EVAL_17740;
  assign _EVAL_18258 = _EVAL_14682 | _EVAL_849;
  assign _EVAL_8872 = _EVAL_15131 == 32'h48;
  assign bpu__EVAL_40 = csr__EVAL_117;
  assign _EVAL_6941 = _EVAL_11162 | _EVAL_8999;
  assign _EVAL_2832 = alu__EVAL_2 & _EVAL_18671;
  assign _EVAL_11596 = _EVAL_13703 & _EVAL_1739;
  assign _EVAL_16866 = _EVAL_2109 & pmp_checker__EVAL_24;
  assign _EVAL_12439 = _EVAL_11162 & _EVAL_8342;
  assign _EVAL_18634 = _EVAL_9383 | _EVAL_8013;
  assign _EVAL_8917 = ~_EVAL_2871;
  assign _EVAL_12191 = _EVAL_8923 | _EVAL_14418;
  assign _EVAL_15755 = {_EVAL_10975,_EVAL_14765};
  assign _EVAL_10778 = _EVAL_12191 | _EVAL_9545;
  assign fetch_pmp_checker__EVAL_17 = csr__EVAL_86;
  assign _EVAL_17705 = _EVAL_805 == 32'h40001010;
  assign _EVAL_18773 = ~_EVAL_14142;
  assign fetch_pmp_checker__EVAL_16 = csr__EVAL_7;
  assign _EVAL_2113 = _EVAL_19013 ? csr__EVAL_34 : 32'h0;
  assign _EVAL_15312 = csr__EVAL_50 & _EVAL_10679;
  assign _EVAL_7407 = _EVAL_10831 & _EVAL_1739;
  assign _EVAL_9658 = 32'h1013 == _EVAL_12413;
  assign _EVAL_3707 = $signed(_EVAL_10019) == 33'sh0;
  assign _EVAL_2100 = _EVAL_15974 ? 24'hffffff : 24'h0;
  assign rf__EVAL = _EVAL_17570 ? _EVAL_9548 : _EVAL_16768;
  assign _EVAL_15411 = _EVAL_18410 | _EVAL_4545;
  assign _EVAL_4467 = _EVAL_17543 | _EVAL_5146;
  assign _EVAL_7689 = ~_EVAL_4450;
  assign _EVAL_10156 = 32'h2000033 == _EVAL_12413;
  assign _EVAL_15453 = _EVAL_17605 | _EVAL_4619;
  assign _EVAL_4189 = $signed(_EVAL_8187) == 33'sh0;
  assign _EVAL_15785 = csr__EVAL_49 ? csr__EVAL_30 : _EVAL_11443;
  assign _EVAL_5933 = _EVAL_423[1:0];
  assign bpu__EVAL_18 = csr__EVAL_71;
  assign _EVAL_62 = _EVAL_13133;
  assign fetch_pmp_checker__EVAL_9 = csr__EVAL_102;
  assign _EVAL_11607 = _EVAL_11480 & 32'h2000074;
  assign _EVAL_16867 = _EVAL_9843 ^ 32'h80000000;
  assign _EVAL_17211 = _EVAL_9449 & csr__EVAL_59;
  assign _EVAL_7862 = _EVAL_5589 | _EVAL_17352;
  assign _EVAL_16692 = _EVAL_15759 ? _EVAL_10894 : _EVAL_15785;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_2097 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_2215 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_2667 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_2751 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_3051 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_3130 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_4297 = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_4377 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_5301 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_5564 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_5900 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_6190 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_6538 = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_6647 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_6792 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_7693 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_8342 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_8580 = _RAND_17[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_8631 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_8874 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_8999 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_9119 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_9429 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_9449 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_9510 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_10347 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_10353 = _RAND_26[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_10468 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_10593 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_10894 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_11162 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_12371 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _EVAL_12379 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _EVAL_12498 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _EVAL_12508 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _EVAL_12724 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _EVAL_13327 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _EVAL_14160 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _EVAL_14184 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _EVAL_14478 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _EVAL_14896 = _RAND_40[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _EVAL_15545 = _RAND_41[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _EVAL_15759 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _EVAL_16030 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _EVAL_16096 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _EVAL_16207 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _EVAL_16543 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _EVAL_16644 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _EVAL_16733 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _EVAL_16768 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _EVAL_17371 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _EVAL_17801 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _EVAL_18514 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _EVAL_19551 = _RAND_53[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_36) begin
    if (_EVAL_3611) begin
      _EVAL_2097 <= _EVAL_17997;
    end
    if (_EVAL_3611) begin
      _EVAL_2215 <= _EVAL_15396;
    end
    if (_EVAL_8339) begin
      if (~_EVAL_15768) begin
        _EVAL_2667 <= _EVAL_15097;
      end
    end
    if (_EVAL_8339) begin
      if (_EVAL_15768) begin
        _EVAL_2751 <= _EVAL_14920;
      end
    end
    if (_EVAL_3611) begin
      _EVAL_3051 <= _EVAL_641;
    end
    _EVAL_3130 <= _EVAL_17570 & _EVAL_16096;
    if (_EVAL_8339) begin
      if (~_EVAL_15768) begin
        _EVAL_4297 <= _EVAL_14920;
      end
    end
    if (_EVAL_3611) begin
      _EVAL_4377 <= _EVAL_19090;
    end
    if (_EVAL_64) begin
      _EVAL_5301 <= 1'h0;
    end else if (_EVAL_13144) begin
      _EVAL_5301 <= 1'h0;
    end else begin
      _EVAL_5301 <= _EVAL_3820;
    end
    if (_EVAL_64) begin
      _EVAL_5564 <= 1'h0;
    end else begin
      _EVAL_5564 <= _EVAL_2872;
    end
    if (_EVAL_8339) begin
      if (~_EVAL_15768) begin
        _EVAL_5900 <= _EVAL_127;
      end
    end
    _EVAL_6190 <= csr__EVAL_91;
    _EVAL_6538 <= fetch__EVAL_7;
    if (_EVAL_8339) begin
      if (_EVAL_15768) begin
        _EVAL_6647 <= _EVAL_3117;
      end
    end
    if (_EVAL_3611) begin
      _EVAL_6792 <= _EVAL_13133;
    end
    if (_EVAL_8339) begin
      if (_EVAL_15768) begin
        _EVAL_7693 <= _EVAL_15097;
      end
    end
    if (_EVAL_8339) begin
      if (~_EVAL_15768) begin
        _EVAL_8342 <= _EVAL_17140;
      end
    end
    _EVAL_8580 <= fetch__EVAL_3;
    if (_EVAL_2743) begin
      _EVAL_8631 <= _EVAL_16768;
    end else if (_EVAL_8892) begin
      _EVAL_8631 <= 32'h0;
    end else begin
      _EVAL_8631 <= rf__EVAL_2;
    end
    if (_EVAL_8339) begin
      if (_EVAL_15768) begin
        _EVAL_8874 <= _EVAL_10111;
      end
    end
    if (_EVAL_64) begin
      _EVAL_8999 <= 1'h0;
    end else if (_EVAL_13371) begin
      if (_EVAL_1801) begin
        _EVAL_8999 <= 1'h0;
      end else if (_EVAL_8339) begin
        _EVAL_8999 <= _EVAL_8110;
      end
    end else if (_EVAL_8339) begin
      _EVAL_8999 <= _EVAL_8110;
    end
    _EVAL_9119 <= csr__EVAL_75;
    if (_EVAL_64) begin
      _EVAL_9429 <= 1'h0;
    end else if (_EVAL_9378) begin
      _EVAL_9429 <= _EVAL_3170;
    end else if (_EVAL_9429) begin
      _EVAL_9429 <= 1'h0;
    end else begin
      _EVAL_9429 <= _EVAL_3170;
    end
    if (_EVAL_64) begin
      _EVAL_9449 <= 1'h0;
    end else begin
      _EVAL_9449 <= _EVAL_4688;
    end
    if (_EVAL_8339) begin
      if (~_EVAL_15768) begin
        _EVAL_9510 <= _EVAL_13139;
      end
    end
    if (_EVAL_16030) begin
      _EVAL_10347 <= _EVAL_51;
    end else if (_EVAL_17211) begin
      _EVAL_10347 <= csr__EVAL_85;
    end else if (_EVAL_639) begin
      if (_EVAL_19529) begin
        _EVAL_10347 <= csr__EVAL_85;
      end else if (_EVAL_5146) begin
        _EVAL_10347 <= fetch__EVAL_21;
      end else begin
        _EVAL_10347 <= _EVAL_5622;
      end
    end
    if (_EVAL_9061) begin
      _EVAL_10353 <= _EVAL_14920;
    end
    if (_EVAL_3611) begin
      _EVAL_10468 <= _EVAL_3607;
    end
    if (_EVAL_16647) begin
      _EVAL_10593 <= _EVAL_7156;
    end
    if (_EVAL_3611) begin
      _EVAL_10894 <= _EVAL_6400;
    end
    if (_EVAL_64) begin
      _EVAL_11162 <= 1'h0;
    end else if (_EVAL_13371) begin
      if (~_EVAL_1801) begin
        _EVAL_11162 <= 1'h0;
      end else if (_EVAL_8339) begin
        _EVAL_11162 <= _EVAL_18247;
      end
    end else if (_EVAL_8339) begin
      _EVAL_11162 <= _EVAL_18247;
    end
    if (_EVAL_8339) begin
      if (_EVAL_15768) begin
        _EVAL_12371 <= _EVAL_13139;
      end
    end
    if (_EVAL_8339) begin
      if (~_EVAL_15768) begin
        _EVAL_12379 <= _EVAL_3117;
      end
    end
    if (_EVAL_16647) begin
      _EVAL_12498 <= _EVAL_10371;
    end
    if (_EVAL_8339) begin
      if (~_EVAL_15768) begin
        _EVAL_12508 <= _EVAL_10111;
      end
    end
    if (_EVAL_6270) begin
      _EVAL_12724 <= _EVAL_16768;
    end else if (_EVAL_3741) begin
      _EVAL_12724 <= 32'h0;
    end else begin
      _EVAL_12724 <= rf__EVAL_0;
    end
    _EVAL_13327 <= csr__EVAL_84;
    if (_EVAL_8339) begin
      if (_EVAL_15768) begin
        _EVAL_14160 <= _EVAL_17140;
      end
    end
    if (_EVAL_16647) begin
      _EVAL_14184 <= _EVAL_15053;
    end
    if (_EVAL_64) begin
      _EVAL_14478 <= 1'h0;
    end else begin
      _EVAL_14478 <= _EVAL_7137;
    end
    if (!(_EVAL_9378)) begin
      if (_EVAL_9429) begin
        _EVAL_14896 <= _EVAL_10353;
      end else if (_EVAL_5512) begin
        _EVAL_14896 <= _EVAL_14920;
      end
    end
    _EVAL_15545 <= fetch__EVAL_2;
    if (_EVAL_64) begin
      _EVAL_15759 <= 1'h0;
    end else begin
      _EVAL_15759 <= _EVAL_4090;
    end
    _EVAL_16030 <= _EVAL_64 | _EVAL_15467;
    if (_EVAL_13047) begin
      _EVAL_16096 <= 1'h0;
    end else begin
      _EVAL_16096 <= _EVAL_10051;
    end
    if (_EVAL_9061) begin
      _EVAL_16207 <= _EVAL_10480;
    end
    if (_EVAL_64) begin
      _EVAL_16543 <= 1'h0;
    end else begin
      _EVAL_16543 <= _EVAL_18942;
    end
    _EVAL_16644 <= csr__EVAL_26;
    if (_EVAL_3611) begin
      _EVAL_16733 <= _EVAL_15768;
    end
    if (!(_EVAL_9378)) begin
      if (_EVAL_9429) begin
        _EVAL_16768 <= _EVAL_16207;
      end else if (_EVAL_5512) begin
        _EVAL_16768 <= _EVAL_10480;
      end
    end
    if (_EVAL_64) begin
      _EVAL_17371 <= 1'h0;
    end else begin
      _EVAL_17371 <= _EVAL_15656;
    end
    if (_EVAL_8339) begin
      _EVAL_17801 <= _EVAL_10928;
    end
    if (_EVAL_17886) begin
      _EVAL_18514 <= _EVAL_15648;
    end else begin
      _EVAL_18514 <= _EVAL_2225;
    end
    if (_EVAL_8339) begin
      if (_EVAL_15768) begin
        _EVAL_19551 <= _EVAL_127;
      end
    end
  end
endmodule
