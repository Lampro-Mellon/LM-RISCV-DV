//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_46_assert(
  input         _EVAL,
  input         _EVAL_0,
  input  [31:0] _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [3:0]  _EVAL_6,
  input  [1:0]  _EVAL_7,
  input  [3:0]  _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [2:0]  _EVAL_14,
  input  [3:0]  _EVAL_15
);
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire [6:0] _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire [5:0] _EVAL_22;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_23;
  reg [3:0] _EVAL_24;
  reg [31:0] _RAND_0;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire [31:0] _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire [5:0] _EVAL_36;
  reg  _EVAL_37;
  reg [31:0] _RAND_1;
  wire [32:0] _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire [32:0] _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire [32:0] _EVAL_49;
  wire [1:0] _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  reg [31:0] _EVAL_53;
  reg [31:0] _RAND_2;
  wire [32:0] _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire [31:0] _EVAL_58;
  wire  _EVAL_59;
  wire [7:0] _EVAL_60;
  wire [5:0] _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_65;
  wire [32:0] _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire [32:0] _EVAL_71;
  wire [32:0] _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire [31:0] _EVAL_79;
  wire  _EVAL_80;
  wire [32:0] _EVAL_81;
  wire  _EVAL_82;
  wire [1:0] _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire [32:0] _EVAL_88;
  wire  _EVAL_90;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire [32:0] _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire [3:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire [1:0] _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire [3:0] _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_119;
  wire [5:0] _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_124;
  wire [7:0] _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire [6:0] _EVAL_130;
  wire  _EVAL_131;
  wire [31:0] _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire [32:0] _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire [1:0] _EVAL_144;
  wire [22:0] _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire [31:0] _EVAL_161;
  wire [7:0] _EVAL_162;
  wire [31:0] _EVAL_163;
  wire  _EVAL_165;
  reg [2:0] _EVAL_166;
  reg [31:0] _RAND_3;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire [32:0] _EVAL_179;
  wire  _EVAL_180;
  wire [32:0] _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire [31:0] _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire [7:0] _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  reg [3:0] _EVAL_195;
  reg [31:0] _RAND_4;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  reg [5:0] _EVAL_200;
  reg [31:0] _RAND_5;
  wire  _EVAL_201;
  reg  _EVAL_202;
  reg [31:0] _RAND_6;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire [3:0] _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  reg  _EVAL_210;
  reg [31:0] _RAND_7;
  reg [1:0] _EVAL_211;
  reg [31:0] _RAND_8;
  wire [6:0] _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire [5:0] _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire [5:0] _EVAL_221;
  wire [31:0] _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire [32:0] _EVAL_229;
  wire  _EVAL_230;
  wire [6:0] _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire [32:0] _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  reg [31:0] _EVAL_241;
  reg [31:0] _RAND_9;
  wire [32:0] _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire [1:0] _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire [32:0] _EVAL_253;
  wire  _EVAL_254;
  wire [3:0] _EVAL_255;
  wire  _EVAL_256;
  reg [2:0] _EVAL_257;
  reg [31:0] _RAND_10;
  wire  _EVAL_258;
  wire  _EVAL_259;
  reg [5:0] _EVAL_260;
  reg [31:0] _RAND_11;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  reg [5:0] _EVAL_267;
  reg [31:0] _RAND_12;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire [22:0] _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire [32:0] _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  reg  _EVAL_280;
  reg [31:0] _RAND_13;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire [32:0] _EVAL_288;
  reg [5:0] _EVAL_289;
  reg [31:0] _RAND_14;
  wire  _EVAL_290;
  wire  _EVAL_291;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_25 = ~_EVAL_131;
  assign _EVAL_229 = $signed(_EVAL_253) & -33'sh1000;
  assign _EVAL_184 = _EVAL_1 ^ 32'h2000000;
  assign _EVAL_263 = _EVAL_173 & _EVAL_204;
  assign _EVAL_174 = _EVAL_3 & _EVAL_183;
  assign _EVAL_40 = $signed(_EVAL_81) == 33'sh0;
  assign _EVAL_22 = _EVAL_130[5:0];
  assign _EVAL_139 = {1'b0,$signed(_EVAL_184)};
  assign _EVAL_131 = _EVAL_198 | _EVAL_9;
  assign _EVAL_179 = $signed(_EVAL_71) & -33'sh2000;
  assign _EVAL_276 = ~_EVAL_258;
  assign _EVAL_279 = _EVAL_11 == 3'h6;
  assign _EVAL_256 = _EVAL_241 < plusarg_reader_out;
  assign _EVAL_18 = _EVAL_5 & _EVAL_239;
  assign _EVAL_196 = _EVAL == _EVAL_202;
  assign _EVAL_46 = _EVAL_1 == _EVAL_53;
  assign _EVAL_235 = _EVAL_47 & _EVAL_193;
  assign _EVAL_206 = _EVAL_250[0];
  assign _EVAL_265 = _EVAL_238 | _EVAL_106;
  assign _EVAL_274 = _EVAL_148 | _EVAL_77;
  assign _EVAL_194 = _EVAL_35 | _EVAL_9;
  assign _EVAL_17 = $signed(_EVAL_49) == 33'sh0;
  assign _EVAL_212 = _EVAL_289 - 6'h1;
  assign _EVAL_255 = _EVAL_8 & _EVAL_207;
  assign _EVAL_259 = _EVAL_261 | _EVAL_124;
  assign _EVAL_63 = _EVAL_201 | _EVAL_280;
  assign _EVAL_134 = _EVAL_27 | _EVAL_51;
  assign _EVAL_159 = ~_EVAL_65;
  assign _EVAL_271 = _EVAL_30 | _EVAL_124;
  assign _EVAL_94 = {1'b0,$signed(_EVAL_161)};
  assign _EVAL_185 = _EVAL_46 | _EVAL_9;
  assign _EVAL_219 = _EVAL_171 | _EVAL_9;
  assign _EVAL_264 = _EVAL_290 | _EVAL_9;
  assign _EVAL_155 = _EVAL_282 | _EVAL_9;
  assign _EVAL_268 = _EVAL_3 & _EVAL_78;
  assign _EVAL_65 = _EVAL_287 | _EVAL_9;
  assign _EVAL_42 = _EVAL_234;
  assign _EVAL_197 = _EVAL_289 == 6'h0;
  assign _EVAL_90 = _EVAL_7 == _EVAL_211;
  assign _EVAL_74 = _EVAL_44 | _EVAL_9;
  assign _EVAL_48 = ~_EVAL;
  assign _EVAL_136 = ~_EVAL_76;
  assign _EVAL_277 = _EVAL_229;
  assign _EVAL_284 = ~_EVAL_74;
  assign _EVAL_163 = _EVAL_1 & _EVAL_28;
  assign _EVAL_114 = {_EVAL_265,_EVAL_251,_EVAL_191,_EVAL_141};
  assign _EVAL_77 = plusarg_reader_out == 32'h0;
  assign _EVAL_232 = ~_EVAL_133;
  assign _EVAL_55 = ~_EVAL_194;
  assign _EVAL_69 = _EVAL_280 | _EVAL_201;
  assign _EVAL_43 = _EVAL_6 <= 4'h8;
  assign _EVAL_182 = _EVAL_273 | _EVAL_9;
  assign _EVAL_251 = _EVAL_238 | _EVAL_246;
  assign _EVAL_190 = ~_EVAL_125;
  assign _EVAL_239 = _EVAL_14 == 3'h4;
  assign _EVAL_154 = _EVAL_14 == 3'h1;
  assign _EVAL_175 = _EVAL_153 & _EVAL_220;
  assign _EVAL_108 = _EVAL_275 | _EVAL_9;
  assign _EVAL_61 = _EVAL_231[5:0];
  assign _EVAL_161 = _EVAL_1 ^ 32'h20000000;
  assign _EVAL_49 = _EVAL_67;
  assign _EVAL_192 = _EVAL_3 & _EVAL_45;
  assign _EVAL_100 = _EVAL_271 | _EVAL_40;
  assign _EVAL_60 = ~_EVAL_162;
  assign _EVAL_176 = _EVAL_158 & _EVAL_209;
  assign _EVAL_193 = _EVAL_1[1];
  assign _EVAL_218 = ~_EVAL_86;
  assign _EVAL_168 = _EVAL_3 & _EVAL_279;
  assign _EVAL_162 = _EVAL_145[7:0];
  assign _EVAL_28 = {{24'd0}, _EVAL_190};
  assign _EVAL_99 = _EVAL_3 & _EVAL_157;
  assign _EVAL_20 = ~_EVAL_169;
  assign _EVAL_171 = _EVAL_134 | _EVAL_101;
  assign _EVAL_85 = _EVAL_6 >= 4'h2;
  assign _EVAL_110 = _EVAL_14 == 3'h5;
  assign _EVAL_244 = _EVAL_201 != _EVAL_206;
  assign _EVAL_150 = _EVAL_85 | _EVAL_70;
  assign _EVAL_128 = _EVAL_153 & _EVAL_263;
  assign _EVAL_275 = _EVAL_2 == _EVAL_37;
  assign _EVAL_58 = _EVAL_1 ^ 32'h80000000;
  assign _EVAL_157 = _EVAL_11 == 3'h5;
  assign _EVAL_249 = _EVAL_0 & _EVAL_3;
  assign _EVAL_243 = ~_EVAL_151;
  assign _EVAL_95 = _EVAL_158 | _EVAL_249;
  assign _EVAL_237 = _EVAL_249 & _EVAL_178;
  assign _EVAL_32 = _EVAL_172 | _EVAL_12;
  assign _EVAL_68 = _EVAL_14 == _EVAL_166;
  assign _EVAL_26 = ~_EVAL_138;
  assign _EVAL_266 = _EVAL_5 & _EVAL_154;
  assign _EVAL_87 = _EVAL_15 >= 4'h2;
  assign _EVAL_38 = $signed(_EVAL_139) & -33'sh1000000;
  assign _EVAL_252 = _EVAL_11 == 3'h2;
  assign _EVAL_133 = _EVAL_227 | _EVAL_9;
  assign _EVAL_213 = _EVAL_6 == _EVAL_195;
  assign _EVAL_30 = $signed(_EVAL_42) == 33'sh0;
  assign _EVAL_21 = _EVAL_259 | _EVAL_40;
  assign _EVAL_207 = ~_EVAL_114;
  assign _EVAL_209 = _EVAL_260 == 6'h0;
  assign _EVAL_73 = _EVAL_11 == 3'h0;
  assign _EVAL_247 = _EVAL_5 & _EVAL_93;
  assign _EVAL_98 = _EVAL_122 | _EVAL_9;
  assign _EVAL_285 = ~_EVAL_219;
  assign _EVAL_31 = _EVAL_112 | _EVAL_9;
  assign _EVAL_201 = _EVAL_50[0];
  assign _EVAL_148 = ~_EVAL_280;
  assign _EVAL_35 = _EVAL_15 == _EVAL_24;
  assign _EVAL_27 = _EVAL_137 & _EVAL_281;
  assign _EVAL_230 = ~_EVAL_185;
  assign _EVAL_67 = $signed(_EVAL_94) & -33'sh2000;
  assign _EVAL_165 = _EVAL_237 & _EVAL_199;
  assign _EVAL_81 = _EVAL_54;
  assign _EVAL_33 = _EVAL_172 | _EVAL_9;
  assign _EVAL_19 = _EVAL_260 - 6'h1;
  assign _EVAL_51 = _EVAL_117 & _EVAL_278;
  assign _EVAL_222 = _EVAL_88[31:0];
  assign _EVAL_142 = ~_EVAL_31;
  assign _EVAL_96 = _EVAL_269 | _EVAL_9;
  assign _EVAL_145 = 23'hff << _EVAL_15;
  assign _EVAL_129 = _EVAL_59 | _EVAL_9;
  assign _EVAL_39 = _EVAL_116 | _EVAL_9;
  assign _EVAL_203 = _EVAL_51 | _EVAL_101;
  assign _EVAL_269 = _EVAL_7 <= 2'h2;
  assign _EVAL_103 = ~_EVAL_8;
  assign _EVAL_167 = _EVAL_121 | _EVAL_9;
  assign _EVAL_188 = _EVAL_249 & _EVAL_186;
  assign _EVAL_160 = _EVAL_48 | _EVAL_9;
  assign _EVAL_125 = _EVAL_270[7:0];
  assign _EVAL_187 = _EVAL_11[0];
  assign _EVAL_121 = _EVAL_255 == 4'h0;
  assign _EVAL_225 = _EVAL_158 & _EVAL_197;
  assign _EVAL_227 = _EVAL_137 & _EVAL_126;
  assign _EVAL_158 = _EVAL_13 & _EVAL_5;
  assign _EVAL_270 = 23'hff << _EVAL_6;
  assign _EVAL_16 = _EVAL_137 & _EVAL_17;
  assign _EVAL_92 = _EVAL_137 & _EVAL_100;
  assign _EVAL_116 = _EVAL_274 | _EVAL_256;
  assign _EVAL_62 = _EVAL_11 == _EVAL_257;
  assign _EVAL_221 = _EVAL_190[7:2];
  assign _EVAL_41 = _EVAL_90 | _EVAL_9;
  assign _EVAL_278 = $signed(_EVAL_242) == 33'sh0;
  assign _EVAL_82 = _EVAL_148 | _EVAL_9;
  assign _EVAL_57 = ~_EVAL_155;
  assign _EVAL_189 = _EVAL_5 & _EVAL_105;
  assign _EVAL_215 = ~_EVAL_52;
  assign _EVAL_258 = _EVAL_224 | _EVAL_9;
  assign _EVAL_105 = _EVAL_14 == 3'h3;
  assign _EVAL_205 = _EVAL_14 == 3'h0;
  assign _EVAL_169 = _EVAL_68 | _EVAL_9;
  assign _EVAL_117 = _EVAL_6 <= 4'h6;
  assign _EVAL_199 = ~_EVAL_279;
  assign _EVAL_262 = ~_EVAL_264;
  assign _EVAL_254 = _EVAL_3 & _EVAL_73;
  assign _EVAL_253 = {1'b0,$signed(_EVAL_79)};
  assign _EVAL_80 = _EVAL_1[0];
  assign _EVAL_204 = ~_EVAL_80;
  assign _EVAL_178 = _EVAL_200 == 6'h0;
  assign _EVAL_233 = _EVAL_203 | _EVAL_16;
  assign _EVAL_88 = _EVAL_241 + 32'h1;
  assign _EVAL_246 = _EVAL_153 & _EVAL_143;
  assign _EVAL_214 = ~_EVAL_201;
  assign _EVAL_101 = _EVAL_43 & _EVAL_261;
  assign _EVAL_56 = _EVAL_3 & _EVAL_252;
  assign _EVAL_290 = _EVAL_7 != 2'h2;
  assign _EVAL_186 = _EVAL_267 == 6'h0;
  assign _EVAL_152 = _EVAL_5 & _EVAL_177;
  assign _EVAL_130 = _EVAL_200 - 6'h1;
  assign _EVAL_93 = ~_EVAL_197;
  assign _EVAL_141 = _EVAL_150 | _EVAL_128;
  assign _EVAL_111 = 2'h1 << _EVAL_223;
  assign _EVAL_273 = _EVAL_11 <= 3'h6;
  assign _EVAL_138 = _EVAL_213 | _EVAL_9;
  assign _EVAL_181 = {1'b0,$signed(_EVAL_1)};
  assign _EVAL_144 = _EVAL_111 | 2'h1;
  assign _EVAL_47 = _EVAL_144[1];
  assign _EVAL_217 = _EVAL_212[5:0];
  assign _EVAL_78 = ~_EVAL_186;
  assign _EVAL_59 = ~_EVAL_12;
  assign _EVAL_238 = _EVAL_85 | _EVAL_235;
  assign _EVAL_170 = ~_EVAL_206;
  assign _EVAL_172 = ~_EVAL_4;
  assign _EVAL_29 = _EVAL_14 == 3'h6;
  assign _EVAL_198 = _EVAL_7 == 2'h0;
  assign _EVAL_151 = _EVAL_119 | _EVAL_9;
  assign _EVAL_23 = ~_EVAL_160;
  assign _EVAL_124 = $signed(_EVAL_72) == 33'sh0;
  assign _EVAL_231 = _EVAL_267 - 6'h1;
  assign _EVAL_261 = $signed(_EVAL_277) == 33'sh0;
  assign _EVAL_224 = _EVAL_103 == 4'h0;
  assign _EVAL_220 = _EVAL_173 & _EVAL_80;
  assign _EVAL_286 = _EVAL_87 | _EVAL_9;
  assign _EVAL_75 = ~_EVAL_41;
  assign _EVAL_191 = _EVAL_150 | _EVAL_175;
  assign _EVAL_248 = ~_EVAL_182;
  assign _EVAL_208 = ~_EVAL_33;
  assign _EVAL_71 = {1'b0,$signed(_EVAL_132)};
  assign _EVAL_149 = ~_EVAL_98;
  assign _EVAL_120 = _EVAL_60[7:2];
  assign _EVAL_240 = _EVAL_5 & _EVAL_110;
  assign _EVAL_282 = _EVAL_163 == 32'h0;
  assign _EVAL_177 = _EVAL_14 == 3'h7;
  assign _EVAL_236 = ~_EVAL_245;
  assign _EVAL_34 = ~_EVAL_108;
  assign _EVAL_234 = $signed(_EVAL_288) & -33'shc000;
  assign _EVAL_50 = _EVAL_176 ? 2'h1 : 2'h0;
  assign _EVAL_137 = _EVAL_6 <= 4'h2;
  assign _EVAL_226 = ~_EVAL_286;
  assign _EVAL_84 = ~_EVAL_82;
  assign _EVAL_180 = _EVAL_14 == 3'h2;
  assign _EVAL_115 = ~_EVAL_9;
  assign _EVAL_102 = _EVAL_5 & _EVAL_29;
  assign _EVAL_183 = _EVAL_11 == 3'h1;
  assign _EVAL_106 = _EVAL_153 & _EVAL_147;
  assign _EVAL_54 = $signed(_EVAL_181) & -33'sh5000;
  assign _EVAL_122 = _EVAL_244 | _EVAL_214;
  assign _EVAL_250 = _EVAL_165 ? _EVAL_83 : 2'h0;
  assign _EVAL_83 = 2'h1 << _EVAL;
  assign _EVAL_291 = ~_EVAL_129;
  assign _EVAL_242 = _EVAL_179;
  assign _EVAL_156 = ~_EVAL_113;
  assign _EVAL_143 = _EVAL_193 & _EVAL_204;
  assign _EVAL_173 = ~_EVAL_193;
  assign _EVAL_223 = _EVAL_6[0];
  assign _EVAL_44 = _EVAL_92 | _EVAL_101;
  assign _EVAL_97 = _EVAL_69 & _EVAL_170;
  assign _EVAL_86 = _EVAL_14[2];
  assign _EVAL_153 = _EVAL_144[0];
  assign _EVAL_283 = ~_EVAL_167;
  assign _EVAL_70 = _EVAL_47 & _EVAL_173;
  assign _EVAL_245 = _EVAL_196 | _EVAL_9;
  assign _EVAL_287 = _EVAL_4 == _EVAL_210;
  assign _EVAL_132 = _EVAL_1 ^ 32'h40000000;
  assign _EVAL_147 = _EVAL_193 & _EVAL_80;
  assign _EVAL_109 = _EVAL_5 & _EVAL_180;
  assign _EVAL_107 = _EVAL_5 & _EVAL_205;
  assign _EVAL_281 = _EVAL_100 | _EVAL_17;
  assign _EVAL_72 = _EVAL_38;
  assign _EVAL_288 = {1'b0,$signed(_EVAL_58)};
  assign _EVAL_146 = ~_EVAL_216;
  assign _EVAL_45 = _EVAL_11 == 3'h4;
  assign _EVAL_140 = ~_EVAL_96;
  assign _EVAL_36 = _EVAL_19[5:0];
  assign _EVAL_104 = ~_EVAL_39;
  assign _EVAL_113 = _EVAL_62 | _EVAL_9;
  assign _EVAL_119 = _EVAL_63 >> _EVAL;
  assign _EVAL_76 = _EVAL_32 | _EVAL_9;
  assign _EVAL_112 = _EVAL_8 == _EVAL_114;
  assign _EVAL_52 = _EVAL_85 | _EVAL_9;
  assign _EVAL_216 = _EVAL_233 | _EVAL_9;
  assign _EVAL_79 = _EVAL_1 ^ 32'h3000;
  assign _EVAL_126 = _EVAL_21 | _EVAL_17;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_24 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_37 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_53 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_166 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_195 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_200 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_202 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_210 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_211 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_241 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_257 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_260 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_267 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_280 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_289 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_10) begin
    if (_EVAL_188) begin
      _EVAL_24 <= _EVAL_15;
    end
    if (_EVAL_188) begin
      _EVAL_37 <= _EVAL_2;
    end
    if (_EVAL_225) begin
      _EVAL_53 <= _EVAL_1;
    end
    if (_EVAL_225) begin
      _EVAL_166 <= _EVAL_14;
    end
    if (_EVAL_225) begin
      _EVAL_195 <= _EVAL_6;
    end
    if (_EVAL_9) begin
      _EVAL_200 <= 6'h0;
    end else if (_EVAL_249) begin
      if (_EVAL_178) begin
        if (_EVAL_187) begin
          _EVAL_200 <= _EVAL_120;
        end else begin
          _EVAL_200 <= 6'h0;
        end
      end else begin
        _EVAL_200 <= _EVAL_22;
      end
    end
    if (_EVAL_188) begin
      _EVAL_202 <= _EVAL;
    end
    if (_EVAL_188) begin
      _EVAL_210 <= _EVAL_4;
    end
    if (_EVAL_188) begin
      _EVAL_211 <= _EVAL_7;
    end
    if (_EVAL_9) begin
      _EVAL_241 <= 32'h0;
    end else if (_EVAL_95) begin
      _EVAL_241 <= 32'h0;
    end else begin
      _EVAL_241 <= _EVAL_222;
    end
    if (_EVAL_188) begin
      _EVAL_257 <= _EVAL_11;
    end
    if (_EVAL_9) begin
      _EVAL_260 <= 6'h0;
    end else if (_EVAL_158) begin
      if (_EVAL_209) begin
        if (_EVAL_218) begin
          _EVAL_260 <= _EVAL_221;
        end else begin
          _EVAL_260 <= 6'h0;
        end
      end else begin
        _EVAL_260 <= _EVAL_36;
      end
    end
    if (_EVAL_9) begin
      _EVAL_267 <= 6'h0;
    end else if (_EVAL_249) begin
      if (_EVAL_186) begin
        if (_EVAL_187) begin
          _EVAL_267 <= _EVAL_120;
        end else begin
          _EVAL_267 <= 6'h0;
        end
      end else begin
        _EVAL_267 <= _EVAL_61;
      end
    end
    if (_EVAL_9) begin
      _EVAL_280 <= 1'h0;
    end else begin
      _EVAL_280 <= _EVAL_97;
    end
    if (_EVAL_9) begin
      _EVAL_289 <= 6'h0;
    end else if (_EVAL_158) begin
      if (_EVAL_197) begin
        if (_EVAL_218) begin
          _EVAL_289 <= _EVAL_221;
        end else begin
          _EVAL_289 <= 6'h0;
        end
      end else begin
        _EVAL_289 <= _EVAL_217;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5942d6d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50c505b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(450d0da8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9da5e44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2872fe00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ec653e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af7afdc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5648994b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22ed4b70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33a8f0da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c15d74f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0d27379)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3aa6af1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acbf4c9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b4816a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(339bf430)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(657847d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f08bef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61618f1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b8b9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a590fcf5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7da474dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7e60bb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_3 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_149) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40632d74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5757adc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a919e41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(924e0efa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9c14acd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7530587)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff54f275)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57e34b63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_284) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(494503c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(629d8356)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15d79730)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e40bbbf6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a4ce842)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f6280f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2e3ba4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7f49dd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75dcb2f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd44d8d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c92f39a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2034838c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be686a00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e4f9fc4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6190c07c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf46123)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cc50ac6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5663f248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a82b11ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fa12848)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7f4b122)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3ca29d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a9cb649)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bf57c3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9748143b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c509b289)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(674fd831)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfc6c14d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e604ef03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b5eb294)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77120798)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2181f2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ed214b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_284) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b07d5c58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(449ce347)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8918395)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db7901dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e637b13d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
