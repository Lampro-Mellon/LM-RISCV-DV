//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_4_assert(
  input         _EVAL_0,
  input  [3:0]  _EVAL_7,
  input         _EVAL_14,
  input         _EVAL_28,
  input         _EVAL_45,
  input         _EVAL_48,
  input  [31:0] _EVAL_50,
  input  [3:0]  _EVAL_52,
  input  [31:0] _EVAL_58,
  input  [3:0]  _EVAL_61,
  input         _EVAL_69,
  input  [2:0]  _EVAL_79,
  input  [2:0]  _EVAL_86,
  input  [2:0]  _EVAL_87,
  input  [2:0]  _EVAL_89,
  input         _EVAL_91,
  input         _EVAL_97,
  input  [3:0]  _EVAL_115,
  input  [3:0]  _EVAL_120,
  input         _EVAL_122,
  input         _EVAL_125,
  input  [2:0]  _EVAL_128,
  input  [2:0]  _EVAL_135,
  input  [31:0] _EVAL_136,
  input  [3:0]  _EVAL_141,
  input         _EVAL_154,
  input         _EVAL_155,
  input         _EVAL_162,
  input         _EVAL_163,
  input         _EVAL_176,
  input         _EVAL_205,
  input         _EVAL_226,
  input         _EVAL_249,
  input         _EVAL_258,
  input         _EVAL_271,
  input  [2:0]  _EVAL_286,
  input         _EVAL_291,
  input         _EVAL_300,
  input         _EVAL_354,
  input         _EVAL_358,
  input         _EVAL_359,
  input         _EVAL_363,
  input         _EVAL_378,
  input  [46:0] _EVAL_466,
  input         _EVAL_473,
  input         _EVAL_481,
  input         _EVAL_487,
  input         _EVAL_497,
  input         _EVAL_509,
  input         _EVAL_512,
  input         _EVAL_541,
  input         _EVAL_545,
  input         _EVAL_577,
  input         _EVAL_617,
  input         _EVAL_636,
  input  [46:0] _EVAL_691,
  input         _EVAL_701,
  input         _EVAL_709,
  input         _EVAL_755,
  input  [2:0]  _EVAL_759,
  input         _EVAL_768,
  input         _EVAL_802,
  input         _EVAL_803,
  input  [46:0] _EVAL_836,
  input         _EVAL_846,
  input         _EVAL_866,
  input         _EVAL_881,
  input         _EVAL_882,
  input         _EVAL_883,
  input         _EVAL_900,
  input         _EVAL_915,
  input         _EVAL_923,
  input         _EVAL_934,
  input         _EVAL_940,
  input         _EVAL_964,
  input         _EVAL_988,
  input         _EVAL_1025
);
  wire  _EVAL_166;
  wire  _EVAL_172;
  wire  _EVAL_182;
  wire  _EVAL_189;
  wire  _EVAL_191;
  wire  _EVAL_194;
  wire  _EVAL_215;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_229;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_272;
  wire [3:0] TLMonitor__EVAL;
  wire [3:0] TLMonitor__EVAL_0;
  wire [31:0] TLMonitor__EVAL_1;
  wire  TLMonitor__EVAL_2;
  wire [2:0] TLMonitor__EVAL_3;
  wire  TLMonitor__EVAL_4;
  wire  TLMonitor__EVAL_5;
  wire  TLMonitor__EVAL_6;
  wire [3:0] TLMonitor__EVAL_7;
  wire  TLMonitor__EVAL_8;
  wire  TLMonitor__EVAL_9;
  wire  TLMonitor__EVAL_10;
  wire  TLMonitor__EVAL_11;
  wire [1:0] TLMonitor__EVAL_12;
  wire  TLMonitor__EVAL_13;
  wire  TLMonitor__EVAL_14;
  wire [2:0] TLMonitor__EVAL_15;
  wire  TLMonitor__EVAL_16;
  wire [2:0] TLMonitor__EVAL_17;
  wire  TLMonitor__EVAL_18;
  wire  _EVAL_287;
  wire  _EVAL_293;
  wire  _EVAL_302;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_308;
  wire  _EVAL_317;
  wire  _EVAL_335;
  wire  _EVAL_336;
  wire  _EVAL_337;
  wire  _EVAL_339;
  wire  _EVAL_350;
  wire  _EVAL_352;
  wire  _EVAL_360;
  wire  _EVAL_365;
  wire  _EVAL_372;
  wire  _EVAL_390;
  wire  _EVAL_395;
  wire  _EVAL_400;
  wire  _EVAL_407;
  wire  _EVAL_412;
  wire  _EVAL_419;
  wire  _EVAL_423;
  wire  _EVAL_426;
  wire  _EVAL_428;
  wire [3:0] TLMonitor_1__EVAL;
  wire [3:0] TLMonitor_1__EVAL_0;
  wire [31:0] TLMonitor_1__EVAL_1;
  wire  TLMonitor_1__EVAL_2;
  wire [2:0] TLMonitor_1__EVAL_3;
  wire  TLMonitor_1__EVAL_4;
  wire  TLMonitor_1__EVAL_5;
  wire  TLMonitor_1__EVAL_6;
  wire [3:0] TLMonitor_1__EVAL_7;
  wire  TLMonitor_1__EVAL_8;
  wire  TLMonitor_1__EVAL_9;
  wire  TLMonitor_1__EVAL_10;
  wire  TLMonitor_1__EVAL_11;
  wire [1:0] TLMonitor_1__EVAL_12;
  wire  TLMonitor_1__EVAL_13;
  wire  TLMonitor_1__EVAL_14;
  wire [2:0] TLMonitor_1__EVAL_15;
  wire  TLMonitor_1__EVAL_16;
  wire [2:0] TLMonitor_1__EVAL_17;
  wire  TLMonitor_1__EVAL_18;
  wire  _EVAL_431;
  wire  _EVAL_436;
  wire  _EVAL_445;
  wire  _EVAL_446;
  wire  _EVAL_449;
  wire  _EVAL_475;
  wire  _EVAL_484;
  wire  _EVAL_505;
  wire  _EVAL_521;
  wire  _EVAL_533;
  wire  _EVAL_535;
  wire  _EVAL_547;
  wire  _EVAL_549;
  wire  _EVAL_556;
  wire  _EVAL_561;
  wire  _EVAL_576;
  wire  _EVAL_581;
  wire  _EVAL_582;
  wire  _EVAL_588;
  wire  _EVAL_589;
  wire  _EVAL_591;
  wire  _EVAL_604;
  wire  _EVAL_647;
  wire  _EVAL_663;
  wire  _EVAL_688;
  wire  _EVAL_692;
  wire  _EVAL_699;
  wire  _EVAL_713;
  wire  _EVAL_719;
  wire  _EVAL_725;
  wire  _EVAL_734;
  wire  _EVAL_736;
  wire  _EVAL_741;
  wire  _EVAL_745;
  wire  _EVAL_748;
  wire  _EVAL_764;
  wire  _EVAL_774;
  wire  _EVAL_775;
  wire  _EVAL_780;
  wire  _EVAL_782;
  wire  _EVAL_795;
  wire  _EVAL_800;
  wire  _EVAL_801;
  wire  _EVAL_807;
  wire  _EVAL_812;
  wire  _EVAL_815;
  wire  _EVAL_816;
  wire  _EVAL_827;
  wire  _EVAL_831;
  wire  _EVAL_844;
  wire  _EVAL_856;
  wire  _EVAL_858;
  wire  _EVAL_864;
  wire  _EVAL_867;
  wire  _EVAL_873;
  wire  _EVAL_875;
  wire  _EVAL_880;
  wire  _EVAL_897;
  wire  _EVAL_902;
  wire  _EVAL_910;
  wire  _EVAL_913;
  wire  _EVAL_916;
  wire  TLMonitor_2__EVAL;
  wire  TLMonitor_2__EVAL_0;
  wire  TLMonitor_2__EVAL_1;
  wire [2:0] TLMonitor_2__EVAL_2;
  wire  TLMonitor_2__EVAL_3;
  wire [31:0] TLMonitor_2__EVAL_4;
  wire  TLMonitor_2__EVAL_5;
  wire [1:0] TLMonitor_2__EVAL_6;
  wire [2:0] TLMonitor_2__EVAL_7;
  wire  TLMonitor_2__EVAL_8;
  wire [3:0] TLMonitor_2__EVAL_9;
  wire [3:0] TLMonitor_2__EVAL_10;
  wire  TLMonitor_2__EVAL_11;
  wire [2:0] TLMonitor_2__EVAL_12;
  wire  TLMonitor_2__EVAL_13;
  wire  TLMonitor_2__EVAL_14;
  wire  TLMonitor_2__EVAL_15;
  wire  TLMonitor_2__EVAL_16;
  wire [3:0] TLMonitor_2__EVAL_17;
  wire  _EVAL_928;
  wire  _EVAL_930;
  wire  _EVAL_933;
  wire  _EVAL_935;
  wire  _EVAL_948;
  wire  _EVAL_949;
  wire  _EVAL_956;
  wire  _EVAL_970;
  wire  _EVAL_974;
  wire  _EVAL_980;
  wire  _EVAL_986;
  wire  _EVAL_987;
  wire  _EVAL_994;
  wire  _EVAL_1005;
  wire  _EVAL_1007;
  wire  _EVAL_1015;
  wire  _EVAL_1019;
  wire  _EVAL_1020;
  _EVAL_2_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14),
    ._EVAL_15(TLMonitor__EVAL_15),
    ._EVAL_16(TLMonitor__EVAL_16),
    ._EVAL_17(TLMonitor__EVAL_17),
    ._EVAL_18(TLMonitor__EVAL_18)
  );
  _EVAL_2_assert TLMonitor_1 (
    ._EVAL(TLMonitor_1__EVAL),
    ._EVAL_0(TLMonitor_1__EVAL_0),
    ._EVAL_1(TLMonitor_1__EVAL_1),
    ._EVAL_2(TLMonitor_1__EVAL_2),
    ._EVAL_3(TLMonitor_1__EVAL_3),
    ._EVAL_4(TLMonitor_1__EVAL_4),
    ._EVAL_5(TLMonitor_1__EVAL_5),
    ._EVAL_6(TLMonitor_1__EVAL_6),
    ._EVAL_7(TLMonitor_1__EVAL_7),
    ._EVAL_8(TLMonitor_1__EVAL_8),
    ._EVAL_9(TLMonitor_1__EVAL_9),
    ._EVAL_10(TLMonitor_1__EVAL_10),
    ._EVAL_11(TLMonitor_1__EVAL_11),
    ._EVAL_12(TLMonitor_1__EVAL_12),
    ._EVAL_13(TLMonitor_1__EVAL_13),
    ._EVAL_14(TLMonitor_1__EVAL_14),
    ._EVAL_15(TLMonitor_1__EVAL_15),
    ._EVAL_16(TLMonitor_1__EVAL_16),
    ._EVAL_17(TLMonitor_1__EVAL_17),
    ._EVAL_18(TLMonitor_1__EVAL_18)
  );
  _EVAL_3_assert TLMonitor_2 (
    ._EVAL(TLMonitor_2__EVAL),
    ._EVAL_0(TLMonitor_2__EVAL_0),
    ._EVAL_1(TLMonitor_2__EVAL_1),
    ._EVAL_2(TLMonitor_2__EVAL_2),
    ._EVAL_3(TLMonitor_2__EVAL_3),
    ._EVAL_4(TLMonitor_2__EVAL_4),
    ._EVAL_5(TLMonitor_2__EVAL_5),
    ._EVAL_6(TLMonitor_2__EVAL_6),
    ._EVAL_7(TLMonitor_2__EVAL_7),
    ._EVAL_8(TLMonitor_2__EVAL_8),
    ._EVAL_9(TLMonitor_2__EVAL_9),
    ._EVAL_10(TLMonitor_2__EVAL_10),
    ._EVAL_11(TLMonitor_2__EVAL_11),
    ._EVAL_12(TLMonitor_2__EVAL_12),
    ._EVAL_13(TLMonitor_2__EVAL_13),
    ._EVAL_14(TLMonitor_2__EVAL_14),
    ._EVAL_15(TLMonitor_2__EVAL_15),
    ._EVAL_16(TLMonitor_2__EVAL_16),
    ._EVAL_17(TLMonitor_2__EVAL_17)
  );
  assign TLMonitor__EVAL_3 = _EVAL_691[46:44];
  assign _EVAL_774 = ~_EVAL_339;
  assign TLMonitor__EVAL_9 = _EVAL_28;
  assign TLMonitor_1__EVAL_0 = _EVAL_115;
  assign TLMonitor__EVAL_12 = _EVAL_691[43:42];
  assign TLMonitor_2__EVAL = _EVAL_125;
  assign TLMonitor__EVAL_1 = _EVAL_136;
  assign _EVAL_928 = _EVAL_782 | _EVAL_154;
  assign _EVAL_352 = _EVAL_335 & _EVAL_426;
  assign _EVAL_719 = _EVAL_352 | _EVAL_154;
  assign TLMonitor_1__EVAL_8 = _EVAL_836[33];
  assign _EVAL_827 = _EVAL_795 | _EVAL_755;
  assign _EVAL_948 = ~_EVAL_800;
  assign _EVAL_407 = ~_EVAL_701;
  assign TLMonitor_1__EVAL_16 = _EVAL_154;
  assign TLMonitor_2__EVAL_3 = _EVAL_466[0];
  assign _EVAL_734 = _EVAL_774 | _EVAL_449;
  assign _EVAL_604 = _EVAL_218 & _EVAL_994;
  assign _EVAL_816 = ~_EVAL_755;
  assign _EVAL_423 = ~_EVAL_915;
  assign TLMonitor__EVAL_4 = _EVAL_286[0];
  assign _EVAL_930 = ~_EVAL_803;
  assign _EVAL_867 = ~_EVAL_365;
  assign _EVAL_699 = _EVAL_980 | _EVAL_182;
  assign _EVAL_172 = _EVAL_407 | _EVAL_974;
  assign _EVAL_549 = ~_EVAL_795;
  assign TLMonitor__EVAL_11 = _EVAL_122;
  assign _EVAL_949 = ~_EVAL_509;
  assign _EVAL_561 = _EVAL_302 | _EVAL_154;
  assign TLMonitor_2__EVAL_16 = _EVAL_882 | _EVAL_481;
  assign _EVAL_400 = ~_EVAL_484;
  assign TLMonitor__EVAL_15 = _EVAL_86;
  assign TLMonitor_1__EVAL_10 = _EVAL_836[34];
  assign TLMonitor_2__EVAL_17 = _EVAL_61;
  assign _EVAL_1005 = ~_EVAL_272;
  assign _EVAL_916 = _EVAL_336 | _EVAL_556;
  assign TLMonitor_1__EVAL_14 = _EVAL_836[0];
  assign _EVAL_647 = _EVAL_487 | _EVAL_577;
  assign _EVAL_293 = _EVAL_741 | _EVAL_446;
  assign TLMonitor__EVAL_13 = _EVAL_48;
  assign TLMonitor__EVAL = _EVAL_691[41:38];
  assign TLMonitor_1__EVAL_11 = _EVAL_0;
  assign _EVAL_272 = _EVAL_535 | _EVAL_154;
  assign _EVAL_308 = _EVAL_265 & _EVAL_521;
  assign _EVAL_1019 = ~_EVAL_487;
  assign _EVAL_339 = _EVAL_956 | _EVAL_923;
  assign _EVAL_521 = _EVAL_287 | _EVAL_930;
  assign _EVAL_182 = _EVAL_191 | _EVAL_636;
  assign _EVAL_745 = _EVAL_549 | _EVAL_816;
  assign _EVAL_475 = _EVAL_604 | _EVAL_154;
  assign _EVAL_1015 = _EVAL_395 | _EVAL_154;
  assign TLMonitor_1__EVAL_15 = _EVAL_128;
  assign _EVAL_412 = ~_EVAL_768;
  assign TLMonitor_1__EVAL_17 = _EVAL_79;
  assign _EVAL_431 = _EVAL_484 | _EVAL_709;
  assign TLMonitor_1__EVAL_4 = _EVAL_759[0];
  assign TLMonitor_1__EVAL_18 = _EVAL_497 ? _EVAL_701 : _EVAL_541;
  assign TLMonitor_2__EVAL_9 = _EVAL_141;
  assign _EVAL_725 = _EVAL_589 & _EVAL_745;
  assign _EVAL_215 = ~_EVAL_359;
  assign _EVAL_265 = _EVAL_831 | _EVAL_390;
  assign _EVAL_741 = ~_EVAL_258;
  assign TLMonitor__EVAL_18 = _EVAL_940 ? _EVAL_205 : _EVAL_964;
  assign TLMonitor__EVAL_8 = _EVAL_691[33];
  assign _EVAL_317 = ~_EVAL_636;
  assign _EVAL_589 = _EVAL_436 | _EVAL_547;
  assign _EVAL_166 = ~_EVAL_194;
  assign _EVAL_372 = ~_EVAL_473;
  assign _EVAL_194 = _EVAL_172 | _EVAL_154;
  assign TLMonitor_1__EVAL_5 = _EVAL_162;
  assign TLMonitor__EVAL_17 = _EVAL_135;
  assign _EVAL_831 = ~_EVAL_378;
  assign _EVAL_801 = _EVAL_293 | _EVAL_154;
  assign _EVAL_880 = ~_EVAL_577;
  assign _EVAL_780 = ~_EVAL_913;
  assign _EVAL_897 = _EVAL_308 & _EVAL_305;
  assign _EVAL_390 = ~_EVAL_354;
  assign _EVAL_419 = _EVAL_934 | _EVAL_271;
  assign _EVAL_556 = ~_EVAL_176;
  assign TLMonitor_2__EVAL_6 = _EVAL_466[43:42];
  assign TLMonitor__EVAL_6 = _EVAL_883 | _EVAL_363;
  assign _EVAL_336 = ~_EVAL_582;
  assign TLMonitor_1__EVAL_2 = _EVAL_14;
  assign TLMonitor__EVAL_10 = _EVAL_691[34];
  assign _EVAL_713 = _EVAL_400 | _EVAL_237;
  assign _EVAL_970 = _EVAL_229 | _EVAL_154;
  assign TLMonitor_2__EVAL_0 = _EVAL_162;
  assign _EVAL_445 = ~_EVAL_934;
  assign _EVAL_864 = _EVAL_915 | _EVAL_473;
  assign TLMonitor_1__EVAL_1 = _EVAL_58;
  assign _EVAL_902 = ~_EVAL_928;
  assign _EVAL_446 = _EVAL_864 | _EVAL_300;
  assign TLMonitor_1__EVAL = _EVAL_836[41:38];
  assign TLMonitor_1__EVAL_13 = _EVAL_155;
  assign _EVAL_748 = _EVAL_699 | _EVAL_154;
  assign _EVAL_974 = _EVAL_339 | _EVAL_846;
  assign _EVAL_935 = _EVAL_505 | _EVAL_217;
  assign _EVAL_663 = _EVAL_647 | _EVAL_881;
  assign _EVAL_535 = _EVAL_807 | _EVAL_350;
  assign _EVAL_266 = ~_EVAL_475;
  assign TLMonitor__EVAL_2 = _EVAL_69;
  assign TLMonitor_1__EVAL_9 = _EVAL_45;
  assign TLMonitor_2__EVAL_5 = _EVAL_91;
  assign _EVAL_873 = ~_EVAL_512;
  assign _EVAL_844 = ~_EVAL_647;
  assign TLMonitor_2__EVAL_13 = _EVAL_466[33];
  assign _EVAL_428 = _EVAL_445 | _EVAL_588;
  assign _EVAL_337 = ~_EVAL_864;
  assign _EVAL_395 = _EVAL_1020 | _EVAL_663;
  assign TLMonitor_2__EVAL_4 = _EVAL_50;
  assign _EVAL_533 = ~_EVAL_866;
  assign _EVAL_305 = _EVAL_591 | _EVAL_317;
  assign _EVAL_812 = _EVAL_533 | _EVAL_873;
  assign _EVAL_807 = ~_EVAL_900;
  assign _EVAL_217 = ~_EVAL_923;
  assign _EVAL_581 = ~_EVAL_226;
  assign _EVAL_365 = _EVAL_238 | _EVAL_154;
  assign TLMonitor__EVAL_5 = _EVAL_162;
  assign _EVAL_449 = ~_EVAL_846;
  assign _EVAL_591 = ~_EVAL_191;
  assign _EVAL_815 = ~_EVAL_875;
  assign _EVAL_956 = _EVAL_866 | _EVAL_512;
  assign _EVAL_436 = ~_EVAL_249;
  assign TLMonitor_2__EVAL_14 = _EVAL_291 ? _EVAL_900 : _EVAL_988;
  assign TLMonitor_1__EVAL_12 = _EVAL_836[43:42];
  assign _EVAL_688 = _EVAL_428 & _EVAL_360;
  assign _EVAL_764 = ~_EVAL_881;
  assign _EVAL_547 = ~_EVAL_1025;
  assign _EVAL_986 = ~_EVAL_300;
  assign _EVAL_987 = ~_EVAL_748;
  assign _EVAL_910 = ~_EVAL_561;
  assign _EVAL_856 = _EVAL_304 & _EVAL_734;
  assign TLMonitor_1__EVAL_6 = _EVAL_545 | _EVAL_358;
  assign _EVAL_484 = _EVAL_768 | _EVAL_359;
  assign TLMonitor_2__EVAL_11 = _EVAL_466[34];
  assign TLMonitor_2__EVAL_7 = _EVAL_87;
  assign _EVAL_287 = ~_EVAL_736;
  assign TLMonitor__EVAL_14 = _EVAL_691[0];
  assign _EVAL_800 = _EVAL_856 | _EVAL_154;
  assign _EVAL_304 = _EVAL_812 & _EVAL_935;
  assign _EVAL_218 = _EVAL_1019 | _EVAL_880;
  assign _EVAL_229 = _EVAL_581 | _EVAL_431;
  assign _EVAL_795 = _EVAL_249 | _EVAL_1025;
  assign TLMonitor_2__EVAL_10 = _EVAL_466[41:38];
  assign _EVAL_782 = _EVAL_688 & _EVAL_916;
  assign _EVAL_576 = ~_EVAL_719;
  assign TLMonitor__EVAL_0 = _EVAL_7;
  assign TLMonitor_2__EVAL_15 = _EVAL_97;
  assign TLMonitor__EVAL_16 = _EVAL_154;
  assign _EVAL_505 = ~_EVAL_956;
  assign _EVAL_692 = ~_EVAL_617;
  assign TLMonitor_2__EVAL_12 = _EVAL_89;
  assign _EVAL_588 = ~_EVAL_271;
  assign _EVAL_582 = _EVAL_419 | _EVAL_617;
  assign _EVAL_191 = _EVAL_736 | _EVAL_803;
  assign _EVAL_335 = _EVAL_423 | _EVAL_372;
  assign _EVAL_360 = _EVAL_775 | _EVAL_692;
  assign _EVAL_1020 = ~_EVAL_802;
  assign TLMonitor_2__EVAL_1 = _EVAL_163;
  assign _EVAL_858 = _EVAL_412 | _EVAL_215;
  assign _EVAL_913 = _EVAL_897 | _EVAL_154;
  assign TLMonitor_1__EVAL_3 = _EVAL_836[46:44];
  assign _EVAL_994 = _EVAL_844 | _EVAL_764;
  assign _EVAL_1007 = ~_EVAL_1015;
  assign TLMonitor_2__EVAL_8 = _EVAL_154;
  assign _EVAL_302 = _EVAL_949 | _EVAL_827;
  assign _EVAL_426 = _EVAL_337 | _EVAL_986;
  assign _EVAL_933 = ~_EVAL_970;
  assign _EVAL_736 = _EVAL_378 | _EVAL_354;
  assign _EVAL_775 = ~_EVAL_419;
  assign TLMonitor__EVAL_7 = _EVAL_120;
  assign _EVAL_238 = _EVAL_858 & _EVAL_713;
  assign TLMonitor_1__EVAL_7 = _EVAL_52;
  assign _EVAL_875 = _EVAL_725 | _EVAL_154;
  assign _EVAL_189 = ~_EVAL_801;
  assign _EVAL_237 = ~_EVAL_709;
  assign TLMonitor_2__EVAL_2 = _EVAL_466[46:44];
  assign _EVAL_350 = _EVAL_582 | _EVAL_176;
  assign _EVAL_980 = ~_EVAL_205;
  always @(posedge _EVAL_162) begin
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_780) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1007) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_815) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3808bb77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_576) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2658285f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_933) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3808bb77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_902) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_902) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2658285f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3808bb77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_576) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_948) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2658285f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_867) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2658285f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2658285f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_867) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_910) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3808bb77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_987) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1007) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3808bb77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_780) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2658285f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_948) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_933) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_910) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_815) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2658285f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1005) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3808bb77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1005) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_987) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3808bb77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
