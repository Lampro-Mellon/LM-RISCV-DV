//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_58_assert(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input  [29:0] _EVAL_5,
  input         _EVAL_6,
  input  [3:0]  _EVAL_7,
  input  [2:0]  _EVAL_8,
  input  [3:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input  [1:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [3:0]  _EVAL_17,
  input  [2:0]  _EVAL_18
);
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire [7:0] _EVAL_23;
  wire  _EVAL_24;
  wire [5:0] _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire [29:0] _EVAL_28;
  reg [4:0] _EVAL_29;
  reg [31:0] _RAND_0;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire [4:0] _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire [4:0] _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire [5:0] _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire [30:0] _EVAL_41;
  wire [30:0] _EVAL_42;
  reg [5:0] _EVAL_43;
  reg [31:0] _RAND_1;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire [22:0] _EVAL_50;
  wire [7:0] _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  reg [2:0] _EVAL_54;
  reg [31:0] _RAND_2;
  wire  _EVAL_55;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire [5:0] _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire [30:0] _EVAL_65;
  wire [7:0] _EVAL_66;
  wire [7:0] _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire [5:0] _EVAL_73;
  wire  _EVAL_74;
  reg [3:0] _EVAL_75;
  reg [31:0] _RAND_3;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire [5:0] _EVAL_79;
  wire [31:0] plusarg_reader_out;
  wire [30:0] _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire [1:0] _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire [7:0] _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire [4:0] _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire [7:0] _EVAL_113;
  wire  _EVAL_114;
  wire [4:0] _EVAL_115;
  wire [30:0] _EVAL_116;
  wire [31:0] _EVAL_117;
  wire  _EVAL_118;
  reg [3:0] _EVAL_119;
  reg [31:0] _RAND_4;
  wire  _EVAL_120;
  wire  _EVAL_121;
  reg [29:0] _EVAL_122;
  reg [31:0] _RAND_5;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire [30:0] _EVAL_125;
  wire  _EVAL_126;
  wire [29:0] _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire [30:0] _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire [5:0] _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire [6:0] _EVAL_148;
  wire  _EVAL_149;
  wire [30:0] _EVAL_150;
  wire [30:0] _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire [7:0] _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  reg [2:0] _EVAL_162;
  reg [31:0] _RAND_6;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire [3:0] _EVAL_169;
  wire [4:0] _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [29:0] _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire [6:0] _EVAL_178;
  wire  _EVAL_179;
  wire [29:0] _EVAL_180;
  wire  _EVAL_181;
  wire [3:0] _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  reg [1:0] _EVAL_185;
  reg [31:0] _RAND_7;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire [32:0] _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_203;
  reg [2:0] _EVAL_204;
  reg [31:0] _RAND_8;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire [1:0] _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_212;
  wire [4:0] _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire [7:0] _EVAL_217;
  wire [6:0] _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  reg [5:0] _EVAL_225;
  reg [31:0] _RAND_9;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  reg [5:0] _EVAL_232;
  reg [31:0] _RAND_10;
  wire [3:0] _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire [22:0] _EVAL_237;
  reg  _EVAL_238;
  reg [31:0] _RAND_11;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  reg  _EVAL_258;
  reg [31:0] _RAND_12;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  reg [5:0] _EVAL_263;
  reg [31:0] _RAND_13;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire [1:0] _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  reg [31:0] _EVAL_274;
  reg [31:0] _RAND_14;
  wire  _EVAL_275;
  reg [2:0] _EVAL_276;
  reg [31:0] _RAND_15;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire [30:0] _EVAL_289;
  reg [2:0] _EVAL_290;
  reg [31:0] _RAND_16;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire [29:0] _EVAL_294;
  wire  _EVAL_295;
  wire [4:0] _EVAL_296;
  wire  _EVAL_297;
  wire [4:0] _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_307;
  wire [30:0] _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire [1:0] _EVAL_312;
  wire [6:0] _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire [30:0] _EVAL_318;
  wire [3:0] _EVAL_319;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_168 = _EVAL_173 & _EVAL_171;
  assign _EVAL_293 = ~_EVAL_2;
  assign _EVAL_206 = _EVAL_184 | _EVAL_14;
  assign _EVAL_242 = _EVAL_84 == 2'h0;
  assign _EVAL_105 = _EVAL_17 >= 4'h2;
  assign _EVAL_141 = ~_EVAL_98;
  assign _EVAL_250 = ~_EVAL_6;
  assign _EVAL_131 = _EVAL_15 & _EVAL_175;
  assign _EVAL_39 = ~_EVAL_85;
  assign _EVAL_59 = _EVAL_17 == _EVAL_119;
  assign _EVAL_146 = _EVAL_205 | _EVAL_282;
  assign _EVAL_86 = _EVAL_11 == _EVAL_238;
  assign _EVAL_157 = ~_EVAL_11;
  assign _EVAL_27 = ~_EVAL_279;
  assign _EVAL_136 = _EVAL_314 & _EVAL_24;
  assign _EVAL_62 = _EVAL_217[7:2];
  assign _EVAL_165 = _EVAL_21 | _EVAL_14;
  assign _EVAL_236 = _EVAL_53 | _EVAL_286;
  assign _EVAL_120 = ~_EVAL_206;
  assign _EVAL_142 = _EVAL_114 | _EVAL_14;
  assign _EVAL_60 = ~_EVAL_44;
  assign _EVAL_291 = _EVAL_15 & _EVAL_307;
  assign _EVAL_271 = _EVAL_312 | 2'h1;
  assign _EVAL_78 = ~_EVAL_207;
  assign _EVAL_198 = ~_EVAL_33;
  assign _EVAL_25 = _EVAL_218[5:0];
  assign _EVAL_177 = ~_EVAL_106;
  assign _EVAL_190 = _EVAL_8 == 3'h4;
  assign _EVAL_184 = _EVAL_12 != 2'h2;
  assign _EVAL_210 = _EVAL_9 == _EVAL_75;
  assign _EVAL_156 = _EVAL_208 == 2'h1;
  assign _EVAL_73 = _EVAL_67[7:2];
  assign _EVAL_314 = _EVAL_216 & _EVAL_310;
  assign _EVAL_123 = _EVAL_222 | _EVAL_186;
  assign _EVAL_124 = _EVAL_3 == 3'h1;
  assign _EVAL_265 = _EVAL_152 | _EVAL_70;
  assign _EVAL_79 = _EVAL_313[5:0];
  assign _EVAL_280 = _EVAL_15 & _EVAL_81;
  assign _EVAL_107 = ~_EVAL_296;
  assign _EVAL_32 = _EVAL_51[4:0];
  assign _EVAL_244 = _EVAL_3 == 3'h6;
  assign _EVAL_68 = _EVAL_154 | _EVAL_14;
  assign _EVAL_50 = 23'hff << _EVAL_9;
  assign _EVAL_117 = _EVAL_194[31:0];
  assign _EVAL_61 = _EVAL_274 < plusarg_reader_out;
  assign _EVAL_275 = ~_EVAL_161;
  assign _EVAL_226 = _EVAL_103 | _EVAL_255;
  assign _EVAL_317 = ~_EVAL_203;
  assign _EVAL_182 = ~_EVAL_169;
  assign _EVAL_167 = _EVAL_263 == 6'h0;
  assign _EVAL_48 = _EVAL_139 & _EVAL_187;
  assign _EVAL_218 = _EVAL_232 - 6'h1;
  assign _EVAL_135 = _EVAL_173 & _EVAL_265;
  assign _EVAL_84 = _EVAL_10[2:1];
  assign _EVAL_212 = ~_EVAL_300;
  assign _EVAL_245 = ~_EVAL_46;
  assign _EVAL_298 = _EVAL_29 | _EVAL_32;
  assign _EVAL_102 = _EVAL_43 == 6'h0;
  assign _EVAL_224 = _EVAL_302 & _EVAL_106;
  assign _EVAL_166 = ~_EVAL_95;
  assign _EVAL_313 = _EVAL_43 - 6'h1;
  assign _EVAL_112 = _EVAL_17 <= 4'h8;
  assign _EVAL_150 = $signed(_EVAL_151) & -31'sh1000000;
  assign _EVAL_20 = ~_EVAL_234;
  assign _EVAL_172 = ~_EVAL_102;
  assign _EVAL_115 = _EVAL_32 | _EVAL_29;
  assign _EVAL_216 = _EVAL_16 & _EVAL_13;
  assign _EVAL_286 = _EVAL_173 & _EVAL_240;
  assign _EVAL_240 = _EVAL_265 | _EVAL_171;
  assign _EVAL_103 = ~_EVAL_259;
  assign _EVAL_256 = ~_EVAL_145;
  assign _EVAL_229 = ~_EVAL_45;
  assign _EVAL_259 = _EVAL_29 != 5'h0;
  assign _EVAL_260 = _EVAL_157 | _EVAL_6;
  assign _EVAL_55 = ~_EVAL_121;
  assign _EVAL_305 = _EVAL_8[2];
  assign _EVAL_151 = {1'b0,$signed(_EVAL_294)};
  assign _EVAL_292 = _EVAL_132 | _EVAL_14;
  assign _EVAL_46 = _EVAL_309 | _EVAL_14;
  assign _EVAL_254 = ~_EVAL_165;
  assign _EVAL_139 = _EVAL_4 & _EVAL_15;
  assign _EVAL_127 = {{22'd0}, _EVAL_217};
  assign _EVAL_159 = _EVAL_50[7:0];
  assign _EVAL_205 = _EVAL_40 | _EVAL_242;
  assign _EVAL_308 = _EVAL_42;
  assign _EVAL_213 = _EVAL_29 >> _EVAL_10;
  assign _EVAL_297 = ~_EVAL_219;
  assign _EVAL_312 = 2'h1 << _EVAL_155;
  assign _EVAL_309 = _EVAL_5 == _EVAL_122;
  assign _EVAL_284 = _EVAL_13 & _EVAL_140;
  assign _EVAL_294 = _EVAL_5 ^ 30'h2000000;
  assign _EVAL_22 = _EVAL_15 & _EVAL_269;
  assign _EVAL_181 = _EVAL_3[0];
  assign _EVAL_174 = _EVAL_5 ^ 30'h20000000;
  assign _EVAL_281 = _EVAL_264 | _EVAL_278;
  assign _EVAL_228 = _EVAL_287 | _EVAL_14;
  assign _EVAL_129 = _EVAL <= 3'h1;
  assign _EVAL_267 = _EVAL <= 3'h4;
  assign _EVAL_132 = _EVAL_8 == _EVAL_290;
  assign _EVAL_262 = $signed(_EVAL_318) == 31'sh0;
  assign _EVAL_128 = ~_EVAL_266;
  assign _EVAL_149 = _EVAL_3 == 3'h4;
  assign _EVAL_287 = _EVAL != 3'h0;
  assign _EVAL_247 = _EVAL_213[0];
  assign _EVAL_282 = _EVAL_10 == 3'h4;
  assign _EVAL_195 = _EVAL_105 | _EVAL_14;
  assign _EVAL_110 = ~_EVAL_215;
  assign _EVAL_66 = 8'h1 << _EVAL_18;
  assign _EVAL_24 = ~_EVAL_244;
  assign _EVAL_121 = _EVAL_147 | _EVAL_14;
  assign _EVAL_140 = _EVAL_3 == 3'h0;
  assign _EVAL_311 = ~_EVAL_305;
  assign _EVAL_169 = {_EVAL_123,_EVAL_99,_EVAL_97,_EVAL_281};
  assign _EVAL_178 = _EVAL_263 - 6'h1;
  assign _EVAL_197 = _EVAL_3 == 3'h2;
  assign _EVAL_35 = _EVAL_298 & _EVAL_107;
  assign _EVAL_230 = _EVAL_18 == 3'h4;
  assign _EVAL_246 = _EVAL_208 == 2'h0;
  assign _EVAL_186 = _EVAL_188 & _EVAL_224;
  assign _EVAL_187 = _EVAL_232 == 6'h0;
  assign _EVAL_176 = _EVAL_283 | _EVAL_14;
  assign _EVAL_97 = _EVAL_264 | _EVAL_315;
  assign _EVAL_268 = ~_EVAL_68;
  assign _EVAL_288 = _EVAL_302 & _EVAL_177;
  assign _EVAL_158 = _EVAL_249 | _EVAL_230;
  assign _EVAL_37 = ~_EVAL_118;
  assign _EVAL_249 = _EVAL_156 | _EVAL_246;
  assign _EVAL_114 = _EVAL_3 == _EVAL_204;
  assign _EVAL_34 = _EVAL_130 | _EVAL_14;
  assign _EVAL_235 = _EVAL_13 & _EVAL_197;
  assign _EVAL_170 = _EVAL_115 >> _EVAL_18;
  assign _EVAL_130 = _EVAL_28 == 30'h0;
  assign _EVAL_278 = _EVAL_188 & _EVAL_100;
  assign _EVAL_101 = _EVAL_86 | _EVAL_14;
  assign _EVAL_164 = _EVAL_15 & _EVAL_76;
  assign _EVAL_45 = _EVAL_146 | _EVAL_14;
  assign _EVAL_301 = _EVAL_8 == 3'h5;
  assign _EVAL_41 = {1'b0,$signed(_EVAL_5)};
  assign _EVAL_180 = _EVAL_5 ^ 30'h3000;
  assign _EVAL_200 = _EVAL_31 | _EVAL_14;
  assign _EVAL_98 = _EVAL_210 | _EVAL_14;
  assign _EVAL_38 = _EVAL_148[5:0];
  assign _EVAL_100 = _EVAL_52 & _EVAL_177;
  assign _EVAL_52 = ~_EVAL_302;
  assign _EVAL_295 = ~_EVAL_239;
  assign _EVAL_108 = ~_EVAL_34;
  assign _EVAL_302 = _EVAL_5[1];
  assign _EVAL_223 = _EVAL_226 | _EVAL_61;
  assign _EVAL_319 = ~_EVAL_7;
  assign _EVAL_215 = _EVAL_199 | _EVAL_14;
  assign _EVAL_83 = _EVAL_18 == _EVAL_162;
  assign _EVAL_36 = ~_EVAL_200;
  assign _EVAL_81 = _EVAL_8 == 3'h7;
  assign _EVAL_145 = _EVAL_26 | _EVAL_14;
  assign _EVAL_77 = _EVAL_0 == _EVAL_258;
  assign _EVAL_58 = _EVAL_3 <= 3'h6;
  assign _EVAL_143 = _EVAL_191 & _EVAL_52;
  assign _EVAL_318 = _EVAL_133;
  assign _EVAL_171 = $signed(_EVAL_125) == 31'sh0;
  assign _EVAL_183 = _EVAL_13 & _EVAL_134;
  assign _EVAL_152 = $signed(_EVAL_116) == 31'sh0;
  assign _EVAL_88 = ~_EVAL_72;
  assign _EVAL_26 = _EVAL_7 == _EVAL_169;
  assign _EVAL_264 = _EVAL_105 | _EVAL_143;
  assign _EVAL_85 = _EVAL_272 | _EVAL_14;
  assign _EVAL_89 = _EVAL_173 & _EVAL_262;
  assign _EVAL_104 = _EVAL_8 == 3'h2;
  assign _EVAL_222 = _EVAL_105 | _EVAL_220;
  assign _EVAL_154 = _EVAL <= 3'h2;
  assign _EVAL_65 = $signed(_EVAL_80) & -31'sh2000;
  assign _EVAL_67 = ~_EVAL_159;
  assign _EVAL_219 = _EVAL_109 | _EVAL_14;
  assign _EVAL_71 = _EVAL_250 | _EVAL_14;
  assign _EVAL_255 = plusarg_reader_out == 32'h0;
  assign _EVAL_42 = $signed(_EVAL_41) & -31'sh5000;
  assign _EVAL_53 = _EVAL_112 & _EVAL_262;
  assign _EVAL_144 = ~_EVAL_64;
  assign _EVAL_199 = _EVAL_12 <= 2'h2;
  assign _EVAL_261 = ~_EVAL_299;
  assign _EVAL_76 = _EVAL_8 == 3'h6;
  assign _EVAL_80 = {1'b0,$signed(_EVAL_174)};
  assign _EVAL_300 = _EVAL_193 | _EVAL_14;
  assign _EVAL_113 = _EVAL_136 ? _EVAL_66 : 8'h0;
  assign _EVAL_233 = _EVAL_7 & _EVAL_182;
  assign _EVAL_188 = _EVAL_271[0];
  assign _EVAL_193 = _EVAL_12 == _EVAL_185;
  assign _EVAL_138 = _EVAL_139 | _EVAL_216;
  assign _EVAL_57 = _EVAL_15 & _EVAL_104;
  assign _EVAL_283 = ~_EVAL_247;
  assign _EVAL_279 = _EVAL_223 | _EVAL_14;
  assign _EVAL_125 = _EVAL_65;
  assign _EVAL_316 = _EVAL_8 == 3'h1;
  assign _EVAL_252 = _EVAL == 3'h0;
  assign _EVAL_173 = _EVAL_17 <= 4'h2;
  assign _EVAL_160 = _EVAL_13 & _EVAL_149;
  assign _EVAL_243 = _EVAL_157 | _EVAL_14;
  assign _EVAL_315 = _EVAL_188 & _EVAL_189;
  assign _EVAL_270 = ~_EVAL_176;
  assign _EVAL_231 = _EVAL_13 & _EVAL_124;
  assign _EVAL_273 = _EVAL_319 == 4'h0;
  assign _EVAL_49 = _EVAL_89 | _EVAL_14;
  assign _EVAL_109 = _EVAL_53 | _EVAL_168;
  assign _EVAL_269 = ~_EVAL_187;
  assign _EVAL_289 = {1'b0,$signed(_EVAL_180)};
  assign _EVAL_189 = _EVAL_52 & _EVAL_106;
  assign _EVAL_93 = _EVAL <= 3'h3;
  assign _EVAL_307 = _EVAL_8 == 3'h0;
  assign _EVAL_28 = _EVAL_5 & _EVAL_127;
  assign _EVAL_99 = _EVAL_222 | _EVAL_201;
  assign _EVAL_116 = _EVAL_150;
  assign _EVAL_194 = _EVAL_274 + 32'h1;
  assign _EVAL_33 = _EVAL_236 | _EVAL_14;
  assign _EVAL_92 = 8'h1 << _EVAL_10;
  assign _EVAL_74 = ~_EVAL_101;
  assign _EVAL_94 = ~_EVAL_251;
  assign _EVAL_82 = _EVAL_13 & _EVAL_172;
  assign _EVAL_63 = ~_EVAL_227;
  assign _EVAL_72 = _EVAL_293 | _EVAL_14;
  assign _EVAL_227 = _EVAL_59 | _EVAL_14;
  assign _EVAL_31 = _EVAL_170[0];
  assign _EVAL_234 = _EVAL_83 | _EVAL_14;
  assign _EVAL_44 = _EVAL_90 | _EVAL_14;
  assign _EVAL_111 = ~_EVAL_14;
  assign _EVAL_221 = _EVAL_15 & _EVAL_301;
  assign _EVAL_106 = _EVAL_5[0];
  assign _EVAL_51 = _EVAL_209 ? _EVAL_92 : 8'h0;
  assign _EVAL_196 = ~_EVAL_243;
  assign _EVAL_253 = ~_EVAL_47;
  assign _EVAL_91 = _EVAL_9 >= 4'h2;
  assign _EVAL_208 = _EVAL_18[2:1];
  assign _EVAL_251 = _EVAL_91 | _EVAL_14;
  assign _EVAL_179 = _EVAL_15 & _EVAL_190;
  assign _EVAL_209 = _EVAL_139 & _EVAL_167;
  assign _EVAL_64 = _EVAL_129 | _EVAL_14;
  assign _EVAL_203 = _EVAL_267 | _EVAL_14;
  assign _EVAL_191 = _EVAL_271[1];
  assign _EVAL_148 = _EVAL_225 - 6'h1;
  assign _EVAL_147 = _EVAL == _EVAL_54;
  assign _EVAL_21 = _EVAL_233 == 4'h0;
  assign _EVAL_30 = _EVAL_10 == _EVAL_276;
  assign _EVAL_90 = _EVAL_53 | _EVAL_135;
  assign _EVAL_272 = _EVAL_12 == 2'h0;
  assign _EVAL_266 = _EVAL_58 | _EVAL_14;
  assign _EVAL_192 = ~_EVAL_71;
  assign _EVAL_201 = _EVAL_188 & _EVAL_288;
  assign _EVAL_133 = $signed(_EVAL_289) & -31'sh1000;
  assign _EVAL_299 = _EVAL_93 | _EVAL_14;
  assign _EVAL_47 = _EVAL_260 | _EVAL_14;
  assign _EVAL_285 = ~_EVAL_228;
  assign _EVAL_23 = _EVAL_237[7:0];
  assign _EVAL_310 = _EVAL_225 == 6'h0;
  assign _EVAL_70 = $signed(_EVAL_308) == 31'sh0;
  assign _EVAL_126 = ~_EVAL_142;
  assign _EVAL_175 = _EVAL_8 == 3'h3;
  assign _EVAL_69 = ~_EVAL_195;
  assign _EVAL_40 = _EVAL_84 == 2'h1;
  assign _EVAL_118 = _EVAL_77 | _EVAL_14;
  assign _EVAL_155 = _EVAL_17[0];
  assign _EVAL_241 = _EVAL_216 & _EVAL_102;
  assign _EVAL_239 = _EVAL_273 | _EVAL_14;
  assign _EVAL_304 = _EVAL_13 & _EVAL_244;
  assign _EVAL_237 = 23'hff << _EVAL_17;
  assign _EVAL_134 = _EVAL_3 == 3'h5;
  assign _EVAL_87 = _EVAL_15 & _EVAL_316;
  assign _EVAL_296 = _EVAL_113[4:0];
  assign _EVAL_217 = ~_EVAL_23;
  assign _EVAL_95 = _EVAL_158 | _EVAL_14;
  assign _EVAL_220 = _EVAL_191 & _EVAL_302;
  assign _EVAL_207 = _EVAL_30 | _EVAL_14;
  assign _EVAL_96 = ~_EVAL_49;
  assign _EVAL_161 = _EVAL_252 | _EVAL_14;
  assign _EVAL_137 = _EVAL_178[5:0];
  assign _EVAL_214 = ~_EVAL_292;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_29 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_43 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_54 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_75 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_119 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_122 = _RAND_5[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_162 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_185 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_204 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_225 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_232 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_238 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_258 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_263 = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_274 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_276 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_290 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_1) begin
    if (_EVAL_14) begin
      _EVAL_29 <= 5'h0;
    end else begin
      _EVAL_29 <= _EVAL_35;
    end
    if (_EVAL_14) begin
      _EVAL_43 <= 6'h0;
    end else if (_EVAL_216) begin
      if (_EVAL_102) begin
        if (_EVAL_181) begin
          _EVAL_43 <= _EVAL_73;
        end else begin
          _EVAL_43 <= 6'h0;
        end
      end else begin
        _EVAL_43 <= _EVAL_79;
      end
    end
    if (_EVAL_48) begin
      _EVAL_54 <= _EVAL;
    end
    if (_EVAL_241) begin
      _EVAL_75 <= _EVAL_9;
    end
    if (_EVAL_48) begin
      _EVAL_119 <= _EVAL_17;
    end
    if (_EVAL_48) begin
      _EVAL_122 <= _EVAL_5;
    end
    if (_EVAL_241) begin
      _EVAL_162 <= _EVAL_18;
    end
    if (_EVAL_241) begin
      _EVAL_185 <= _EVAL_12;
    end
    if (_EVAL_241) begin
      _EVAL_204 <= _EVAL_3;
    end
    if (_EVAL_14) begin
      _EVAL_225 <= 6'h0;
    end else if (_EVAL_216) begin
      if (_EVAL_310) begin
        if (_EVAL_181) begin
          _EVAL_225 <= _EVAL_73;
        end else begin
          _EVAL_225 <= 6'h0;
        end
      end else begin
        _EVAL_225 <= _EVAL_38;
      end
    end
    if (_EVAL_14) begin
      _EVAL_232 <= 6'h0;
    end else if (_EVAL_139) begin
      if (_EVAL_187) begin
        if (_EVAL_311) begin
          _EVAL_232 <= _EVAL_62;
        end else begin
          _EVAL_232 <= 6'h0;
        end
      end else begin
        _EVAL_232 <= _EVAL_25;
      end
    end
    if (_EVAL_241) begin
      _EVAL_238 <= _EVAL_11;
    end
    if (_EVAL_241) begin
      _EVAL_258 <= _EVAL_0;
    end
    if (_EVAL_14) begin
      _EVAL_263 <= 6'h0;
    end else if (_EVAL_139) begin
      if (_EVAL_167) begin
        if (_EVAL_311) begin
          _EVAL_263 <= _EVAL_62;
        end else begin
          _EVAL_263 <= 6'h0;
        end
      end else begin
        _EVAL_263 <= _EVAL_137;
      end
    end
    if (_EVAL_14) begin
      _EVAL_274 <= 32'h0;
    end else if (_EVAL_138) begin
      _EVAL_274 <= 32'h0;
    end else begin
      _EVAL_274 <= _EVAL_117;
    end
    if (_EVAL_48) begin
      _EVAL_276 <= _EVAL_10;
    end
    if (_EVAL_48) begin
      _EVAL_290 <= _EVAL_8;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81ab1b84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_275) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c91a0bb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1743c99a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1efb899)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77977237)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d64ce61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ce9aef3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c083ff5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faf7e6eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b574bc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_275) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5aa13bd3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ebb9939)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fe87ab8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d9e1c5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4269b393)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ac8af54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df4858e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b633091)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c316d4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffeb3334)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(670f841a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90ba03b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7e6cfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(505a0c71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b013734)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f79737c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab9251a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc4eda89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bb99045)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(735fb90f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c27bd29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f26c22c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac6a7ed2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(341d39fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e42c1aa4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfb29309)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90d7a104)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c444d709)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd9cb9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bf9e47a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fedf99bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(578290dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ed1e18b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1372d294)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(398923d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f279574b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6aacce2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cd45ef8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cf4b831)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c087f95e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5655b1ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(345139d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f476a99b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_275) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22eebcbf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6faaecb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f50632dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c541eb72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f599f77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56e82bcd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8769578)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58ab3a7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(514e568f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa6de6ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9663dabe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b8c7cc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8983155d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(388e4651)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdce1346)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26260fdb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(441e8e48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd3239ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe9fdec8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5941dffa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11b6d235)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee1a7b85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9aa78a7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48f8da1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab788afc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ad7b9a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_275) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f66d9247)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_275) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c117bfa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_275) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27d2af5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(474adda0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0d9cb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5d4da15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff0583e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b648dc36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64ee269e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e72b65c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79733141)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
