//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_26(
  output [31:0] _EVAL,
  output        _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [31:0] _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  output        _EVAL_5,
  input         _EVAL_6,
  output [2:0]  _EVAL_7,
  input  [2:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [1:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  output        _EVAL_17,
  input         _EVAL_18,
  input  [31:0] _EVAL_19,
  output [2:0]  _EVAL_20,
  output [2:0]  _EVAL_21,
  input         _EVAL_22,
  output        _EVAL_23,
  output [1:0]  _EVAL_24,
  output [2:0]  _EVAL_25,
  input  [2:0]  _EVAL_26,
  output        _EVAL_27,
  input         _EVAL_28,
  input  [3:0]  _EVAL_29,
  output [2:0]  _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  output [30:0] _EVAL_33,
  output        _EVAL_34,
  output [2:0]  _EVAL_35,
  output        _EVAL_36,
  input  [30:0] _EVAL_37,
  output        _EVAL_38,
  input  [2:0]  _EVAL_39,
  input         _EVAL_40,
  output        _EVAL_41,
  output        _EVAL_42,
  output [31:0] _EVAL_43,
  output        _EVAL_44,
  output [2:0]  _EVAL_45,
  input         _EVAL_46,
  output [3:0]  _EVAL_47,
  output        _EVAL_48
);
  assign _EVAL = _EVAL_19;
  assign _EVAL_34 = _EVAL_16;
  assign _EVAL_23 = _EVAL_15;
  assign _EVAL_24 = _EVAL_11;
  assign _EVAL_47 = _EVAL_29;
  assign _EVAL_35 = _EVAL_10;
  assign _EVAL_30 = _EVAL_4;
  assign _EVAL_38 = _EVAL_40;
  assign _EVAL_42 = _EVAL_13;
  assign _EVAL_7 = _EVAL_39;
  assign _EVAL_45 = _EVAL_1;
  assign _EVAL_21 = _EVAL_8;
  assign _EVAL_48 = _EVAL_31;
  assign _EVAL_25 = _EVAL_9;
  assign _EVAL_43 = _EVAL_2;
  assign _EVAL_0 = _EVAL_12;
  assign _EVAL_17 = _EVAL_14;
  assign _EVAL_44 = _EVAL_6;
  assign _EVAL_20 = _EVAL_26;
  assign _EVAL_5 = _EVAL_18;
  assign _EVAL_33 = _EVAL_37;
  assign _EVAL_36 = _EVAL_46;
  assign _EVAL_27 = _EVAL_3;
  assign _EVAL_41 = _EVAL_28;
endmodule
