//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_66(
  output        _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  output        _EVAL_4,
  input         _EVAL_5,
  output [3:0]  _EVAL_6,
  input         _EVAL_7,
  output [1:0]  _EVAL_8,
  input  [31:0] _EVAL_9,
  input  [1:0]  _EVAL_10,
  output [31:0] _EVAL_11,
  output [2:0]  _EVAL_12,
  input  [3:0]  _EVAL_13,
  output        _EVAL_14,
  output        _EVAL_15,
  output [2:0]  _EVAL_16,
  output        _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  input  [2:0]  _EVAL_20
);
  reg  _EVAL_21 [0:1];
  reg [31:0] _RAND_0;
  wire  _EVAL_21__EVAL_22_data;
  wire  _EVAL_21__EVAL_22_addr;
  wire  _EVAL_21__EVAL_23_data;
  wire  _EVAL_21__EVAL_23_addr;
  wire  _EVAL_21__EVAL_23_mask;
  wire  _EVAL_21__EVAL_23_en;
  wire  _EVAL_24;
  reg [3:0] _EVAL_25 [0:1];
  reg [31:0] _RAND_1;
  wire [3:0] _EVAL_25__EVAL_26_data;
  wire  _EVAL_25__EVAL_26_addr;
  wire [3:0] _EVAL_25__EVAL_27_data;
  wire  _EVAL_25__EVAL_27_addr;
  wire  _EVAL_25__EVAL_27_mask;
  wire  _EVAL_25__EVAL_27_en;
  reg  _EVAL_29;
  reg [31:0] _RAND_2;
  wire  _EVAL_30;
  reg  _EVAL_31;
  reg [31:0] _RAND_3;
  reg  _EVAL_32;
  reg [31:0] _RAND_4;
  wire  _EVAL_34;
  wire  _EVAL_35;
  reg  _EVAL_37 [0:1];
  reg [31:0] _RAND_5;
  wire  _EVAL_37__EVAL_38_data;
  wire  _EVAL_37__EVAL_38_addr;
  wire  _EVAL_37__EVAL_39_data;
  wire  _EVAL_37__EVAL_39_addr;
  wire  _EVAL_37__EVAL_39_mask;
  wire  _EVAL_37__EVAL_39_en;
  reg [2:0] _EVAL_40 [0:1];
  reg [31:0] _RAND_6;
  wire [2:0] _EVAL_40__EVAL_41_data;
  wire  _EVAL_40__EVAL_41_addr;
  wire [2:0] _EVAL_40__EVAL_42_data;
  wire  _EVAL_40__EVAL_42_addr;
  wire  _EVAL_40__EVAL_42_mask;
  wire  _EVAL_40__EVAL_42_en;
  reg [2:0] _EVAL_43 [0:1];
  reg [31:0] _RAND_7;
  wire [2:0] _EVAL_43__EVAL_44_data;
  wire  _EVAL_43__EVAL_44_addr;
  wire [2:0] _EVAL_43__EVAL_45_data;
  wire  _EVAL_43__EVAL_45_addr;
  wire  _EVAL_43__EVAL_45_mask;
  wire  _EVAL_43__EVAL_45_en;
  wire  _EVAL_46;
  wire [1:0] _EVAL_47;
  wire  _EVAL_48;
  reg [1:0] _EVAL_49 [0:1];
  reg [31:0] _RAND_8;
  wire [1:0] _EVAL_49__EVAL_50_data;
  wire  _EVAL_49__EVAL_50_addr;
  wire [1:0] _EVAL_49__EVAL_51_data;
  wire  _EVAL_49__EVAL_51_addr;
  wire  _EVAL_49__EVAL_51_mask;
  wire  _EVAL_49__EVAL_51_en;
  wire  _EVAL_52;
  reg  _EVAL_53 [0:1];
  reg [31:0] _RAND_9;
  wire  _EVAL_53__EVAL_54_data;
  wire  _EVAL_53__EVAL_54_addr;
  wire  _EVAL_53__EVAL_55_data;
  wire  _EVAL_53__EVAL_55_addr;
  wire  _EVAL_53__EVAL_55_mask;
  wire  _EVAL_53__EVAL_55_en;
  wire  _EVAL_56;
  wire  _EVAL_57;
  reg [31:0] _EVAL_58 [0:1];
  reg [31:0] _RAND_10;
  wire [31:0] _EVAL_58__EVAL_59_data;
  wire  _EVAL_58__EVAL_59_addr;
  wire [31:0] _EVAL_58__EVAL_60_data;
  wire  _EVAL_58__EVAL_60_addr;
  wire  _EVAL_58__EVAL_60_mask;
  wire  _EVAL_58__EVAL_60_en;
  wire [1:0] _EVAL_61;
  assign _EVAL_21__EVAL_22_addr = _EVAL_32;
  assign _EVAL_21__EVAL_22_data = _EVAL_21[_EVAL_21__EVAL_22_addr];
  assign _EVAL_21__EVAL_23_data = _EVAL_7;
  assign _EVAL_21__EVAL_23_addr = _EVAL_29;
  assign _EVAL_21__EVAL_23_mask = 1'h1;
  assign _EVAL_21__EVAL_23_en = _EVAL_17 & _EVAL_1;
  assign _EVAL_25__EVAL_26_addr = _EVAL_32;
  assign _EVAL_25__EVAL_26_data = _EVAL_25[_EVAL_25__EVAL_26_addr];
  assign _EVAL_25__EVAL_27_data = _EVAL_13;
  assign _EVAL_25__EVAL_27_addr = _EVAL_29;
  assign _EVAL_25__EVAL_27_mask = 1'h1;
  assign _EVAL_25__EVAL_27_en = _EVAL_17 & _EVAL_1;
  assign _EVAL_37__EVAL_38_addr = _EVAL_32;
  assign _EVAL_37__EVAL_38_data = _EVAL_37[_EVAL_37__EVAL_38_addr];
  assign _EVAL_37__EVAL_39_data = _EVAL_2;
  assign _EVAL_37__EVAL_39_addr = _EVAL_29;
  assign _EVAL_37__EVAL_39_mask = 1'h1;
  assign _EVAL_37__EVAL_39_en = _EVAL_17 & _EVAL_1;
  assign _EVAL_40__EVAL_41_addr = _EVAL_32;
  assign _EVAL_40__EVAL_41_data = _EVAL_40[_EVAL_40__EVAL_41_addr];
  assign _EVAL_40__EVAL_42_data = _EVAL_0;
  assign _EVAL_40__EVAL_42_addr = _EVAL_29;
  assign _EVAL_40__EVAL_42_mask = 1'h1;
  assign _EVAL_40__EVAL_42_en = _EVAL_17 & _EVAL_1;
  assign _EVAL_43__EVAL_44_addr = _EVAL_32;
  assign _EVAL_43__EVAL_44_data = _EVAL_43[_EVAL_43__EVAL_44_addr];
  assign _EVAL_43__EVAL_45_data = _EVAL_20;
  assign _EVAL_43__EVAL_45_addr = _EVAL_29;
  assign _EVAL_43__EVAL_45_mask = 1'h1;
  assign _EVAL_43__EVAL_45_en = _EVAL_17 & _EVAL_1;
  assign _EVAL_49__EVAL_50_addr = _EVAL_32;
  assign _EVAL_49__EVAL_50_data = _EVAL_49[_EVAL_49__EVAL_50_addr];
  assign _EVAL_49__EVAL_51_data = _EVAL_10;
  assign _EVAL_49__EVAL_51_addr = _EVAL_29;
  assign _EVAL_49__EVAL_51_mask = 1'h1;
  assign _EVAL_49__EVAL_51_en = _EVAL_17 & _EVAL_1;
  assign _EVAL_53__EVAL_54_addr = _EVAL_32;
  assign _EVAL_53__EVAL_54_data = _EVAL_53[_EVAL_53__EVAL_54_addr];
  assign _EVAL_53__EVAL_55_data = _EVAL_19;
  assign _EVAL_53__EVAL_55_addr = _EVAL_29;
  assign _EVAL_53__EVAL_55_mask = 1'h1;
  assign _EVAL_53__EVAL_55_en = _EVAL_17 & _EVAL_1;
  assign _EVAL_58__EVAL_59_addr = _EVAL_32;
  assign _EVAL_58__EVAL_59_data = _EVAL_58[_EVAL_58__EVAL_59_addr];
  assign _EVAL_58__EVAL_60_data = _EVAL_9;
  assign _EVAL_58__EVAL_60_addr = _EVAL_29;
  assign _EVAL_58__EVAL_60_mask = 1'h1;
  assign _EVAL_58__EVAL_60_en = _EVAL_17 & _EVAL_1;
  assign _EVAL_24 = _EVAL_30 != _EVAL_48;
  assign _EVAL_57 = _EVAL_56 & _EVAL_34;
  assign _EVAL_17 = ~_EVAL_46;
  assign _EVAL_8 = _EVAL_49__EVAL_50_data;
  assign _EVAL_14 = _EVAL_53__EVAL_54_data;
  assign _EVAL_46 = _EVAL_56 & _EVAL_31;
  assign _EVAL_56 = _EVAL_29 == _EVAL_32;
  assign _EVAL_6 = _EVAL_25__EVAL_26_data;
  assign _EVAL_12 = _EVAL_43__EVAL_44_data;
  assign _EVAL_16 = _EVAL_40__EVAL_41_data;
  assign _EVAL_61 = _EVAL_29 + 1'h1;
  assign _EVAL_4 = ~_EVAL_57;
  assign _EVAL_48 = _EVAL_5 & _EVAL_4;
  assign _EVAL_30 = _EVAL_17 & _EVAL_1;
  assign _EVAL_47 = _EVAL_32 + 1'h1;
  assign _EVAL_34 = ~_EVAL_31;
  assign _EVAL_11 = _EVAL_58__EVAL_59_data;
  assign _EVAL_35 = _EVAL_47[0];
  assign _EVAL_52 = _EVAL_61[0];
  assign _EVAL_15 = _EVAL_37__EVAL_38_data;
  assign _EVAL = _EVAL_21__EVAL_22_data;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_21[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_25[initvar] = _RAND_1[3:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_29 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_31 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_32 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_37[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_40[initvar] = _RAND_6[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_43[initvar] = _RAND_7[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_49[initvar] = _RAND_8[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_53[initvar] = _RAND_9[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_58[initvar] = _RAND_10[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_18) begin
    if(_EVAL_21__EVAL_23_en & _EVAL_21__EVAL_23_mask) begin
      _EVAL_21[_EVAL_21__EVAL_23_addr] <= _EVAL_21__EVAL_23_data;
    end
    if(_EVAL_25__EVAL_27_en & _EVAL_25__EVAL_27_mask) begin
      _EVAL_25[_EVAL_25__EVAL_27_addr] <= _EVAL_25__EVAL_27_data;
    end
    if (_EVAL_3) begin
      _EVAL_29 <= 1'h0;
    end else if (_EVAL_30) begin
      _EVAL_29 <= _EVAL_52;
    end
    if (_EVAL_3) begin
      _EVAL_31 <= 1'h0;
    end else if (_EVAL_24) begin
      _EVAL_31 <= _EVAL_30;
    end
    if (_EVAL_3) begin
      _EVAL_32 <= 1'h0;
    end else if (_EVAL_48) begin
      _EVAL_32 <= _EVAL_35;
    end
    if(_EVAL_37__EVAL_39_en & _EVAL_37__EVAL_39_mask) begin
      _EVAL_37[_EVAL_37__EVAL_39_addr] <= _EVAL_37__EVAL_39_data;
    end
    if(_EVAL_40__EVAL_42_en & _EVAL_40__EVAL_42_mask) begin
      _EVAL_40[_EVAL_40__EVAL_42_addr] <= _EVAL_40__EVAL_42_data;
    end
    if(_EVAL_43__EVAL_45_en & _EVAL_43__EVAL_45_mask) begin
      _EVAL_43[_EVAL_43__EVAL_45_addr] <= _EVAL_43__EVAL_45_data;
    end
    if(_EVAL_49__EVAL_51_en & _EVAL_49__EVAL_51_mask) begin
      _EVAL_49[_EVAL_49__EVAL_51_addr] <= _EVAL_49__EVAL_51_data;
    end
    if(_EVAL_53__EVAL_55_en & _EVAL_53__EVAL_55_mask) begin
      _EVAL_53[_EVAL_53__EVAL_55_addr] <= _EVAL_53__EVAL_55_data;
    end
    if(_EVAL_58__EVAL_60_en & _EVAL_58__EVAL_60_mask) begin
      _EVAL_58[_EVAL_58__EVAL_60_addr] <= _EVAL_58__EVAL_60_data;
    end
  end
endmodule
