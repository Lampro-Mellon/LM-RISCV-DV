//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_67_assert(
  input         _EVAL_1,
  input  [2:0]  _EVAL_5,
  input         _EVAL_12,
  input         _EVAL_16,
  input  [2:0]  _EVAL_17,
  input  [3:0]  _EVAL_23,
  input         _EVAL_32,
  input  [29:0] _EVAL_36,
  input  [3:0]  _EVAL_37,
  input  [2:0]  _EVAL_41,
  input         _EVAL_43,
  input         Queue_1__EVAL_4,
  input  [2:0]  Queue_1__EVAL_16,
  input  [3:0]  Queue_1__EVAL_6,
  input  [1:0]  Queue_1__EVAL_8,
  input         Queue_1__EVAL_15,
  input         Queue__EVAL_11,
  input         Queue_1__EVAL,
  input         Queue_1__EVAL_14,
  input  [2:0]  Queue_1__EVAL_12
);
  wire [2:0] TLMonitor__EVAL;
  wire [2:0] TLMonitor__EVAL_0;
  wire [3:0] TLMonitor__EVAL_1;
  wire [2:0] TLMonitor__EVAL_2;
  wire [3:0] TLMonitor__EVAL_3;
  wire  TLMonitor__EVAL_4;
  wire  TLMonitor__EVAL_5;
  wire [1:0] TLMonitor__EVAL_6;
  wire  TLMonitor__EVAL_7;
  wire  TLMonitor__EVAL_8;
  wire  TLMonitor__EVAL_9;
  wire  TLMonitor__EVAL_10;
  wire  TLMonitor__EVAL_11;
  wire  TLMonitor__EVAL_12;
  wire [2:0] TLMonitor__EVAL_13;
  wire  TLMonitor__EVAL_14;
  wire  TLMonitor__EVAL_15;
  wire [2:0] TLMonitor__EVAL_16;
  wire [29:0] TLMonitor__EVAL_17;
  wire [3:0] TLMonitor__EVAL_18;
  _EVAL_64_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14),
    ._EVAL_15(TLMonitor__EVAL_15),
    ._EVAL_16(TLMonitor__EVAL_16),
    ._EVAL_17(TLMonitor__EVAL_17),
    ._EVAL_18(TLMonitor__EVAL_18)
  );
  assign TLMonitor__EVAL_5 = Queue_1__EVAL_4;
  assign TLMonitor__EVAL_2 = _EVAL_17;
  assign TLMonitor__EVAL_1 = _EVAL_37;
  assign TLMonitor__EVAL_13 = Queue_1__EVAL_16;
  assign TLMonitor__EVAL_18 = Queue_1__EVAL_6;
  assign TLMonitor__EVAL_6 = Queue_1__EVAL_8;
  assign TLMonitor__EVAL = _EVAL_5;
  assign TLMonitor__EVAL_17 = _EVAL_36;
  assign TLMonitor__EVAL_10 = Queue_1__EVAL_15;
  assign TLMonitor__EVAL_9 = _EVAL_12;
  assign TLMonitor__EVAL_7 = Queue__EVAL_11;
  assign TLMonitor__EVAL_4 = Queue_1__EVAL;
  assign TLMonitor__EVAL_12 = Queue_1__EVAL_14;
  assign TLMonitor__EVAL_3 = _EVAL_23;
  assign TLMonitor__EVAL_15 = _EVAL_43;
  assign TLMonitor__EVAL_0 = Queue_1__EVAL_12;
  assign TLMonitor__EVAL_14 = _EVAL_16;
  assign TLMonitor__EVAL_8 = _EVAL_32;
  assign TLMonitor__EVAL_16 = _EVAL_41;
  assign TLMonitor__EVAL_11 = _EVAL_1;

endmodule
