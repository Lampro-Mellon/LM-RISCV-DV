//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_141(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  output [1:0]  _EVAL_1,
  input         _EVAL_2,
  input  [9:0]  _EVAL_3,
  output [2:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  output        _EVAL_6,
  input         _EVAL_7,
  output        _EVAL_8,
  output [31:0] _EVAL_9,
  output [31:0] _EVAL_10,
  input  [31:0] _EVAL_11,
  input         _EVAL_12,
  input  [2:0]  _EVAL_13,
  input  [1:0]  _EVAL_14,
  input  [2:0]  _EVAL_15,
  output        _EVAL_16,
  output        _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  input         _EVAL_20,
  input  [8:0]  _EVAL_21,
  input         _EVAL_22,
  output [1:0]  _EVAL_23,
  output [2:0]  _EVAL_24,
  input         _EVAL_25,
  input  [31:0] _EVAL_26,
  output        _EVAL_27,
  input  [3:0]  _EVAL_28,
  input  [3:0]  _EVAL_29,
  input         _EVAL_30,
  output [2:0]  _EVAL_31,
  input         _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_34,
  output        _EVAL_35,
  input  [11:0] _EVAL_36,
  output        _EVAL_37,
  input         _EVAL_38,
  input  [2:0]  _EVAL_39,
  input  [1:0]  _EVAL_40,
  input         _EVAL_41
);
  wire  _EVAL_45;
  wire [31:0] _EVAL_49;
  wire [31:0] _EVAL_51;
  wire [31:0] _EVAL_54;
  wire [31:0] _EVAL_55;
  wire  _EVAL_56;
  wire [31:0] _EVAL_58;
  wire [15:0] _EVAL_61;
  wire [31:0] _EVAL_63;
  wire  _EVAL_65;
  wire [31:0] _EVAL_66;
  reg [7:0] _EVAL_67;
  reg [31:0] _RAND_0;
  wire  _EVAL_71;
  wire [31:0] _EVAL_72;
  wire  _EVAL_76;
  wire [31:0] _EVAL_78;
  wire  _EVAL_79;
  wire [31:0] _EVAL_83;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_90;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire [7:0] _EVAL_95;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire [31:0] _EVAL_102;
  wire [31:0] _EVAL_109;
  wire [31:0] _EVAL_110;
  wire [31:0] _EVAL_111;
  wire  _EVAL_113;
  wire  _EVAL_115;
  wire  _EVAL_117;
  wire [31:0] _EVAL_118;
  wire  _EVAL_121;
  wire [31:0] _EVAL_123;
  wire  _EVAL_124;
  wire [31:0] _EVAL_125;
  wire  _EVAL_126;
  wire [31:0] _EVAL_127;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire [31:0] _EVAL_133;
  wire  _EVAL_139;
  wire [31:0] _EVAL_143;
  wire [22:0] _EVAL_147;
  wire  _EVAL_150;
  wire [31:0] _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_156;
  reg [15:0] _EVAL_167;
  reg [31:0] _RAND_1;
  wire  _EVAL_169;
  wire  _EVAL_171;
  wire [31:0] _EVAL_172;
  wire  _EVAL_174;
  wire [31:0] _EVAL_175;
  wire  _EVAL_178;
  wire [31:0] _EVAL_179;
  wire  _EVAL_180;
  wire [2:0] _EVAL_181;
  wire [31:0] _EVAL_182;
  wire [31:0] _EVAL_184;
  wire  _EVAL_187;
  wire [31:0] _EVAL_191;
  wire [31:0] _EVAL_198;
  wire  _EVAL_200;
  wire  _EVAL_202;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire [31:0] _EVAL_207;
  wire  _EVAL_209;
  wire [31:0] _EVAL_212;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_217;
  wire  _EVAL_219;
  wire [31:0] _EVAL_223;
  wire  _EVAL_225;
  wire [31:0] _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_236;
  wire [31:0] _EVAL_238;
  wire [31:0] _EVAL_239;
  wire  _EVAL_244;
  wire  _EVAL_248;
  wire [31:0] _EVAL_249;
  wire [31:0] _EVAL_251;
  wire [31:0] _EVAL_256;
  wire [31:0] _EVAL_257;
  wire [31:0] _EVAL_258;
  wire [31:0] _EVAL_259;
  wire  _EVAL_265;
  reg [7:0] _EVAL_266;
  reg [31:0] _RAND_2;
  wire [31:0] _EVAL_268;
  wire [31:0] _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_275;
  wire  _EVAL_279;
  wire [16:0] _EVAL_280;
  wire [23:0] _EVAL_282;
  wire  _EVAL_285;
  wire  _EVAL_304;
  wire [9:0] _EVAL_306;
  wire [31:0] _EVAL_308;
  wire [31:0] _EVAL_311;
  wire [31:0] _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_317;
  wire  _EVAL_320;
  wire  _EVAL_323;
  wire [31:0] _EVAL_324;
  wire [31:0] _EVAL_325;
  wire [31:0] _EVAL_327;
  wire  _EVAL_329;
  wire  _EVAL_331;
  wire [31:0] _EVAL_332;
  wire  _EVAL_333;
  wire  _EVAL_334;
  wire  _EVAL_339;
  wire  _EVAL_343;
  wire [31:0] _EVAL_344;
  wire  _EVAL_347;
  reg [7:0] _EVAL_351;
  reg [31:0] _RAND_3;
  wire [31:0] _EVAL_353;
  wire [31:0] _EVAL_354;
  wire  _EVAL_360;
  wire  _EVAL_363;
  wire  _EVAL_365;
  wire  _EVAL_366;
  wire  _EVAL_368;
  wire  _EVAL_370;
  wire  _EVAL_372;
  wire [31:0] _EVAL_374;
  wire  _EVAL_375;
  wire [31:0] _EVAL_377;
  wire  _EVAL_378;
  wire  _EVAL_382;
  wire  _EVAL_384;
  wire  _EVAL_386;
  wire  _EVAL_389;
  wire  _EVAL_392;
  wire [31:0] _EVAL_393;
  wire  _EVAL_397;
  wire  _EVAL_401;
  wire  _EVAL_402;
  wire  _EVAL_403;
  wire  _EVAL_406;
  wire  _EVAL_407;
  wire [31:0] _EVAL_409;
  wire  _EVAL_412;
  wire  _EVAL_415;
  wire [31:0] _EVAL_417;
  wire [31:0] _EVAL_419;
  wire  _EVAL_420;
  wire  _EVAL_421;
  wire  _EVAL_431;
  wire [31:0] _EVAL_432;
  wire [31:0] _EVAL_434;
  wire [31:0] _EVAL_436;
  wire  _EVAL_439;
  wire [31:0] _EVAL_442;
  wire  _EVAL_448;
  wire [31:0] _EVAL_450;
  wire  _EVAL_451;
  wire  _EVAL_458;
  wire  _EVAL_459;
  wire  _EVAL_463;
  wire  _EVAL_464;
  wire  _EVAL_468;
  wire  _EVAL_470;
  wire [31:0] _EVAL_471;
  wire  _EVAL_473;
  wire  _EVAL_474;
  wire  _EVAL_477;
  wire  _EVAL_479;
  wire  _EVAL_480;
  wire  _EVAL_481;
  wire  _EVAL_484;
  wire [31:0] _EVAL_485;
  wire [31:0] _EVAL_486;
  wire  _EVAL_487;
  wire  _EVAL_488;
  wire [31:0] _EVAL_492;
  wire  _EVAL_493;
  wire  _EVAL_497;
  wire  _EVAL_498;
  wire  _EVAL_499;
  wire  _EVAL_502;
  wire  _EVAL_505;
  wire  _EVAL_506;
  wire  _EVAL_509;
  wire  _EVAL_510;
  wire  _EVAL_512;
  wire  _EVAL_514;
  wire  _EVAL_516;
  wire  _EVAL_519;
  wire  _EVAL_526;
  wire [31:0] _EVAL_527;
  wire [7:0] _EVAL_530;
  wire [31:0] _EVAL_533;
  wire [31:0] _EVAL_538;
  wire [31:0] _EVAL_540;
  wire [31:0] _EVAL_541;
  wire  _EVAL_542;
  wire  _EVAL_545;
  wire [31:0] _EVAL_546;
  wire [31:0] _EVAL_547;
  wire  _EVAL_549;
  wire [7:0] _EVAL_551;
  wire [31:0] _EVAL_552;
  wire  _EVAL_554;
  reg [7:0] _EVAL_555;
  reg [31:0] _RAND_4;
  wire  _EVAL_558;
  wire [31:0] _EVAL_559;
  wire  _EVAL_563;
  wire  _EVAL_565;
  wire [31:0] _EVAL_566;
  wire [31:0] _EVAL_567;
  wire  _EVAL_569;
  wire  _EVAL_571;
  wire  _EVAL_572;
  wire [31:0] _EVAL_575;
  wire  _EVAL_577;
  wire  _EVAL_583;
  wire  _EVAL_585;
  wire [31:0] _EVAL_592;
  wire  _EVAL_599;
  wire [31:0] _EVAL_601;
  wire  _EVAL_602;
  wire [31:0] _EVAL_605;
  wire  _EVAL_606;
  wire  _EVAL_607;
  wire [31:0] _EVAL_608;
  wire [31:0] _EVAL_611;
  wire [1:0] _EVAL_612;
  wire [31:0] _EVAL_613;
  wire [31:0] _EVAL_614;
  wire  _EVAL_616;
  wire  _EVAL_617;
  wire  _EVAL_619;
  wire  _EVAL_620;
  wire  _EVAL_622;
  wire  _EVAL_624;
  wire  _EVAL_628;
  wire [31:0] _EVAL_630;
  wire [31:0] _EVAL_634;
  wire  _EVAL_636;
  wire  _EVAL_638;
  wire  _EVAL_642;
  wire  _EVAL_645;
  wire  _EVAL_649;
  wire  _EVAL_650;
  wire  _EVAL_651;
  wire [31:0] _EVAL_653;
  wire  _EVAL_654;
  wire  _EVAL_659;
  wire [31:0] _EVAL_662;
  wire [31:0] _EVAL_669;
  wire  _EVAL_674;
  wire  _EVAL_679;
  wire  _EVAL_683;
  wire  _EVAL_685;
  wire [31:0] _EVAL_686;
  wire  _EVAL_689;
  wire [31:0] _EVAL_692;
  wire  _EVAL_696;
  wire  _EVAL_697;
  wire  _EVAL_699;
  wire  _EVAL_700;
  wire [31:0] _EVAL_702;
  wire  _EVAL_705;
  wire [31:0] _EVAL_707;
  wire  _EVAL_710;
  wire  _EVAL_711;
  wire  _EVAL_713;
  wire  _EVAL_719;
  wire  _EVAL_721;
  wire [31:0] _EVAL_722;
  wire [31:0] _EVAL_723;
  wire  _EVAL_724;
  wire  _EVAL_725;
  wire [31:0] _EVAL_727;
  wire  _EVAL_728;
  wire  _EVAL_730;
  wire  _EVAL_734;
  wire [31:0] _EVAL_735;
  wire  _EVAL_736;
  wire  _EVAL_739;
  wire  _EVAL_744;
  wire  _EVAL_748;
  wire [31:0] _EVAL_751;
  wire  _EVAL_752;
  wire  _EVAL_753;
  wire  _EVAL_754;
  wire  _EVAL_757;
  wire  _EVAL_759;
  wire  _EVAL_760;
  wire  _EVAL_762;
  wire  _EVAL_763;
  wire [31:0] _EVAL_765;
  wire [31:0] _EVAL_766;
  wire  _EVAL_768;
  wire  _EVAL_769;
  wire  _EVAL_771;
  wire  _EVAL_774;
  wire  _EVAL_784;
  wire  _EVAL_785;
  wire  _EVAL_788;
  wire [31:0] _EVAL_789;
  wire [31:0] _EVAL_790;
  wire  _EVAL_792;
  wire  _EVAL_793;
  wire  _EVAL_795;
  wire  _EVAL_797;
  wire [31:0] _EVAL_799;
  wire  _EVAL_802;
  wire  _EVAL_808;
  wire [31:0] _EVAL_809;
  wire [31:0] _EVAL_815;
  wire  _EVAL_817;
  reg [23:0] _EVAL_819;
  reg [31:0] _RAND_5;
  wire [31:0] _EVAL_820;
  wire  _EVAL_822;
  wire  _EVAL_829;
  wire  _EVAL_832;
  wire  _EVAL_833;
  wire [31:0] _EVAL_835;
  wire  _EVAL_836;
  wire [31:0] _EVAL_837;
  wire [31:0] _EVAL_841;
  wire  _EVAL_842;
  wire  _EVAL_846;
  wire  _EVAL_847;
  wire [31:0] _EVAL_849;
  wire  _EVAL_851;
  wire  _EVAL_857;
  wire [31:0] _EVAL_858;
  wire [23:0] _EVAL_859;
  wire  _EVAL_861;
  wire  _EVAL_863;
  wire  _EVAL_866;
  wire  _EVAL_867;
  wire  _EVAL_868;
  wire [31:0] _EVAL_869;
  wire [9:0] _EVAL_870;
  wire  _EVAL_876;
  wire  _EVAL_879;
  wire  _EVAL_881;
  wire [31:0] _EVAL_882;
  wire  _EVAL_886;
  wire  _EVAL_890;
  wire [31:0] _EVAL_891;
  wire  _EVAL_895;
  wire  _EVAL_900;
  wire  _EVAL_906;
  wire [31:0] _EVAL_908;
  wire [31:0] _EVAL_909;
  wire [31:0] _EVAL_910;
  wire [31:0] _EVAL_912;
  wire  _EVAL_916;
  wire  _EVAL_921;
  wire [31:0] _EVAL_922;
  wire  _EVAL_926;
  wire [31:0] _EVAL_930;
  wire [31:0] _EVAL_931;
  wire  _EVAL_934;
  wire  _EVAL_941;
  wire [31:0] _EVAL_942;
  wire [31:0] _EVAL_943;
  wire [31:0] _EVAL_946;
  wire [31:0] _EVAL_949;
  wire  _EVAL_951;
  wire  _EVAL_952;
  wire [31:0] _EVAL_956;
  wire [4:0] _EVAL_957;
  wire [4:0] _EVAL_958;
  wire  _EVAL_959;
  wire [31:0] _EVAL_960;
  wire [31:0] _EVAL_963;
  wire [31:0] _EVAL_964;
  wire  _EVAL_965;
  wire [31:0] _EVAL_967;
  wire  _EVAL_968;
  wire  _EVAL_969;
  wire [31:0] _EVAL_972;
  wire  _EVAL_982;
  wire  _EVAL_984;
  wire  _EVAL_985;
  wire  _EVAL_987;
  wire [31:0] _EVAL_990;
  wire [7:0] _EVAL_991;
  wire [31:0] _EVAL_993;
  wire [31:0] _EVAL_995;
  wire  _EVAL_996;
  wire  _EVAL_997;
  wire [31:0] _EVAL_1000;
  wire [31:0] _EVAL_1003;
  wire [31:0] _EVAL_1004;
  wire [31:0] _EVAL_1007;
  wire  _EVAL_1008;
  wire  _EVAL_1010;
  wire [31:0] _EVAL_1012;
  wire  _EVAL_1014;
  wire [31:0] _EVAL_1015;
  wire  _EVAL_1018;
  wire [31:0] _EVAL_1019;
  wire  _EVAL_1020;
  wire  _EVAL_1021;
  wire  _EVAL_1023;
  wire [31:0] _EVAL_1026;
  wire [31:0] _EVAL_1030;
  wire  _EVAL_1031;
  wire  _EVAL_1034;
  wire  _EVAL_1035;
  wire [31:0] _EVAL_1036;
  wire  _EVAL_1037;
  wire  _EVAL_1038;
  wire  _EVAL_1039;
  wire  _EVAL_1040;
  wire [31:0] _EVAL_1041;
  wire  _EVAL_1044;
  wire  _EVAL_1045;
  wire  _EVAL_1046;
  wire  _EVAL_1047;
  wire  _EVAL_1049;
  wire  _EVAL_1050;
  wire  _EVAL_1051;
  wire  _EVAL_1052;
  wire  _EVAL_1057;
  wire  _EVAL_1066;
  wire  _EVAL_1069;
  wire  _EVAL_1071;
  wire [31:0] _EVAL_1073;
  wire  _EVAL_1077;
  wire  _EVAL_1081;
  wire  _EVAL_1082;
  wire [31:0] _EVAL_1084;
  wire [31:0] _EVAL_1087;
  wire  _EVAL_1089;
  wire  _EVAL_1095;
  wire [31:0] _EVAL_1096;
  wire  _EVAL_1097;
  wire  _EVAL_1098;
  wire  _EVAL_1099;
  wire  _EVAL_1101;
  wire [31:0] _EVAL_1104;
  wire [31:0] _EVAL_1109;
  wire  _EVAL_1110;
  wire  _EVAL_1114;
  wire  _EVAL_1115;
  wire  _EVAL_1116;
  wire  _EVAL_1121;
  wire  _EVAL_1123;
  wire  _EVAL_1124;
  wire [31:0] _EVAL_1125;
  wire  _EVAL_1127;
  wire  _EVAL_1132;
  wire [31:0] _EVAL_1133;
  wire  _EVAL_1135;
  wire  _EVAL_1136;
  wire  _EVAL_1138;
  wire [31:0] _EVAL_1139;
  wire [31:0] _EVAL_1140;
  wire  _EVAL_1145;
  wire [31:0] _EVAL_1147;
  wire  _EVAL_1149;
  wire [31:0] _EVAL_1150;
  wire  _EVAL_1151;
  wire  _EVAL_1152;
  wire [31:0] _EVAL_1154;
  wire  _EVAL_1155;
  wire  _EVAL_1159;
  wire  _EVAL_1160;
  wire  _EVAL_1163;
  wire  _EVAL_1166;
  wire [31:0] _EVAL_1167;
  wire [31:0] _EVAL_1170;
  wire  _EVAL_1174;
  wire  _EVAL_1175;
  wire  _EVAL_1176;
  wire  _EVAL_1177;
  wire  _EVAL_1181;
  wire  _EVAL_1182;
  wire  _EVAL_1183;
  wire  _EVAL_1184;
  wire  _EVAL_1185;
  wire  _EVAL_1186;
  wire  _EVAL_1191;
  wire  _EVAL_1194;
  wire [31:0] _EVAL_1196;
  wire  _EVAL_1198;
  wire [31:0] _EVAL_1200;
  wire  _EVAL_1206;
  wire  _EVAL_1211;
  wire [31:0] _EVAL_1213;
  wire  _EVAL_1215;
  wire  _EVAL_1217;
  wire [17:0] _EVAL_1218;
  wire [31:0] _EVAL_1219;
  wire  _EVAL_1220;
  wire [31:0] _EVAL_1221;
  wire  _EVAL_1224;
  wire  _EVAL_1226;
  wire  _EVAL_1228;
  wire  _EVAL_1230;
  wire  _EVAL_1231;
  wire  _EVAL_1237;
  wire  _EVAL_1238;
  wire  _EVAL_1240;
  wire [31:0] _EVAL_1243;
  wire [31:0] _EVAL_1244;
  wire  _EVAL_1251;
  wire [31:0] _EVAL_1257;
  wire  _EVAL_1258;
  wire  _EVAL_1261;
  wire  _EVAL_1268;
  wire [31:0] _EVAL_1269;
  wire [31:0] _EVAL_1270;
  wire  _EVAL_1271;
  wire  _EVAL_1273;
  wire  _EVAL_1274;
  wire  _EVAL_1275;
  wire [31:0] _EVAL_1276;
  wire [31:0] _EVAL_1285;
  wire [31:0] _EVAL_1290;
  wire [31:0] _EVAL_1297;
  wire  _EVAL_1303;
  wire  _EVAL_1304;
  wire  _EVAL_1307;
  wire  _EVAL_1311;
  wire [31:0] _EVAL_1312;
  wire  _EVAL_1314;
  wire [7:0] _EVAL_1319;
  wire  _EVAL_1321;
  wire [31:0] _EVAL_1324;
  wire [31:0] _EVAL_1325;
  wire  _EVAL_1326;
  wire [31:0] _EVAL_1328;
  wire [31:0] _EVAL_1331;
  wire  _EVAL_1332;
  wire  _EVAL_1334;
  wire  _EVAL_1335;
  wire  _EVAL_1337;
  wire [11:0] _EVAL_1339;
  wire  _EVAL_1341;
  wire [31:0] _EVAL_1343;
  wire  _EVAL_1347;
  wire  _EVAL_1348;
  wire [31:0] _EVAL_1350;
  wire [31:0] _EVAL_1351;
  wire  _EVAL_1357;
  wire  _EVAL_1358;
  wire  _EVAL_1360;
  wire  _EVAL_1362;
  wire [31:0] _EVAL_1365;
  wire [31:0] _EVAL_1366;
  wire  _EVAL_1367;
  wire  _EVAL_1368;
  wire [31:0] _EVAL_1370;
  wire  _EVAL_1374;
  wire  _EVAL_1375;
  wire  _EVAL_1376;
  wire [31:0] _EVAL_1377;
  wire  _EVAL_1380;
  wire [31:0] _EVAL_1383;
  wire  _EVAL_1390;
  wire [31:0] _EVAL_1392;
  wire [31:0] _EVAL_1395;
  wire [8:0] _EVAL_1399;
  wire  _EVAL_1400;
  wire [31:0] _EVAL_1401;
  wire  _EVAL_1407;
  wire  _EVAL_1408;
  wire [31:0] _EVAL_1410;
  wire [31:0] _EVAL_1419;
  wire  _EVAL_1420;
  wire  _EVAL_1422;
  wire  _EVAL_1423;
  wire  _EVAL_1425;
  wire  _EVAL_1426;
  wire  _EVAL_1429;
  wire  _EVAL_1433;
  wire [31:0] _EVAL_1435;
  wire [31:0] _EVAL_1436;
  wire  _EVAL_1437;
  wire  _EVAL_1441;
  wire  _EVAL_1445;
  wire  _EVAL_1448;
  wire  _EVAL_1450;
  wire  _EVAL_1460;
  wire  _EVAL_1461;
  wire [31:0] _EVAL_1462;
  wire [31:0] _EVAL_1465;
  wire  _EVAL_1467;
  wire [31:0] _EVAL_1469;
  wire [31:0] _EVAL_1470;
  wire  _EVAL_1471;
  wire  _EVAL_1472;
  wire  _EVAL_1475;
  wire  _EVAL_1476;
  wire [31:0] _EVAL_1477;
  wire [31:0] _EVAL_1478;
  wire  _EVAL_1480;
  wire  _EVAL_1486;
  wire  _EVAL_1487;
  wire [31:0] _EVAL_1490;
  wire  _EVAL_1493;
  wire  _EVAL_1494;
  wire [31:0] _EVAL_1495;
  wire  _EVAL_1496;
  wire  _EVAL_1506;
  wire  _EVAL_1507;
  wire  _EVAL_1508;
  wire  _EVAL_1512;
  wire [31:0] _EVAL_1513;
  wire [31:0] _EVAL_1514;
  wire [31:0] _EVAL_1516;
  wire  _EVAL_1517;
  wire  _EVAL_1518;
  wire  _EVAL_1523;
  wire [31:0] _EVAL_1525;
  wire [31:0] _EVAL_1527;
  wire  _EVAL_1528;
  wire [31:0] _EVAL_1530;
  wire [31:0] _EVAL_1532;
  wire  _EVAL_1538;
  wire  _EVAL_1540;
  wire  _EVAL_1541;
  wire  _EVAL_1544;
  wire [31:0] _EVAL_1545;
  wire [31:0] _EVAL_1547;
  wire  _EVAL_1549;
  wire [7:0] _EVAL_1552;
  wire  _EVAL_1553;
  wire [31:0] _EVAL_1556;
  wire  _EVAL_1557;
  wire  _EVAL_1561;
  wire  _EVAL_1562;
  wire  _EVAL_1564;
  wire  _EVAL_1567;
  wire  _EVAL_1568;
  wire  _EVAL_1569;
  wire [31:0] _EVAL_1571;
  wire  _EVAL_1572;
  wire  _EVAL_1575;
  wire [31:0] _EVAL_1576;
  wire [31:0] _EVAL_1578;
  wire [31:0] _EVAL_1583;
  wire [31:0] _EVAL_1587;
  wire  _EVAL_1589;
  wire  _EVAL_1590;
  wire [31:0] _EVAL_1591;
  wire [21:0] _EVAL_1592;
  wire [31:0] _EVAL_1593;
  wire  _EVAL_1594;
  wire  _EVAL_1597;
  wire [31:0] _EVAL_1598;
  wire  _EVAL_1599;
  wire  _EVAL_1603;
  wire  _EVAL_1606;
  wire  _EVAL_1611;
  wire [31:0] _EVAL_1613;
  wire [31:0] _EVAL_1615;
  wire  _EVAL_1620;
  wire [31:0] _EVAL_1622;
  wire  _EVAL_1631;
  wire [31:0] _EVAL_1633;
  wire [31:0] _EVAL_1639;
  wire [31:0] _EVAL_1641;
  wire  _EVAL_1646;
  wire  _EVAL_1650;
  wire [31:0] _EVAL_1653;
  wire  _EVAL_1654;
  wire [31:0] _EVAL_1658;
  wire  _EVAL_1659;
  wire  _EVAL_1665;
  wire  _EVAL_1666;
  wire  _EVAL_1669;
  wire [31:0] _EVAL_1672;
  wire  _EVAL_1675;
  wire [31:0] _EVAL_1677;
  wire  _EVAL_1681;
  wire [9:0] _EVAL_1682;
  wire  _EVAL_1684;
  wire [31:0] _EVAL_1685;
  wire  _EVAL_1687;
  wire  _EVAL_1693;
  wire [31:0] _EVAL_1697;
  wire  _EVAL_1699;
  wire  _EVAL_1701;
  wire  _EVAL_1706;
  wire [31:0] _EVAL_1710;
  wire  _EVAL_1713;
  wire [31:0] _EVAL_1718;
  wire  _EVAL_1720;
  wire  _EVAL_1721;
  wire  debug_hartReset_0__EVAL;
  wire  debug_hartReset_0__EVAL_0;
  wire  debug_hartReset_0__EVAL_1;
  wire  debug_hartReset_0__EVAL_2;
  wire [31:0] _EVAL_1723;
  wire [31:0] _EVAL_1724;
  wire [31:0] _EVAL_1725;
  wire  _EVAL_1728;
  wire [31:0] _EVAL_1731;
  wire [31:0] _EVAL_1732;
  wire  _EVAL_1734;
  wire [31:0] _EVAL_1736;
  wire [31:0] _EVAL_1738;
  wire  _EVAL_1742;
  wire  _EVAL_1746;
  wire  _EVAL_1747;
  wire  _EVAL_1752;
  wire  _EVAL_1754;
  wire [31:0] _EVAL_1755;
  wire  _EVAL_1758;
  wire  _EVAL_1759;
  wire  _EVAL_1761;
  wire  _EVAL_1767;
  wire  _EVAL_1769;
  wire  _EVAL_1771;
  wire  _EVAL_1773;
  wire [31:0] _EVAL_1774;
  reg [11:0] _EVAL_1778;
  reg [31:0] _RAND_6;
  wire [31:0] _EVAL_1779;
  wire [31:0] _EVAL_1787;
  wire  _EVAL_1789;
  wire  _EVAL_1790;
  wire [31:0] _EVAL_1795;
  wire  _EVAL_1798;
  wire [31:0] _EVAL_1799;
  wire  _EVAL_1803;
  wire  _EVAL_1804;
  reg [7:0] _EVAL_1805;
  reg [31:0] _RAND_7;
  wire [31:0] _EVAL_1806;
  wire [31:0] _EVAL_1807;
  wire  _EVAL_1812;
  wire [31:0] _EVAL_1813;
  wire  _EVAL_1815;
  wire  _EVAL_1821;
  wire  _EVAL_1822;
  wire [31:0] _EVAL_1823;
  wire  _EVAL_1824;
  wire  _EVAL_1830;
  wire [31:0] _EVAL_1832;
  wire  _EVAL_1833;
  wire  _EVAL_1834;
  wire  _EVAL_1835;
  wire  _EVAL_1838;
  wire  _EVAL_1839;
  wire  _EVAL_1841;
  wire [31:0] _EVAL_1842;
  wire [31:0] _EVAL_1844;
  wire  _EVAL_1846;
  wire [31:0] _EVAL_1849;
  wire [31:0] _EVAL_1853;
  wire  _EVAL_1856;
  wire  _EVAL_1859;
  wire  _EVAL_1860;
  wire  _EVAL_1863;
  wire  _EVAL_1867;
  wire  _EVAL_1869;
  wire  _EVAL_1871;
  wire  _EVAL_1872;
  wire  _EVAL_1873;
  wire [31:0] _EVAL_1875;
  wire  _EVAL_1880;
  wire  _EVAL_1881;
  wire  _EVAL_1883;
  wire  _EVAL_1884;
  wire  _EVAL_1887;
  wire  _EVAL_1888;
  wire  _EVAL_1891;
  wire  _EVAL_1893;
  reg [7:0] _EVAL_1894;
  reg [31:0] _RAND_8;
  wire  _EVAL_1896;
  wire  _EVAL_1897;
  wire [31:0] _EVAL_1900;
  wire [31:0] _EVAL_1902;
  wire [13:0] _EVAL_1905;
  wire  _EVAL_1911;
  wire  _EVAL_1913;
  wire  _EVAL_1914;
  wire  _EVAL_1921;
  wire [31:0] _EVAL_1925;
  wire  _EVAL_1928;
  wire  _EVAL_1931;
  wire [31:0] _EVAL_1933;
  wire [31:0] _EVAL_1934;
  wire  _EVAL_1935;
  wire  _EVAL_1936;
  wire [31:0] _EVAL_1937;
  wire  _EVAL_1939;
  wire [31:0] _EVAL_1941;
  wire [31:0] _EVAL_1942;
  wire  _EVAL_1944;
  wire  _EVAL_1945;
  wire  _EVAL_1953;
  wire  _EVAL_1957;
  wire [31:0] _EVAL_1958;
  wire  _EVAL_1965;
  wire [31:0] _EVAL_1968;
  wire  _EVAL_1972;
  wire  _EVAL_1975;
  wire [31:0] _EVAL_1977;
  wire [15:0] _EVAL_1978;
  wire  _EVAL_1979;
  wire [31:0] _EVAL_1982;
  wire  _EVAL_1983;
  wire [31:0] _EVAL_1985;
  reg [1:0] _EVAL_1987;
  reg [31:0] _RAND_9;
  wire  _EVAL_1989;
  wire  _EVAL_1991;
  wire [31:0] _EVAL_1992;
  wire  _EVAL_1993;
  wire [31:0] _EVAL_1994;
  wire [31:0] _EVAL_2001;
  wire [31:0] _EVAL_2002;
  wire  _EVAL_2004;
  wire  _EVAL_2005;
  wire [31:0] _EVAL_2006;
  wire  _EVAL_2008;
  reg [2:0] _EVAL_2012;
  reg [31:0] _RAND_10;
  wire  _EVAL_2014;
  wire [31:0] _EVAL_2015;
  wire  _EVAL_2017;
  wire  _EVAL_2018;
  wire  _EVAL_2021;
  wire [31:0] _EVAL_2024;
  wire  _EVAL_2029;
  wire [31:0] _EVAL_2031;
  wire  _EVAL_2039;
  wire  _EVAL_2040;
  wire  _EVAL_2041;
  wire  _EVAL_2050;
  wire  _EVAL_2051;
  wire [31:0] _EVAL_2052;
  wire  _EVAL_2054;
  wire  _EVAL_2056;
  wire [31:0] _EVAL_2057;
  wire  _EVAL_2061;
  wire [31:0] _EVAL_2063;
  wire [31:0] _EVAL_2066;
  wire  _EVAL_2073;
  wire  _EVAL_2074;
  wire  _EVAL_2075;
  wire  _EVAL_2076;
  wire  _EVAL_2077;
  wire [31:0] _EVAL_2078;
  wire  _EVAL_2079;
  wire  _EVAL_2080;
  wire  _EVAL_2081;
  wire  _EVAL_2083;
  wire [31:0] _EVAL_2086;
  wire [31:0] _EVAL_2089;
  wire  _EVAL_2090;
  wire  _EVAL_2091;
  wire  _EVAL_2092;
  wire [31:0] _EVAL_2095;
  wire [31:0] _EVAL_2096;
  wire  _EVAL_2097;
  wire  _EVAL_2101;
  wire  _EVAL_2102;
  wire  _EVAL_2103;
  wire  _EVAL_2104;
  wire [31:0] _EVAL_2106;
  wire [31:0] _EVAL_2110;
  wire  _EVAL_2111;
  wire  _EVAL_2113;
  wire  _EVAL_2115;
  wire  _EVAL_2116;
  wire  _EVAL_2120;
  wire  _EVAL_2121;
  wire [31:0] _EVAL_2125;
  wire  _EVAL_2128;
  wire [31:0] _EVAL_2130;
  wire  _EVAL_2136;
  wire [2:0] _EVAL_2138;
  wire [31:0] _EVAL_2143;
  wire [31:0] _EVAL_2144;
  wire  _EVAL_2145;
  wire  _EVAL_2149;
  wire  _EVAL_2156;
  wire  _EVAL_2157;
  wire [31:0] _EVAL_2160;
  wire  _EVAL_2162;
  wire [15:0] _EVAL_2163;
  wire  _EVAL_2166;
  wire  _EVAL_2168;
  wire [31:0] _EVAL_2173;
  wire  _EVAL_2174;
  wire  _EVAL_2175;
  wire  _EVAL_2177;
  wire  _EVAL_2178;
  wire  _EVAL_2183;
  wire  _EVAL_2185;
  wire  _EVAL_2188;
  wire  _EVAL_2190;
  wire [31:0] _EVAL_2193;
  wire [31:0] _EVAL_2194;
  wire  _EVAL_2196;
  wire  _EVAL_2207;
  wire [31:0] _EVAL_2210;
  wire  _EVAL_2211;
  wire [31:0] _EVAL_2216;
  wire [31:0] _EVAL_2217;
  reg  _EVAL_2218;
  reg [31:0] _RAND_11;
  wire  _EVAL_2219;
  wire  _EVAL_2220;
  wire [31:0] _EVAL_2222;
  wire [31:0] _EVAL_2223;
  wire [31:0] _EVAL_2224;
  wire [31:0] _EVAL_2233;
  wire  _EVAL_2235;
  wire  _EVAL_2237;
  wire [31:0] _EVAL_2238;
  wire  _EVAL_2246;
  wire [31:0] _EVAL_2247;
  wire [31:0] _EVAL_2248;
  wire [31:0] _EVAL_2249;
  wire [31:0] _EVAL_2251;
  wire [11:0] _EVAL_2254;
  wire [31:0] _EVAL_2255;
  wire  _EVAL_2256;
  wire [7:0] _EVAL_2261;
  wire  _EVAL_2262;
  wire [7:0] _EVAL_2264;
  wire  _EVAL_2265;
  wire [31:0] _EVAL_2268;
  wire  _EVAL_2272;
  wire [31:0] _EVAL_2274;
  wire [31:0] _EVAL_2277;
  wire  _EVAL_2279;
  wire [7:0] _EVAL_2280;
  wire [31:0] _EVAL_2284;
  wire  _EVAL_2285;
  wire [31:0] _EVAL_2286;
  wire  _EVAL_2290;
  wire  _EVAL_2291;
  wire  _EVAL_2294;
  wire [31:0] _EVAL_2295;
  wire [31:0] _EVAL_2299;
  wire  _EVAL_2302;
  wire [31:0] _EVAL_2306;
  wire  _EVAL_2308;
  wire  _EVAL_2311;
  wire  _EVAL_2312;
  wire [31:0] _EVAL_2314;
  wire  _EVAL_2317;
  wire  _EVAL_2318;
  wire  _EVAL_2324;
  wire  _EVAL_2325;
  wire [31:0] _EVAL_2326;
  wire  _EVAL_2332;
  wire  _EVAL_2333;
  wire [31:0] _EVAL_2334;
  wire  _EVAL_2336;
  wire  _EVAL_2339;
  wire  _EVAL_2340;
  wire  _EVAL_2343;
  wire [7:0] _EVAL_2344;
  wire  _EVAL_2347;
  wire [31:0] _EVAL_2351;
  wire  _EVAL_2354;
  wire  _EVAL_2358;
  wire  _EVAL_2359;
  wire [31:0] _EVAL_2360;
  wire [31:0] _EVAL_2363;
  wire [31:0] _EVAL_2365;
  wire  _EVAL_2366;
  wire [31:0] _EVAL_2367;
  wire [31:0] _EVAL_2368;
  wire [31:0] _EVAL_2371;
  wire  _EVAL_2373;
  wire [31:0] _EVAL_2378;
  wire  _EVAL_2379;
  wire  _EVAL_2383;
  wire [31:0] _EVAL_2384;
  wire  _EVAL_2387;
  wire  _EVAL_2390;
  wire [31:0] _EVAL_2392;
  wire  _EVAL_2395;
  wire  _EVAL_2398;
  wire [31:0] _EVAL_2399;
  wire  _EVAL_2400;
  wire  _EVAL_2402;
  wire  _EVAL_2403;
  wire  _EVAL_2410;
  wire  _EVAL_2411;
  wire  _EVAL_2412;
  wire  _EVAL_2414;
  wire [31:0] _EVAL_2417;
  wire  _EVAL_2418;
  wire  _EVAL_2419;
  wire [7:0] _EVAL_2420;
  wire  _EVAL_2422;
  wire [31:0] _EVAL_2429;
  wire [31:0] _EVAL_2432;
  wire  _EVAL_2437;
  wire  _EVAL_2438;
  wire [31:0] _EVAL_2440;
  wire  _EVAL_2445;
  wire [31:0] _EVAL_2447;
  wire  _EVAL_2451;
  wire [31:0] _EVAL_2452;
  wire  _EVAL_2453;
  wire  _EVAL_2455;
  wire [31:0] _EVAL_2456;
  wire [31:0] _EVAL_2457;
  wire [23:0] _EVAL_2458;
  wire [31:0] _EVAL_2459;
  wire [31:0] _EVAL_2463;
  wire [31:0] _EVAL_2471;
  wire  _EVAL_2472;
  wire [31:0] _EVAL_2476;
  wire  _EVAL_2479;
  wire [31:0] _EVAL_2480;
  wire  _EVAL_2481;
  wire [31:0] _EVAL_2482;
  wire  _EVAL_2484;
  wire  _EVAL_2485;
  wire  _EVAL_2486;
  wire [28:0] _EVAL_2487;
  wire  _EVAL_2488;
  wire [31:0] _EVAL_2489;
  wire  _EVAL_2491;
  wire [31:0] _EVAL_2494;
  wire [31:0] _EVAL_2495;
  wire [31:0] _EVAL_2496;
  wire  _EVAL_2497;
  wire  _EVAL_2499;
  wire  _EVAL_2501;
  wire [31:0] _EVAL_2503;
  wire  _EVAL_2504;
  wire [31:0] _EVAL_2506;
  wire [31:0] _EVAL_2508;
  wire [31:0] _EVAL_2512;
  wire [31:0] _EVAL_2517;
  wire  _EVAL_2519;
  wire  _EVAL_2520;
  wire  _EVAL_2522;
  wire  _EVAL_2524;
  wire  _EVAL_2527;
  wire  _EVAL_2532;
  wire  _EVAL_2533;
  wire [1:0] _EVAL_2538;
  wire  _EVAL_2540;
  wire [31:0] _EVAL_2544;
  wire  _EVAL_2552;
  wire [31:0] _EVAL_2558;
  wire  _EVAL_2560;
  wire  _EVAL_2565;
  wire  _EVAL_2566;
  wire  _EVAL_2569;
  wire [31:0] _EVAL_2570;
  wire  _EVAL_2571;
  wire  _EVAL_2573;
  wire [31:0] _EVAL_2578;
  wire  _EVAL_2581;
  wire  _EVAL_2583;
  wire [31:0] _EVAL_2584;
  wire [31:0] _EVAL_2588;
  wire  _EVAL_2589;
  wire  _EVAL_2590;
  wire [31:0] _EVAL_2591;
  wire  _EVAL_2593;
  wire  _EVAL_2594;
  wire  _EVAL_2595;
  wire  _EVAL_2598;
  wire  _EVAL_2602;
  wire  _EVAL_2604;
  wire  _EVAL_2610;
  wire [31:0] _EVAL_2611;
  wire [31:0] _EVAL_2615;
  wire [31:0] _EVAL_2616;
  wire [31:0] _EVAL_2619;
  wire  _EVAL_2623;
  wire [2:0] _EVAL_2624;
  wire  _EVAL_2627;
  wire [2:0] _EVAL_2628;
  wire  _EVAL_2629;
  wire  _EVAL_2631;
  wire  _EVAL_2635;
  wire  _EVAL_2636;
  wire  _EVAL_2641;
  wire  _EVAL_2642;
  wire  _EVAL_2643;
  wire  _EVAL_2648;
  wire  _EVAL_2650;
  wire  _EVAL_2651;
  wire [31:0] _EVAL_2653;
  wire  _EVAL_2655;
  wire [31:0] _EVAL_2659;
  wire [7:0] _EVAL_2662;
  wire  _EVAL_2673;
  wire  _EVAL_2674;
  wire  _EVAL_2683;
  wire  _EVAL_2684;
  wire [31:0] _EVAL_2686;
  wire [31:0] _EVAL_2687;
  wire  _EVAL_2688;
  wire  _EVAL_2689;
  wire  _EVAL_2691;
  wire  _EVAL_2695;
  wire [31:0] _EVAL_2697;
  wire  _EVAL_2698;
  wire [31:0] _EVAL_2699;
  wire  _EVAL_2700;
  wire  _EVAL_2703;
  wire  _EVAL_2704;
  wire  _EVAL_2705;
  wire [31:0] _EVAL_2706;
  wire  _EVAL_2707;
  wire  _EVAL_2709;
  wire [7:0] _EVAL_2711;
  wire  _EVAL_2712;
  wire  _EVAL_2713;
  wire  _EVAL_2714;
  wire  _EVAL_2716;
  reg [7:0] _EVAL_2720;
  reg [31:0] _RAND_12;
  wire  _EVAL_2721;
  wire  _EVAL_2724;
  wire  _EVAL_2725;
  wire [7:0] _EVAL_2727;
  wire [31:0] _EVAL_2730;
  wire  _EVAL_2731;
  wire  _EVAL_2732;
  wire [31:0] _EVAL_2735;
  wire [31:0] _EVAL_2736;
  wire [31:0] _EVAL_2737;
  wire  _EVAL_2741;
  wire  _EVAL_2742;
  wire [511:0] _EVAL_2743;
  wire  _EVAL_2744;
  wire  _EVAL_2746;
  wire  _EVAL_2749;
  wire [31:0] _EVAL_2750;
  wire [31:0] _EVAL_2755;
  wire  _EVAL_2756;
  reg [7:0] _EVAL_2757;
  reg [31:0] _RAND_13;
  wire  _EVAL_2758;
  wire  _EVAL_2759;
  wire  _EVAL_2761;
  wire [7:0] _EVAL_2763;
  wire  _EVAL_2769;
  wire [31:0] _EVAL_2770;
  wire  _EVAL_2771;
  wire  _EVAL_2774;
  wire [31:0] _EVAL_2775;
  wire  _EVAL_2777;
  wire [31:0] _EVAL_2780;
  wire  _EVAL_2781;
  wire  _EVAL_2786;
  wire  _EVAL_2788;
  wire [31:0] _EVAL_2789;
  wire [31:0] _EVAL_2791;
  wire [31:0] _EVAL_2794;
  wire  _EVAL_2797;
  wire  _EVAL_2801;
  wire [31:0] _EVAL_2804;
  wire  _EVAL_2807;
  wire [31:0] _EVAL_2809;
  wire  _EVAL_2810;
  wire  _EVAL_2811;
  wire [31:0] _EVAL_2812;
  wire [31:0] _EVAL_2816;
  wire [31:0] _EVAL_2818;
  wire  _EVAL_2819;
  wire [31:0] _EVAL_2820;
  wire [31:0] _EVAL_2821;
  wire  _EVAL_2822;
  wire  _EVAL_2828;
  wire [31:0] _EVAL_2829;
  wire  _EVAL_2831;
  wire  _EVAL_2836;
  wire  _EVAL_2837;
  wire  _EVAL_2838;
  wire  _EVAL_2840;
  wire  _EVAL_2841;
  wire [31:0] _EVAL_2842;
  wire  _EVAL_2843;
  wire  _EVAL_2845;
  wire  _EVAL_2847;
  wire [31:0] _EVAL_2850;
  wire  _EVAL_2851;
  wire  _EVAL_2853;
  wire [31:0] _EVAL_2854;
  wire  _EVAL_2855;
  wire  _EVAL_2858;
  wire [2:0] _EVAL_2861;
  wire  _EVAL_2862;
  wire [7:0] _EVAL_2864;
  wire [31:0] _EVAL_2870;
  wire  _EVAL_2871;
  wire  _EVAL_2878;
  wire  _EVAL_2879;
  wire  _EVAL_2881;
  wire [31:0] _EVAL_2882;
  wire  _EVAL_2883;
  wire  _EVAL_2885;
  wire  _EVAL_2886;
  wire  _EVAL_2887;
  wire  _EVAL_2888;
  wire [31:0] _EVAL_2890;
  wire  _EVAL_2893;
  wire [31:0] _EVAL_2894;
  wire [31:0] _EVAL_2895;
  wire  _EVAL_2896;
  wire  _EVAL_2899;
  reg [7:0] _EVAL_2905;
  reg [31:0] _RAND_14;
  wire [31:0] _EVAL_2908;
  wire  _EVAL_2911;
  wire [31:0] _EVAL_2913;
  wire [31:0] _EVAL_2915;
  wire  _EVAL_2920;
  wire  _EVAL_2921;
  wire [31:0] _EVAL_2927;
  wire [31:0] _EVAL_2928;
  wire  _EVAL_2929;
  wire [31:0] _EVAL_2932;
  wire [31:0] _EVAL_2934;
  wire  _EVAL_2937;
  wire [31:0] _EVAL_2938;
  wire  _EVAL_2939;
  wire [31:0] _EVAL_2945;
  wire [20:0] _EVAL_2948;
  wire  _EVAL_2951;
  wire  _EVAL_2955;
  wire  _EVAL_2956;
  wire [15:0] _EVAL_2957;
  wire  _EVAL_2958;
  wire  _EVAL_2959;
  wire  _EVAL_2961;
  wire  _EVAL_2964;
  wire  _EVAL_2965;
  wire  _EVAL_2970;
  wire  _EVAL_2974;
  wire [31:0] _EVAL_2977;
  reg  _EVAL_2978;
  reg [31:0] _RAND_15;
  wire [31:0] _EVAL_2979;
  wire  _EVAL_2986;
  reg  _EVAL_2987;
  reg [31:0] _RAND_16;
  wire  _EVAL_2988;
  wire [31:0] _EVAL_2989;
  wire  _EVAL_2992;
  wire  _EVAL_2994;
  wire [31:0] _EVAL_2995;
  wire  _EVAL_2996;
  reg [31:0] _EVAL_3000;
  reg [31:0] _RAND_17;
  wire  _EVAL_3001;
  wire [31:0] _EVAL_3002;
  wire  _EVAL_3003;
  wire [31:0] _EVAL_3004;
  wire  _EVAL_3005;
  wire  _EVAL_3009;
  wire  _EVAL_3011;
  wire [31:0] _EVAL_3013;
  wire [31:0] _EVAL_3017;
  wire  _EVAL_3020;
  wire [31:0] _EVAL_3021;
  wire  _EVAL_3022;
  wire  _EVAL_3023;
  wire [31:0] _EVAL_3025;
  wire  _EVAL_3026;
  wire  _EVAL_3027;
  wire  _EVAL_3030;
  wire [31:0] _EVAL_3031;
  wire [31:0] _EVAL_3035;
  wire  _EVAL_3038;
  wire  _EVAL_3039;
  wire  _EVAL_3043;
  wire  _EVAL_3045;
  wire  _EVAL_3046;
  wire  _EVAL_3047;
  reg [7:0] _EVAL_3050;
  reg [31:0] _RAND_18;
  wire [31:0] _EVAL_3052;
  wire [31:0] _EVAL_3059;
  wire [31:0] _EVAL_3061;
  wire [31:0] _EVAL_3064;
  wire  _EVAL_3065;
  reg  _EVAL_3066;
  reg [31:0] _RAND_19;
  wire [31:0] _EVAL_3067;
  wire  _EVAL_3068;
  wire  _EVAL_3069;
  wire  _EVAL_3070;
  wire [31:0] _EVAL_3071;
  wire [31:0] _EVAL_3073;
  wire  _EVAL_3076;
  wire [31:0] _EVAL_3083;
  wire  _EVAL_3085;
  wire [31:0] _EVAL_3087;
  wire [31:0] _EVAL_3088;
  wire  _EVAL_3090;
  wire [31:0] _EVAL_3093;
  wire  _EVAL_3094;
  wire [31:0] _EVAL_3095;
  wire  _EVAL_3096;
  wire [31:0] _EVAL_3097;
  wire  _EVAL_3100;
  wire  _EVAL_3101;
  wire [7:0] _EVAL_3102;
  wire  _EVAL_3103;
  wire  _EVAL_3104;
  reg  _EVAL_3105;
  reg [31:0] _RAND_20;
  wire  _EVAL_3106;
  wire [7:0] _EVAL_3113;
  wire  _EVAL_3115;
  wire [7:0] _EVAL_3116;
  wire  _EVAL_3119;
  wire  _EVAL_3122;
  wire [31:0] _EVAL_3123;
  wire  _EVAL_3127;
  wire  _EVAL_3128;
  wire  _EVAL_3129;
  wire  _EVAL_3132;
  wire  _EVAL_3134;
  wire  _EVAL_3135;
  reg [7:0] _EVAL_3138;
  reg [31:0] _RAND_21;
  wire [31:0] _EVAL_3140;
  wire [7:0] _EVAL_3143;
  wire  _EVAL_3144;
  wire [31:0] _EVAL_3145;
  wire [31:0] _EVAL_3146;
  wire  _EVAL_3148;
  wire [15:0] _EVAL_3152;
  wire  _EVAL_3154;
  wire  _EVAL_3155;
  wire [31:0] _EVAL_3157;
  wire  _EVAL_3159;
  wire  _EVAL_3160;
  wire  _EVAL_3165;
  wire  _EVAL_3169;
  wire  _EVAL_3171;
  wire [31:0] _EVAL_3173;
  wire  _EVAL_3174;
  wire  _EVAL_3176;
  wire  _EVAL_3177;
  wire  _EVAL_3178;
  wire [31:0] _EVAL_3179;
  wire  _EVAL_3182;
  wire  _EVAL_3183;
  wire [31:0] _EVAL_3187;
  wire  _EVAL_3189;
  wire [31:0] _EVAL_3193;
  wire [31:0] _EVAL_3194;
  wire  _EVAL_3195;
  wire  _EVAL_3196;
  wire [31:0] _EVAL_3200;
  wire  _EVAL_3203;
  wire [31:0] _EVAL_3207;
  wire  _EVAL_3209;
  wire  _EVAL_3212;
  wire  _EVAL_3217;
  wire [31:0] _EVAL_3219;
  wire [31:0] _EVAL_3220;
  wire  _EVAL_3221;
  wire  _EVAL_3223;
  wire  _EVAL_3227;
  wire [31:0] _EVAL_3228;
  wire  _EVAL_3230;
  wire [31:0] _EVAL_3231;
  wire  _EVAL_3233;
  wire  _EVAL_3234;
  wire  _EVAL_3235;
  wire  _EVAL_3236;
  wire  _EVAL_3237;
  wire  _EVAL_3238;
  wire [31:0] _EVAL_3239;
  wire  _EVAL_3241;
  wire [7:0] _EVAL_3244;
  wire  _EVAL_3246;
  wire  _EVAL_3247;
  wire  _EVAL_3249;
  wire [31:0] _EVAL_3250;
  wire  _EVAL_3251;
  wire  _EVAL_3252;
  wire  _EVAL_3254;
  wire  _EVAL_3259;
  wire  _EVAL_3262;
  wire  _EVAL_3264;
  wire [31:0] _EVAL_3265;
  wire  _EVAL_3268;
  wire [31:0] _EVAL_3270;
  wire [31:0] _EVAL_3271;
  wire [31:0] _EVAL_3275;
  wire [31:0] _EVAL_3276;
  wire [31:0] _EVAL_3279;
  wire  _EVAL_3280;
  wire  _EVAL_3281;
  wire  _EVAL_3283;
  wire [31:0] _EVAL_3288;
  wire  _EVAL_3290;
  wire [31:0] _EVAL_3295;
  wire  _EVAL_3298;
  wire  _EVAL_3299;
  wire [31:0] _EVAL_3302;
  wire  _EVAL_3306;
  wire [31:0] _EVAL_3309;
  wire  _EVAL_3310;
  wire [31:0] _EVAL_3316;
  wire [31:0] _EVAL_3318;
  wire [31:0] _EVAL_3320;
  wire [31:0] _EVAL_3321;
  wire  _EVAL_3322;
  wire  _EVAL_3323;
  wire  _EVAL_3325;
  wire [31:0] _EVAL_3326;
  wire  _EVAL_3328;
  wire [31:0] _EVAL_3329;
  wire  _EVAL_3331;
  wire [6:0] _EVAL_3337;
  wire  _EVAL_3338;
  wire  _EVAL_3339;
  wire  _EVAL_3342;
  wire  _EVAL_3343;
  reg [31:0] _EVAL_3348;
  reg [31:0] _RAND_22;
  wire [31:0] _EVAL_3349;
  wire  _EVAL_3356;
  wire [31:0] _EVAL_3359;
  wire  _EVAL_3366;
  wire  _EVAL_3369;
  wire [31:0] _EVAL_3372;
  wire [31:0] _EVAL_3377;
  wire  _EVAL_3379;
  wire  _EVAL_3385;
  wire [31:0] _EVAL_3387;
  wire  _EVAL_3388;
  wire  _EVAL_3389;
  wire [7:0] _EVAL_3390;
  wire  _EVAL_3393;
  wire  _EVAL_3395;
  reg  _EVAL_3402;
  reg [31:0] _RAND_23;
  wire [31:0] _EVAL_3403;
  wire [31:0] _EVAL_3404;
  wire  _EVAL_3408;
  wire [31:0] _EVAL_3409;
  wire [31:0] _EVAL_3411;
  wire  _EVAL_3417;
  wire  _EVAL_3418;
  wire  _EVAL_3420;
  wire [31:0] _EVAL_3421;
  wire  _EVAL_3423;
  wire  _EVAL_3425;
  wire  _EVAL_3426;
  wire  _EVAL_3427;
  wire [31:0] _EVAL_3428;
  wire  _EVAL_3429;
  wire  _EVAL_3431;
  reg [7:0] _EVAL_3433;
  reg [31:0] _RAND_24;
  wire  _EVAL_3436;
  wire  _EVAL_3442;
  wire  _EVAL_3444;
  wire  _EVAL_3447;
  wire  _EVAL_3448;
  wire  _EVAL_3452;
  wire [31:0] _EVAL_3454;
  wire  _EVAL_3456;
  wire  _EVAL_3457;
  wire  _EVAL_3458;
  wire [31:0] _EVAL_3459;
  wire  _EVAL_3461;
  wire [31:0] _EVAL_3464;
  wire  _EVAL_3465;
  wire [31:0] _EVAL_3469;
  wire  _EVAL_3470;
  wire  _EVAL_3472;
  wire [7:0] _EVAL_3474;
  wire  _EVAL_3475;
  wire [31:0] _EVAL_3476;
  wire  _EVAL_3480;
  wire  _EVAL_3481;
  wire  _EVAL_3482;
  wire  _EVAL_3485;
  wire  _EVAL_3487;
  wire  _EVAL_3490;
  wire [31:0] _EVAL_3493;
  wire [31:0] _EVAL_3495;
  wire  _EVAL_3496;
  wire  _EVAL_3498;
  wire [31:0] _EVAL_3499;
  wire [31:0] _EVAL_3500;
  wire  _EVAL_3502;
  wire [31:0] _EVAL_3504;
  wire [31:0] _EVAL_3506;
  wire  _EVAL_3507;
  wire  _EVAL_3508;
  wire  _EVAL_3509;
  wire  _EVAL_3511;
  wire [31:0] _EVAL_3513;
  wire  _EVAL_3515;
  wire  _EVAL_3517;
  wire [1:0] _EVAL_3518;
  wire  _EVAL_3519;
  wire [31:0] _EVAL_3520;
  wire  _EVAL_3524;
  wire [31:0] _EVAL_3526;
  wire  _EVAL_3530;
  wire  _EVAL_3531;
  wire  _EVAL_3535;
  wire  _EVAL_3537;
  wire [31:0] _EVAL_3539;
  wire  _EVAL_3540;
  wire  _EVAL_3541;
  wire [31:0] _EVAL_3542;
  wire  _EVAL_3545;
  wire [31:0] _EVAL_3549;
  wire  _EVAL_3551;
  wire  _EVAL_3555;
  wire  _EVAL_3557;
  wire [6:0] _EVAL_3558;
  wire [31:0] _EVAL_3566;
  wire  _EVAL_3567;
  wire  _EVAL_3568;
  wire  _EVAL_3569;
  wire  _EVAL_3574;
  wire  _EVAL_3576;
  wire  _EVAL_3577;
  wire [31:0] _EVAL_3583;
  wire  _EVAL_3586;
  wire  _EVAL_3588;
  wire [31:0] _EVAL_3589;
  wire [31:0] _EVAL_3590;
  wire [31:0] _EVAL_3591;
  wire  _EVAL_3593;
  wire  _EVAL_3595;
  wire  _EVAL_3596;
  wire [31:0] _EVAL_3598;
  wire [31:0] _EVAL_3599;
  wire  _EVAL_3600;
  wire  _EVAL_3603;
  wire [31:0] _EVAL_3604;
  wire  _EVAL_3606;
  wire  _EVAL_3609;
  wire  _EVAL_3610;
  wire  _EVAL_3612;
  wire  _EVAL_3613;
  wire  _EVAL_3614;
  wire [31:0] _EVAL_3623;
  wire  _EVAL_3633;
  wire  _EVAL_3634;
  wire [31:0] _EVAL_3637;
  wire  _EVAL_3641;
  wire [31:0] _EVAL_3644;
  wire [31:0] _EVAL_3647;
  wire  _EVAL_3649;
  wire [31:0] _EVAL_3650;
  wire  _EVAL_3651;
  wire  _EVAL_3652;
  wire  _EVAL_3653;
  wire  _EVAL_3654;
  wire [31:0] _EVAL_3657;
  wire [31:0] _EVAL_3661;
  wire  _EVAL_3662;
  wire  _EVAL_3663;
  wire  _EVAL_3666;
  wire  _EVAL_3668;
  wire  _EVAL_3669;
  wire  _EVAL_3670;
  wire [31:0] _EVAL_3671;
  wire  _EVAL_3672;
  wire [31:0] _EVAL_3675;
  wire [31:0] _EVAL_3676;
  wire [31:0] _EVAL_3677;
  wire [31:0] _EVAL_3682;
  wire [31:0] _EVAL_3687;
  wire [31:0] _EVAL_3688;
  wire  _EVAL_3689;
  wire  _EVAL_3694;
  wire [31:0] _EVAL_3695;
  wire  _EVAL_3698;
  wire  _EVAL_3700;
  wire  _EVAL_3701;
  wire [31:0] _EVAL_3703;
  wire  _EVAL_3704;
  wire  _EVAL_3707;
  wire [31:0] _EVAL_3709;
  wire  _EVAL_3710;
  wire  _EVAL_3711;
  wire  _EVAL_3714;
  wire  _EVAL_3717;
  wire  _EVAL_3722;
  wire  _EVAL_3723;
  wire  _EVAL_3724;
  wire  _EVAL_3725;
  wire  _EVAL_3727;
  wire  _EVAL_3731;
  wire  _EVAL_3736;
  wire [31:0] _EVAL_3738;
  wire [31:0] _EVAL_3739;
  wire [31:0] _EVAL_3741;
  wire  _EVAL_3742;
  wire  _EVAL_3743;
  wire  _EVAL_3745;
  wire  _EVAL_3746;
  wire [31:0] _EVAL_3748;
  wire [7:0] _EVAL_3750;
  wire  _EVAL_3751;
  wire  _EVAL_3753;
  wire [31:0] _EVAL_3754;
  wire  _EVAL_3755;
  wire  _EVAL_3761;
  wire  _EVAL_3762;
  wire  _EVAL_3763;
  wire  _EVAL_3764;
  wire  _EVAL_3769;
  wire [7:0] _EVAL_3770;
  wire  _EVAL_3772;
  wire [31:0] _EVAL_3774;
  wire  _EVAL_3775;
  wire  _EVAL_3776;
  reg [7:0] _EVAL_3777;
  reg [31:0] _RAND_25;
  wire  _EVAL_3782;
  wire  _EVAL_3783;
  wire  _EVAL_3784;
  wire  _EVAL_3788;
  wire [31:0] _EVAL_3791;
  wire  _EVAL_3795;
  wire  _EVAL_3799;
  wire [31:0] _EVAL_3800;
  wire [31:0] _EVAL_3804;
  wire  _EVAL_3806;
  wire  _EVAL_3807;
  wire  _EVAL_3809;
  wire  _EVAL_3811;
  wire  _EVAL_3813;
  wire  _EVAL_3814;
  wire  _EVAL_3815;
  wire  _EVAL_3816;
  wire  _EVAL_3823;
  wire  _EVAL_3824;
  wire  _EVAL_3825;
  wire  _EVAL_3826;
  wire  _EVAL_3829;
  wire [31:0] _EVAL_3830;
  wire  _EVAL_3832;
  wire [31:0] _EVAL_3834;
  wire  _EVAL_3836;
  wire  _EVAL_3837;
  wire  _EVAL_3838;
  wire  _EVAL_3839;
  wire  _EVAL_3841;
  _EVAL_140 debug_hartReset_0 (
    ._EVAL(debug_hartReset_0__EVAL),
    ._EVAL_0(debug_hartReset_0__EVAL_0),
    ._EVAL_1(debug_hartReset_0__EVAL_1),
    ._EVAL_2(debug_hartReset_0__EVAL_2)
  );
  assign _EVAL_2629 = 9'hc7 == _EVAL_1399;
  assign _EVAL_1261 = _EVAL_797 | _EVAL_3431;
  assign _EVAL_1465 = 9'h4c == _EVAL_1399 ? 32'h0 : _EVAL_930;
  assign _EVAL_2929 = 9'h92 == _EVAL_1399;
  assign _EVAL_2636 = 9'h178 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1138;
  assign _EVAL_285 = 9'h136 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3389;
  assign _EVAL_2302 = ~_EVAL_3155;
  assign _EVAL_3238 = 9'h10e == _EVAL_1399 ? _EVAL_1856 : _EVAL_2713;
  assign _EVAL_1989 = 9'h70 == _EVAL_1399;
  assign _EVAL_1071 = 9'h1d6 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2705;
  assign _EVAL_3194 = 9'h128 == _EVAL_1399 ? _EVAL_374 : _EVAL_1377;
  assign _EVAL_1125 = 9'h19 == _EVAL_1399 ? 32'h0 : _EVAL_1547;
  assign _EVAL_3649 = _EVAL_2727 != 8'h0;
  assign _EVAL_542 = 9'h1eb == _EVAL_1399 ? _EVAL_1856 : _EVAL_225;
  assign _EVAL_1871 = _EVAL_642 & _EVAL_473;
  assign _EVAL_334 = 9'h7e == _EVAL_1399;
  assign _EVAL_851 = _EVAL_1972 | _EVAL_1010;
  assign _EVAL_2566 = _EVAL_3634 | _EVAL_3541;
  assign _EVAL_3096 = _EVAL_679 | _EVAL_3127;
  assign _EVAL_3323 = 9'h1bb == _EVAL_1399 ? _EVAL_1856 : _EVAL_2689;
  assign _EVAL_1163 = 9'ha0 == _EVAL_1399;
  assign _EVAL_497 = _EVAL_2290 | _EVAL_3799;
  assign _EVAL_612 = _EVAL_575[17:16];
  assign _EVAL_2438 = 9'h6f == _EVAL_1399;
  assign _EVAL_2697 = 9'h1e9 == _EVAL_1399 ? _EVAL_374 : _EVAL_3083;
  assign _EVAL_1194 = _EVAL_512 | _EVAL_1145;
  assign _EVAL_51 = 9'h14 == _EVAL_1399 ? 32'h100073 : _EVAL_3004;
  assign _EVAL_4 = {{2'd0}, _EVAL_2004};
  assign _EVAL_2168 = _EVAL_2018 | _EVAL_2061;
  assign _EVAL_202 = 9'hcc == _EVAL_1399;
  assign _EVAL_3811 = _EVAL_3283 | _EVAL_2641;
  assign _EVAL_2371 = 9'hc5 == _EVAL_1399 ? 32'h0 : _EVAL_3703;
  assign _EVAL_1622 = 9'hf2 == _EVAL_1399 ? 32'h0 : _EVAL_1392;
  assign _EVAL_3179 = 9'h1a8 == _EVAL_1399 ? _EVAL_374 : _EVAL_2130;
  assign _EVAL_3339 = _EVAL_3672 | _EVAL_3784;
  assign _EVAL_1593 = 9'hb1 == _EVAL_1399 ? 32'h0 : _EVAL_2775;
  assign _EVAL_1844 = 9'h195 == _EVAL_1399 ? _EVAL_374 : _EVAL_58;
  assign _EVAL_3677 = {_EVAL_167,_EVAL_2957};
  assign _EVAL_1021 = 9'hb == _EVAL_1399 ? _EVAL_3670 : _EVAL_1420;
  assign _EVAL_468 = _EVAL_1939 & _EVAL_2749;
  assign _EVAL_3134 = 9'h8f == _EVAL_1399;
  assign _EVAL_2642 = 9'h14 == _EVAL_1399 ? _EVAL_3670 : _EVAL_178;
  assign _EVAL_175 = 9'h4e == _EVAL_1399 ? 32'h0 : _EVAL_1587;
  assign _EVAL_3517 = 9'h6e == _EVAL_1399;
  assign _EVAL_3209 = 9'hed == _EVAL_1399;
  assign _EVAL_3178 = 9'h5d == _EVAL_1399;
  assign _EVAL_2211 = _EVAL_1572 | _EVAL_861;
  assign _EVAL_182 = 9'ha6 == _EVAL_1399 ? 32'h0 : _EVAL_3774;
  assign _EVAL_1018 = ~_EVAL_2673;
  assign _EVAL_605 = 9'hd5 == _EVAL_1399 ? 32'h0 : _EVAL_1832;
  assign _EVAL_270 = 9'hf7 == _EVAL_1399 ? 32'h0 : _EVAL_2791;
  assign _EVAL_233 = 9'h73 == _EVAL_1399;
  assign _EVAL_1334 = 9'h3 == _EVAL_1399 ? _EVAL_3670 : _EVAL_79;
  assign _EVAL_3589 = 9'h1ab == _EVAL_1399 ? _EVAL_374 : _EVAL_2440;
  assign _EVAL_926 = _EVAL_1273 & _EVAL_2836;
  assign _EVAL_3290 = _EVAL_1567 | _EVAL_3237;
  assign _EVAL_1684 = 9'h17 == _EVAL_1399;
  assign _EVAL_3349 = _EVAL_793 ? 32'h111380 : _EVAL_3495;
  assign _EVAL_2429 = 9'h1e == _EVAL_1399 ? 32'h0 : _EVAL_2890;
  assign _EVAL_616 = _EVAL_3207[18];
  assign _EVAL_3343 = 9'hab == _EVAL_1399;
  assign _EVAL_3423 = _EVAL_2403 & _EVAL_3485;
  assign _EVAL_1010 = _EVAL_1304 | _EVAL_3811;
  assign _EVAL_2957 = {{14'd0}, _EVAL_3518};
  assign _EVAL_1084 = 9'h8d == _EVAL_1399 ? 32'h0 : _EVAL_1351;
  assign _EVAL_1931 = 9'hb5 == _EVAL_1399;
  assign _EVAL_3076 = 9'h11a == _EVAL_1399 ? _EVAL_1856 : _EVAL_2648;
  assign _EVAL_2540 = _EVAL_3 == 10'h0;
  assign _EVAL_1603 = 9'hf2 == _EVAL_1399;
  assign _EVAL_3603 = 9'hc0 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2102;
  assign _EVAL_3657 = 9'h2c == _EVAL_1399 ? 32'h0 : _EVAL_2495;
  assign _EVAL_2340 = _EVAL_1251 | _EVAL_2149;
  assign _EVAL_3507 = _EVAL_1367 & _EVAL_1303;
  assign _EVAL_1968 = 9'h57 == _EVAL_1399 ? 32'h0 : _EVAL_611;
  assign _EVAL_448 = 9'hcb == _EVAL_1399;
  assign _EVAL_1863 = _EVAL_554 | _EVAL_1611;
  assign _EVAL_3474 = _EVAL_2363[7:0];
  assign _EVAL_1538 = _EVAL_2285 | _EVAL_759;
  assign _EVAL_2222 = 9'h196 == _EVAL_1399 ? _EVAL_374 : _EVAL_1844;
  assign _EVAL_3761 = _EVAL_2012 == 3'h0;
  assign _EVAL_409 = 9'hab == _EVAL_1399 ? 32'h0 : _EVAL_354;
  assign _EVAL_3070 = 9'h42 == _EVAL_1399 ? _EVAL_1856 : _EVAL_719;
  assign _EVAL_271 = _EVAL_1335 ? 1'h0 : _EVAL_3105;
  assign _EVAL_3476 = 9'h1af == _EVAL_1399 ? _EVAL_374 : _EVAL_949;
  assign _EVAL_533 = 9'h153 == _EVAL_1399 ? _EVAL_374 : _EVAL_2699;
  assign _EVAL_1196 = 9'h1d1 == _EVAL_1399 ? _EVAL_374 : _EVAL_3279;
  assign _EVAL_1273 = _EVAL_1846 & _EVAL_1135;
  assign _EVAL_370 = _EVAL_1326 | _EVAL_1039;
  assign _EVAL_2829 = 9'h52 == _EVAL_1399 ? 32'h0 : _EVAL_3566;
  assign _EVAL_2532 = 9'hb1 == _EVAL_1399;
  assign _EVAL_2014 = _EVAL_248 | _EVAL_2879;
  assign _EVAL_2737 = 9'h190 == _EVAL_1399 ? _EVAL_374 : _EVAL_2770;
  assign _EVAL_847 = 9'h165 == _EVAL_1399 ? _EVAL_1856 : _EVAL_339;
  assign _EVAL_1077 = 9'h18b == _EVAL_1399 ? _EVAL_1856 : _EVAL_2610;
  assign _EVAL_2354 = _EVAL_509 | _EVAL_763;
  assign _EVAL_397 = _EVAL_1183 | _EVAL_3519;
  assign _EVAL_2447 = 9'h160 == _EVAL_1399 ? _EVAL_374 : _EVAL_3329;
  assign _EVAL_795 = 9'h11d == _EVAL_1399 ? _EVAL_1856 : _EVAL_2311;
  assign _EVAL_538 = 9'he3 == _EVAL_1399 ? 32'h0 : _EVAL_2506;
  assign _EVAL_1470 = 9'hee == _EVAL_1399 ? 32'h0 : _EVAL_2015;
  assign _EVAL_1552 = _EVAL_3829 ? 8'hff : 8'h0;
  assign _EVAL_3309 = 9'h39 == _EVAL_1399 ? 32'h0 : _EVAL_3644;
  assign _EVAL_2631 = _EVAL_1666 & _EVAL_2540;
  assign _EVAL_1849 = 9'h73 == _EVAL_1399 ? 32'h0 : _EVAL_3583;
  assign _EVAL_3710 = _EVAL_2174 | _EVAL_1957;
  assign _EVAL_1326 = 9'hd5 == _EVAL_1399;
  assign _EVAL_10 = _EVAL_3420 ? _EVAL_1410 : 32'h0;
  assign _EVAL_3021 = 9'he5 == _EVAL_1399 ? 32'h0 : _EVAL_1641;
  assign _EVAL_1238 = 9'h97 == _EVAL_1399;
  assign _EVAL_3223 = _EVAL_421 & _EVAL_3395;
  assign _EVAL_375 = _EVAL_2235 | _EVAL_2871;
  assign _EVAL_212 = 9'h1c8 == _EVAL_1399 ? _EVAL_374 : _EVAL_1718;
  assign _EVAL_3695 = 9'h189 == _EVAL_1399 ? _EVAL_374 : _EVAL_2334;
  assign _EVAL_3338 = _EVAL_3654 | _EVAL_2742;
  assign _EVAL_3504 = 9'h1e5 == _EVAL_1399 ? _EVAL_374 : _EVAL_179;
  assign _EVAL_912 = 9'ha1 == _EVAL_1399 ? 32'h0 : _EVAL_63;
  assign _EVAL_458 = 9'h14d == _EVAL_1399 ? _EVAL_1856 : _EVAL_2485;
  assign _EVAL_674 = _EVAL_599 | _EVAL_710;
  assign _EVAL_3707 = 9'hd8 == _EVAL_1399;
  assign _EVAL_3183 = 9'h143 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3251;
  assign _EVAL_3189 = 9'h1f0 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3174;
  assign _EVAL_280 = {_EVAL_2336,1'h0,1'h0,1'h0,1'h0,_EVAL_3177,_EVAL_3177,_EVAL_3105,_EVAL_3105,8'ha2};
  assign _EVAL_471 = 9'h7e == _EVAL_1399 ? 32'h0 : _EVAL_1221;
  assign _EVAL_2144 = 9'h10b == _EVAL_1399 ? _EVAL_374 : _EVAL_3321;
  assign _EVAL_2485 = 9'h14c == _EVAL_1399 ? _EVAL_1856 : _EVAL_2565;
  assign _EVAL_559 = 9'h142 == _EVAL_1399 ? _EVAL_374 : _EVAL_2934;
  assign _EVAL_3129 = 9'h36 == _EVAL_1399;
  assign _EVAL_2927 = 9'h16e == _EVAL_1399 ? _EVAL_374 : _EVAL_1133;
  assign _EVAL_822 = 9'h40 == _EVAL_1399 ? _EVAL_1856 : _EVAL_649;
  assign _EVAL_1724 = 9'h165 == _EVAL_1399 ? _EVAL_374 : _EVAL_256;
  assign _EVAL_1759 = 9'h9a == _EVAL_1399;
  assign _EVAL_1097 = 9'h20 == _EVAL_1399;
  assign _EVAL_477 = _EVAL_2939 | _EVAL_2343;
  assign _EVAL_1176 = 5'h9 == _EVAL_958;
  assign _EVAL_1787 = 9'h3d == _EVAL_1399 ? 32'h0 : _EVAL_849;
  assign _EVAL_178 = 9'h13 == _EVAL_1399 ? _EVAL_3670 : _EVAL_3045;
  assign _EVAL_1508 = 9'h1ec == _EVAL_1399 ? _EVAL_1856 : _EVAL_542;
  assign _EVAL_863 = _EVAL_2788 | _EVAL_3106;
  assign _EVAL_1445 = 9'h172 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3586;
  assign _EVAL_1215 = _EVAL_468 & _EVAL_234;
  assign _EVAL_2344 = _EVAL_3085 ? 8'hff : 8'h0;
  assign _EVAL_3654 = 9'h83 == _EVAL_1399;
  assign _EVAL_602 = 9'h109 == _EVAL_1399 ? _EVAL_1856 : _EVAL_730;
  assign _EVAL_257 = 9'h1b9 == _EVAL_1399 ? _EVAL_374 : _EVAL_207;
  assign _EVAL_407 = 9'h3f == _EVAL_1399;
  assign _EVAL_2840 = _EVAL_67 == 8'h0;
  assign _EVAL_3596 = 9'h186 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2744;
  assign _EVAL_3217 = 9'h18c == _EVAL_1399 ? _EVAL_1856 : _EVAL_1077;
  assign _EVAL_2295 = 9'h178 == _EVAL_1399 ? _EVAL_374 : _EVAL_1270;
  assign _EVAL_583 = 9'hd4 == _EVAL_1399;
  assign _EVAL_3574 = 9'ha5 == _EVAL_1399;
  assign _EVAL_607 = 9'hb7 == _EVAL_1399;
  assign _EVAL_3689 = 9'h13e == _EVAL_1399 ? _EVAL_1856 : _EVAL_2899;
  assign _EVAL_1015 = 9'h1bd == _EVAL_1399 ? _EVAL_374 : _EVAL_2006;
  assign _EVAL_722 = 9'h31 == _EVAL_1399 ? 32'h0 : _EVAL_946;
  assign _EVAL_2484 = 9'h17c == _EVAL_1399 ? _EVAL_1856 : _EVAL_431;
  assign _EVAL_1713 = _EVAL_1650 | _EVAL_1423;
  assign _EVAL_1337 = _EVAL_575[0];
  assign _EVAL_2223 = 9'h87 == _EVAL_1399 ? 32'h0 : _EVAL_2913;
  assign _EVAL_434 = 9'h138 == _EVAL_1399 ? _EVAL_374 : _EVAL_2096;
  assign _EVAL_2703 = 9'h104 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2777;
  assign _EVAL_2588 = 9'h67 == _EVAL_1399 ? 32'h0 : _EVAL_2238;
  assign _EVAL_2716 = _EVAL_512 & _EVAL_3610;
  assign _EVAL_2544 = 9'h92 == _EVAL_1399 ? 32'h0 : _EVAL_55;
  assign _EVAL_1358 = _EVAL_1987 != 2'h0;
  assign _EVAL_204 = 9'h9f == _EVAL_1399;
  assign _EVAL_3535 = _EVAL_2631 ? 1'h0 : _EVAL_2987;
  assign _EVAL_1945 = _EVAL_2743[222];
  assign _EVAL_1631 = ~_EVAL_2218;
  assign _EVAL_2383 = 9'h17d == _EVAL_1399 ? _EVAL_1856 : _EVAL_2484;
  assign _EVAL_3165 = 9'hbf == _EVAL_1399;
  assign _EVAL_3230 = _EVAL_1441 | _EVAL_3809;
  assign _EVAL_3389 = 9'h135 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3115;
  assign _EVAL_2519 = 9'h15f == _EVAL_1399 ? _EVAL_1856 : _EVAL_3046;
  assign _EVAL_3227 = 9'h121 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1507;
  assign _EVAL_1587 = 9'h4d == _EVAL_1399 ? 32'h0 : _EVAL_1465;
  assign _EVAL_2591 = 9'he == _EVAL_1399 ? 32'h30000067 : _EVAL_1213;
  assign _EVAL_3322 = 9'h1ee == _EVAL_1399 ? _EVAL_1856 : _EVAL_1461;
  assign _EVAL_3754 = 9'h176 == _EVAL_1399 ? _EVAL_374 : _EVAL_634;
  assign _EVAL_3688 = 9'hb3 == _EVAL_1399 ? 32'h0 : _EVAL_3637;
  assign _EVAL_931 = 9'h182 == _EVAL_1399 ? _EVAL_374 : _EVAL_3231;
  assign _EVAL_1562 = _EVAL_3207[17];
  assign _EVAL_432 = 9'h134 == _EVAL_1399 ? _EVAL_374 : _EVAL_3187;
  assign _EVAL_3480 = 9'h7b == _EVAL_1399;
  assign _EVAL_3241 = 9'h1ce == _EVAL_1399 ? _EVAL_1856 : _EVAL_378;
  assign _EVAL_552 = 9'h159 == _EVAL_1399 ? _EVAL_374 : _EVAL_3830;
  assign _EVAL_3017 = 9'h10 == _EVAL_1399 ? 32'h10802423 : _EVAL_3275;
  assign _EVAL_2584 = 9'h1cc == _EVAL_1399 ? _EVAL_374 : _EVAL_922;
  assign _EVAL_3395 = _EVAL_2840 ? _EVAL_3482 : 1'h1;
  assign _EVAL_1752 = _EVAL_464 & _EVAL_1337;
  assign _EVAL_2964 = 9'h66 == _EVAL_1399;
  assign _EVAL_1958 = 9'h42 == _EVAL_1399 ? 32'h0 : _EVAL_2160;
  assign _EVAL_2029 = _EVAL_642 & _EVAL_1883;
  assign _EVAL_2351 = 9'h154 == _EVAL_1399 ? _EVAL_374 : _EVAL_533;
  assign _EVAL_1191 = _EVAL_642 & _EVAL_1151;
  assign _EVAL_171 = 9'h1cf == _EVAL_1399 ? _EVAL_1856 : _EVAL_3241;
  assign _EVAL_2853 = 9'h1aa == _EVAL_1399 ? _EVAL_1856 : _EVAL_2177;
  assign _EVAL_3807 = _EVAL_3517 | _EVAL_1360;
  assign _EVAL_2673 = _EVAL_3038 & _EVAL_2540;
  assign _EVAL_420 = _EVAL_793 ? _EVAL_2188 : _EVAL_3540;
  assign _EVAL_97 = 9'h1c8 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2801;
  assign _EVAL_2855 = 9'hb9 == _EVAL_1399;
  assign _EVAL_2387 = _EVAL_870[4];
  assign _EVAL_1366 = 9'h24 == _EVAL_1399 ? 32'h0 : _EVAL_1556;
  assign _EVAL_2277 = 9'hcb == _EVAL_1399 ? 32'h0 : _EVAL_3598;
  assign _EVAL_3095 = 9'he8 == _EVAL_1399 ? 32'h0 : _EVAL_3228;
  assign _EVAL_1718 = 9'h1c7 == _EVAL_1399 ? _EVAL_374 : _EVAL_259;
  assign _EVAL_2291 = _EVAL_2402 | _EVAL_2951;
  assign _EVAL_3452 = _EVAL_2743[65];
  assign _EVAL_2106 = 9'h1fa == _EVAL_1399 ? _EVAL_374 : _EVAL_2367;
  assign _EVAL_1965 = 9'h10a == _EVAL_1399 ? _EVAL_1856 : _EVAL_602;
  assign _EVAL_1493 = 9'h56 == _EVAL_1399;
  assign _EVAL_620 = 9'h16b == _EVAL_1399 ? _EVAL_1856 : _EVAL_3176;
  assign _EVAL_66 = 9'h3 == _EVAL_1399 ? 32'hff0000f : _EVAL_3219;
  assign _EVAL_1517 = 9'h1a8 == _EVAL_1399 ? _EVAL_1856 : _EVAL_628;
  assign _EVAL_624 = _EVAL_20 & _EVAL_34;
  assign _EVAL_2707 = 9'he2 == _EVAL_1399;
  assign _EVAL_3623 = 9'hf0 == _EVAL_1399 ? 32'h0 : _EVAL_1477;
  assign _EVAL_3421 = 9'h19f == _EVAL_1399 ? _EVAL_374 : _EVAL_238;
  assign _EVAL_2732 = _EVAL_463 | _EVAL_1541;
  assign _EVAL_1944 = 9'h1fd == _EVAL_1399 ? _EVAL_1856 : _EVAL_2893;
  assign _EVAL_1350 = 9'hfc == _EVAL_1399 ? 32'h0 : _EVAL_1513;
  assign _EVAL_3295 = 9'h1be == _EVAL_1399 ? _EVAL_374 : _EVAL_1015;
  assign _EVAL_1613 = 9'h14c == _EVAL_1399 ? _EVAL_374 : _EVAL_1806;
  assign _EVAL_239 = 9'hba == _EVAL_1399 ? 32'h0 : _EVAL_566;
  assign _EVAL_191 = 9'h50 == _EVAL_1399 ? 32'h0 : _EVAL_223;
  assign _EVAL_3173 = 9'h13b == _EVAL_1399 ? _EVAL_374 : _EVAL_1109;
  assign _EVAL_3465 = 9'hde == _EVAL_1399 ? _EVAL_1856 : _EVAL_2781;
  assign _EVAL_2050 = 9'h1f9 == _EVAL_1399 ? _EVAL_1856 : _EVAL_126;
  assign _EVAL_774 = 9'h1db == _EVAL_1399 ? _EVAL_1856 : _EVAL_519;
  assign _EVAL_968 = 9'h52 == _EVAL_1399;
  assign _EVAL_1530 = 9'hc6 == _EVAL_1399 ? 32'h0 : _EVAL_2371;
  assign _EVAL_1031 = _EVAL_926 | _EVAL_3507;
  assign _EVAL_393 = 9'h104 == _EVAL_1399 ? _EVAL_374 : _EVAL_3513;
  assign _EVAL_2417 = 9'h1ef == _EVAL_1399 ? _EVAL_374 : _EVAL_344;
  assign _EVAL_1506 = _EVAL_2700 | _EVAL_2211;
  assign _EVAL_109 = 9'hc2 == _EVAL_1399 ? 32'h0 : _EVAL_2066;
  assign _EVAL_1240 = 9'h6c == _EVAL_1399;
  assign _EVAL_2066 = 9'hc1 == _EVAL_1399 ? 32'h0 : _EVAL_1677;
  assign _EVAL_1136 = 9'h1f7 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2332;
  assign _EVAL_3746 = _EVAL_334 | _EVAL_754;
  assign _EVAL_3770 = _EVAL_2822 ? 8'hff : 8'h0;
  assign _EVAL_1115 = _EVAL_1472 | _EVAL_2965;
  assign _EVAL_3725 = _EVAL_92 | _EVAL_1928;
  assign _EVAL_3526 = 9'h1f6 == _EVAL_1399 ? _EVAL_374 : _EVAL_2193;
  assign _EVAL_1469 = 9'h29 == _EVAL_1399 ? 32'h0 : _EVAL_3676;
  assign _EVAL_967 = 9'h10d == _EVAL_1399 ? _EVAL_374 : _EVAL_3123;
  assign _EVAL_1549 = 9'hfd == _EVAL_1399;
  assign _EVAL_2883 = 9'h3c == _EVAL_1399;
  assign _EVAL_487 = _EVAL_1589 | _EVAL_1575;
  assign _EVAL_1913 = _EVAL_2743[66];
  assign _EVAL_2286 = 9'h15b == _EVAL_1399 ? _EVAL_374 : _EVAL_417;
  assign _EVAL_1237 = _EVAL_365 | _EVAL_1557;
  assign _EVAL_1742 = 9'h1ca == _EVAL_1399 ? _EVAL_1856 : _EVAL_401;
  assign _EVAL_2004 = _EVAL_13 == 3'h4;
  assign _EVAL_2533 = 9'h1bd == _EVAL_1399 ? _EVAL_1856 : _EVAL_744;
  assign _EVAL_1477 = 9'hef == _EVAL_1399 ? 32'h0 : _EVAL_1470;
  assign _EVAL_463 = 9'hf6 == _EVAL_1399;
  assign _EVAL_2471 = 9'h79 == _EVAL_1399 ? 32'h0 : _EVAL_2482;
  assign _EVAL_1251 = 9'h2b == _EVAL_1399;
  assign _EVAL_2713 = 9'h10d == _EVAL_1399 ? _EVAL_1856 : _EVAL_2520;
  assign _EVAL_991 = _EVAL_1887 ? 8'hff : 8'h0;
  assign _EVAL_2130 = 9'h1a7 == _EVAL_1399 ? _EVAL_374 : _EVAL_2503;
  assign _EVAL_2311 = 9'h11c == _EVAL_1399 ? _EVAL_1856 : _EVAL_2294;
  assign _EVAL_1392 = 9'hf1 == _EVAL_1399 ? 32'h0 : _EVAL_3623;
  assign _EVAL_2487 = {5'h2,_EVAL_282};
  assign _EVAL_2759 = _EVAL_2527 | _EVAL_784;
  assign _EVAL_180 = 9'h127 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2769;
  assign _EVAL_479 = 9'he0 == _EVAL_1399 ? _EVAL_1856 : _EVAL_244;
  assign _EVAL_1887 = _EVAL_29[0];
  assign _EVAL_87 = 9'hf0 == _EVAL_1399;
  assign _EVAL_3837 = 9'h94 == _EVAL_1399;
  assign _EVAL_2843 = 9'h21 == _EVAL_1399;
  assign _EVAL_354 = 9'haa == _EVAL_1399 ? 32'h0 : _EVAL_3316;
  assign _EVAL_3093 = 9'h1fe == _EVAL_1399 ? _EVAL_374 : _EVAL_3302;
  assign _EVAL_1331 = 9'h168 == _EVAL_1399 ? _EVAL_374 : _EVAL_3671;
  assign _EVAL_1269 = 9'h169 == _EVAL_1399 ? _EVAL_374 : _EVAL_1331;
  assign _EVAL_3540 = _EVAL_169 ? _EVAL_2188 : _EVAL_3763;
  assign _EVAL_415 = 9'h118 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2986;
  assign _EVAL_417 = 9'h15a == _EVAL_1399 ? _EVAL_374 : _EVAL_552;
  assign _EVAL_1789 = _EVAL_1174 | _EVAL_3427;
  assign _EVAL_3610 = _EVAL_1778[0];
  assign _EVAL_6 = _EVAL_41;
  assign _EVAL_2102 = _EVAL_3165 | _EVAL_477;
  assign _EVAL_3207 = {_EVAL_67,_EVAL_819};
  assign _EVAL_2002 = 9'h132 == _EVAL_1399 ? _EVAL_374 : _EVAL_1490;
  assign _EVAL_3772 = 9'h58 == _EVAL_1399;
  assign _EVAL_1038 = 9'h163 == _EVAL_1399 ? _EVAL_1856 : _EVAL_846;
  assign _EVAL_3599 = 9'h12b == _EVAL_1399 ? _EVAL_374 : _EVAL_2570;
  assign _EVAL_2570 = 9'h12a == _EVAL_1399 ? _EVAL_374 : _EVAL_1495;
  assign _EVAL_2384 = 9'h3e == _EVAL_1399 ? 32'h0 : _EVAL_1787;
  assign _EVAL_3775 = 5'h10 == _EVAL_958;
  assign _EVAL_1441 = 9'h54 == _EVAL_1399;
  assign _EVAL_519 = 9'h1da == _EVAL_1399 ? _EVAL_1856 : _EVAL_1057;
  assign _EVAL_3104 = _EVAL_1228 ? 1'h0 : 1'h1;
  assign _EVAL_79 = 9'h2 == _EVAL_1399 ? _EVAL_3670 : _EVAL_1175;
  assign _EVAL_1654 = _EVAL_3651 | _EVAL_3448;
  assign _EVAL_1867 = 9'hec == _EVAL_1399;
  assign _EVAL_2018 = _EVAL_3815 & _EVAL_3101;
  assign _EVAL_1244 = 9'h8e == _EVAL_1399 ? 32'h0 : _EVAL_1084;
  assign _EVAL_259 = 9'h1c6 == _EVAL_1399 ? _EVAL_374 : _EVAL_1725;
  assign _EVAL_24 = _EVAL_39;
  assign _EVAL_2828 = _EVAL_563 & _EVAL_3043;
  assign _EVAL_3662 = 5'h8 == _EVAL_958;
  assign _EVAL_3418 = _EVAL_2437 & _EVAL_1913;
  assign _EVAL_2455 = 9'hee == _EVAL_1399;
  assign _EVAL_1121 = _EVAL_3707 | _EVAL_1594;
  assign _EVAL_510 = _EVAL_1759 | _EVAL_2887;
  assign _EVAL_2979 = 9'h17c == _EVAL_1399 ? _EVAL_374 : _EVAL_1755;
  assign _EVAL_1348 = 9'h158 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1407;
  assign _EVAL_3174 = 9'h1ef == _EVAL_1399 ? _EVAL_1856 : _EVAL_3322;
  assign _EVAL_3590 = 9'h6d == _EVAL_1399 ? 32'h0 : _EVAL_2459;
  assign _EVAL_1875 = 9'h17f == _EVAL_1399 ? _EVAL_374 : _EVAL_1150;
  assign _EVAL_3741 = 9'h1a5 == _EVAL_1399 ? _EVAL_374 : _EVAL_3404;
  assign _EVAL_1541 = _EVAL_1833 | _EVAL_1863;
  assign _EVAL_841 = 9'h14f == _EVAL_1399 ? _EVAL_374 : _EVAL_858;
  assign _EVAL_2365 = 9'h6a == _EVAL_1399 ? 32'h0 : _EVAL_2031;
  assign _EVAL_1639 = 9'h6b == _EVAL_1399 ? 32'h0 : _EVAL_2365;
  assign _EVAL_1594 = _EVAL_3704 | _EVAL_832;
  assign _EVAL_1089 = 9'ha9 == _EVAL_1399;
  assign _EVAL_3545 = 9'h16d == _EVAL_1399 ? _EVAL_1856 : _EVAL_569;
  assign _EVAL_1813 = 9'h143 == _EVAL_1399 ? _EVAL_374 : _EVAL_559;
  assign _EVAL_2061 = _EVAL_700 & _EVAL_1380;
  assign _EVAL_2183 = _EVAL_1183 & _EVAL_234;
  assign _EVAL_2001 = 9'hb == _EVAL_1399 ? 32'h40863 : _EVAL_1365;
  assign _EVAL_2552 = 9'h5 == _EVAL_1399 ? _EVAL_3670 : _EVAL_3023;
  assign _EVAL_1583 = 9'h1b == _EVAL_1399 ? 32'h0 : _EVAL_3318;
  assign _EVAL_2249 = 9'h45 == _EVAL_1399 ? 32'h0 : _EVAL_2052;
  assign _EVAL_3128 = 9'h1c4 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3280;
  assign _EVAL_909 = 9'h13e == _EVAL_1399 ? _EVAL_374 : _EVAL_1041;
  assign _EVAL_2602 = 9'h3b == _EVAL_1399;
  assign _EVAL_1045 = _EVAL_320 | _EVAL_867;
  assign _EVAL_1419 = 9'h9a == _EVAL_1399 ? 32'h0 : _EVAL_2457;
  assign _EVAL_1123 = 9'h7c == _EVAL_1399;
  assign _EVAL_2662 = _EVAL_2363[23:16];
  assign _EVAL_2238 = 9'h66 == _EVAL_1399 ? 32'h0 : _EVAL_133;
  assign _EVAL_3557 = 9'h167 == _EVAL_1399 ? _EVAL_1856 : _EVAL_131;
  assign _EVAL_2589 = 9'h159 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1348;
  assign _EVAL_1116 = _EVAL_3551 | _EVAL_1687;
  assign _EVAL_360 = _EVAL_1367 & _EVAL_3649;
  assign _EVAL_3022 = _EVAL_3442 | _EVAL_2851;
  assign _EVAL_1008 = 9'h9b == _EVAL_1399;
  assign _EVAL_2938 = 9'h10f == _EVAL_1399 ? _EVAL_374 : _EVAL_2086;
  assign _EVAL_788 = 9'h191 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3154;
  assign _EVAL_3337 = _EVAL_3558 & 7'h28;
  assign _EVAL_486 = 9'hdc == _EVAL_1399 ? _EVAL_3000 : _EVAL_2611;
  assign _EVAL_1325 = 9'h162 == _EVAL_1399 ? _EVAL_374 : _EVAL_2489;
  assign _EVAL_179 = 9'h1e4 == _EVAL_1399 ? _EVAL_374 : _EVAL_1140;
  assign _EVAL_2363 = {_EVAL_3116,_EVAL_95,_EVAL_1552,_EVAL_2344};
  assign _EVAL_2512 = 9'h9c == _EVAL_1399 ? 32'h0 : _EVAL_419;
  assign _EVAL_2691 = _EVAL_421 ? 1'h0 : _EVAL_275;
  assign _EVAL_1525 = 9'hbb == _EVAL_1399 ? 32'h0 : _EVAL_239;
  assign _EVAL_541 = 9'h144 == _EVAL_1399 ? _EVAL_374 : _EVAL_1813;
  assign _EVAL_1480 = _EVAL_2774 | _EVAL_585;
  assign _EVAL_2948 = {1'h0,_EVAL_2987,_EVAL_2987,_EVAL_2336,_EVAL_280};
  assign _EVAL_132 = _EVAL_3306 | _EVAL_3022;
  assign _EVAL_2113 = 9'h65 == _EVAL_1399;
  assign _EVAL_113 = _EVAL_3402 & _EVAL_2317;
  assign _EVAL_2456 = 9'h1c4 == _EVAL_1399 ? _EVAL_374 : _EVAL_1779;
  assign _EVAL_3268 = _EVAL_1367 & _EVAL_1380;
  assign _EVAL_3499 = 9'h62 == _EVAL_1399 ? 32'h0 : _EVAL_3071;
  assign _EVAL_2714 = _EVAL_3815 & _EVAL_2836;
  assign _EVAL_815 = 9'hc7 == _EVAL_1399 ? 32'h0 : _EVAL_1530;
  assign _EVAL_723 = 9'h13c == _EVAL_1399 ? _EVAL_374 : _EVAL_3173;
  assign _EVAL_3743 = 9'h15b == _EVAL_1399 ? _EVAL_1856 : _EVAL_2054;
  assign _EVAL_3025 = 9'h116 == _EVAL_1399 ? _EVAL_374 : _EVAL_2812;
  assign _EVAL_563 = _EVAL_3182 & _EVAL_1135;
  assign _EVAL_549 = _EVAL_1589 & _EVAL_234;
  assign _EVAL_2017 = _EVAL_2008 | _EVAL_1045;
  assign _EVAL_3700 = _EVAL_1681 | _EVAL_2075;
  assign _EVAL_480 = 9'h49 == _EVAL_1399;
  assign _EVAL_2956 = 9'h43 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3070;
  assign _EVAL_279 = _EVAL_3775 ? _EVAL_2188 : 1'h1;
  assign _EVAL_2520 = 9'h10c == _EVAL_1399 ? _EVAL_1856 : _EVAL_3569;
  assign _EVAL_2489 = 9'h161 == _EVAL_1399 ? _EVAL_374 : _EVAL_2447;
  assign _EVAL_1073 = 9'h9f == _EVAL_1399 ? 32'h0 : _EVAL_3087;
  assign _EVAL_870 = _EVAL_36[11:2];
  assign _EVAL_964 = 9'h43 == _EVAL_1399 ? 32'h0 : _EVAL_1958;
  assign _EVAL_473 = _EVAL_2864 == 8'hff;
  assign _EVAL_1518 = 9'h1c6 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2695;
  assign _EVAL_963 = 9'h109 == _EVAL_1399 ? _EVAL_374 : _EVAL_2820;
  assign _EVAL_577 = _EVAL_2635 | _EVAL_1860;
  assign _EVAL_2651 = _EVAL_3815 & _EVAL_2081;
  assign _EVAL_2079 = 9'h1fa == _EVAL_1399 ? _EVAL_1856 : _EVAL_2050;
  assign _EVAL_957 = _EVAL_3152[4:0];
  assign _EVAL_3444 = _EVAL_3558[2];
  assign _EVAL_3666 = _EVAL_167[1];
  assign _EVAL_331 = _EVAL_2438 | _EVAL_3807;
  assign _EVAL_2928 = 9'h12c == _EVAL_1399 ? _EVAL_374 : _EVAL_3599;
  assign _EVAL_238 = 9'h19e == _EVAL_1399 ? _EVAL_374 : _EVAL_3270;
  assign _EVAL_2410 = 9'h141 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2090;
  assign _EVAL_3026 = _EVAL_870[6];
  assign _EVAL_2420 = _EVAL_26[7:0];
  assign _EVAL_1181 = _EVAL_2643 & _EVAL_502;
  assign _EVAL_2078 = 9'h5e == _EVAL_1399 ? 32'h0 : _EVAL_1532;
  assign _EVAL_3431 = _EVAL_87 | _EVAL_2885;
  assign _EVAL_2265 = 9'h53 == _EVAL_1399;
  assign _EVAL_102 = _EVAL_2246 ? _EVAL_3682 : _EVAL_2248;
  assign _EVAL_622 = 9'h150 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2497;
  assign _EVAL_2786 = _EVAL_1675 & _EVAL_3836;
  assign _EVAL_2896 = _EVAL_421 & _EVAL_3487;
  assign _EVAL_2879 = _EVAL_1549 | _EVAL_3458;
  assign _EVAL_3461 = 9'h44 == _EVAL_1399;
  assign _EVAL_3701 = _EVAL_3498 & _EVAL_2422;
  assign _EVAL_3704 = 9'hd7 == _EVAL_1399;
  assign _EVAL_1435 = _EVAL_1051 ? {{3'd0}, _EVAL_2487} : _EVAL_527;
  assign _EVAL_3031 = {_EVAL_351,_EVAL_2905,_EVAL_1805,_EVAL_3433};
  assign _EVAL_2945 = 9'h198 == _EVAL_1399 ? _EVAL_374 : _EVAL_353;
  assign _EVAL_3265 = 9'h1bb == _EVAL_1399 ? _EVAL_374 : _EVAL_1598;
  assign _EVAL_234 = _EVAL_1987 == 2'h0;
  assign _EVAL_1528 = _EVAL_3234 | _EVAL_3603;
  assign _EVAL_3148 = 9'h1fe == _EVAL_1399 ? _EVAL_1856 : _EVAL_1944;
  assign _EVAL_1666 = _EVAL_3203 & _EVAL_22;
  assign _EVAL_3668 = 9'h1a1 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2390;
  assign _EVAL_1798 = _EVAL_3653 | _EVAL_479;
  assign _EVAL_2503 = 9'h1a6 == _EVAL_1399 ? _EVAL_374 : _EVAL_3741;
  assign _EVAL_450 = 9'h130 == _EVAL_1399 ? _EVAL_374 : _EVAL_1985;
  assign _EVAL_1592 = {{1'd0}, _EVAL_2948};
  assign _EVAL_910 = {{31'd0}, _EVAL_3105};
  assign _EVAL_2977 = 9'h1e6 == _EVAL_1399 ? _EVAL_374 : _EVAL_3504;
  assign _EVAL_3196 = ~_EVAL_959;
  assign _EVAL_268 = 9'hf8 == _EVAL_1399 ? 32'h0 : _EVAL_270;
  assign _EVAL_606 = 9'h1d8 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2560;
  assign _EVAL_2721 = _EVAL_565 | _EVAL_3633;
  assign _EVAL_1591 = 9'h15 == _EVAL_1399 ? 32'h0 : _EVAL_51;
  assign _EVAL_1571 = 9'h1cf == _EVAL_1399 ? _EVAL_374 : _EVAL_990;
  assign _EVAL_1833 = 9'hf5 == _EVAL_1399;
  assign _EVAL_3135 = 9'h28 == _EVAL_1399;
  assign _EVAL_1815 = _EVAL_3249 | _EVAL_487;
  assign _EVAL_1575 = _EVAL_1771 & _EVAL_3649;
  assign _EVAL_61 = {{14'd0}, _EVAL_2538};
  assign _EVAL_3764 = _EVAL_870[8];
  assign _EVAL_1514 = 9'h1f4 == _EVAL_1399 ? _EVAL_374 : _EVAL_3239;
  assign _EVAL_2248 = _EVAL_3662 ? {{14'd0}, _EVAL_1218} : _EVAL_2274;
  assign _EVAL_1000 = 9'hff == _EVAL_1399 ? 32'h0 : _EVAL_3748;
  assign _EVAL_63 = 9'ha0 == _EVAL_1399 ? 32'h0 : _EVAL_1073;
  assign _EVAL_3068 = 9'h100 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1872;
  assign _EVAL_565 = 9'hbb == _EVAL_1399;
  assign _EVAL_3306 = 9'hb0 == _EVAL_1399;
  assign _EVAL_412 = 9'h107 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1812;
  assign _EVAL_1390 = _EVAL_1983 & _EVAL_3485;
  assign _EVAL_1462 = 9'h96 == _EVAL_1399 ? 32'h0 : _EVAL_702;
  assign _EVAL_1124 = 9'h116 == _EVAL_1399 ? _EVAL_1856 : _EVAL_76;
  assign _EVAL_636 = 9'h189 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1429;
  assign _EVAL_585 = _EVAL_1873 | _EVAL_987;
  assign _EVAL_3020 = _EVAL_934 | _EVAL_3310;
  assign _EVAL_2818 = 9'h94 == _EVAL_1399 ? 32'h0 : _EVAL_1527;
  assign _EVAL_3390 = _EVAL_11[7:0];
  assign _EVAL_1553 = _EVAL_2312 | _EVAL_1606;
  assign _EVAL_958 = {_EVAL_2504,_EVAL_748,_EVAL_3444,_EVAL_3385,_EVAL_368};
  assign _EVAL_1154 = 9'h125 == _EVAL_1399 ? _EVAL_374 : _EVAL_2399;
  assign _EVAL_1175 = 9'h1 == _EVAL_1399 ? _EVAL_3670 : _EVAL_3670;
  assign _EVAL_2143 = 9'h1df == _EVAL_1399 ? _EVAL_374 : _EVAL_3454;
  assign _EVAL_2219 = _EVAL_2974 | _EVAL_1115;
  assign _EVAL_1370 = 9'h34 == _EVAL_1399 ? 32'h0 : _EVAL_2057;
  assign _EVAL_2173 = 9'h90 == _EVAL_1399 ? 32'h0 : _EVAL_751;
  assign _EVAL_3342 = _EVAL_2651 | _EVAL_2571;
  assign _EVAL_3252 = _EVAL_769 | _EVAL_2759;
  assign _EVAL_2041 = 9'ha3 == _EVAL_1399;
  assign _EVAL_2495 = 9'h2b == _EVAL_1399 ? 32'h0 : _EVAL_1219;
  assign _EVAL_8 = _EVAL_34;
  assign _EVAL_333 = _EVAL_3574 | _EVAL_2886;
  assign _EVAL_1799 = 9'h1a9 == _EVAL_1399 ? _EVAL_374 : _EVAL_3179;
  assign _EVAL_1109 = 9'h13a == _EVAL_1399 ? _EVAL_374 : _EVAL_869;
  assign _EVAL_857 = 9'h1dc == _EVAL_1399 ? _EVAL_1856 : _EVAL_774;
  assign _EVAL_908 = 9'h110 == _EVAL_1399 ? _EVAL_374 : _EVAL_2938;
  assign _EVAL_56 = 9'h1e0 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2418;
  assign _EVAL_3249 = _EVAL_3369 | _EVAL_397;
  assign _EVAL_757 = _EVAL_3669 | _EVAL_2121;
  assign _EVAL_2711 = _EVAL_26[15:8];
  assign _EVAL_3011 = 9'h24 == _EVAL_1399;
  assign _EVAL_3813 = 9'h3e == _EVAL_1399;
  assign _EVAL_540 = 9'had == _EVAL_1399 ? 32'h0 : _EVAL_3052;
  assign _EVAL_3318 = 9'h1a == _EVAL_1399 ? 32'h0 : _EVAL_1125;
  assign _EVAL_3541 = _EVAL_1684 | _EVAL_3725;
  assign _EVAL_1665 = _EVAL_3090 | _EVAL_3515;
  assign _EVAL_3595 = 9'h31 == _EVAL_1399;
  assign _EVAL_3247 = _EVAL_392 & _EVAL_1856;
  assign _EVAL_3609 = 9'hf9 == _EVAL_1399;
  assign _EVAL_2517 = 9'hbe == _EVAL_1399 ? 32'h0 : _EVAL_2821;
  assign _EVAL_2698 = _EVAL_2797 | _EVAL_577;
  assign _EVAL_3083 = 9'h1e8 == _EVAL_1399 ? _EVAL_374 : _EVAL_3035;
  assign _EVAL_679 = 9'hc9 == _EVAL_1399;
  assign _EVAL_3065 = _EVAL_38;
  assign _EVAL_1019 = 9'ha4 == _EVAL_1399 ? 32'h0 : _EVAL_1383;
  assign _EVAL_2080 = 9'hdb == _EVAL_1399 ? _EVAL_1856 : _EVAL_1569;
  assign _EVAL_922 = 9'h1cb == _EVAL_1399 ? _EVAL_374 : _EVAL_2870;
  assign _EVAL_3454 = 9'h1de == _EVAL_1399 ? _EVAL_374 : _EVAL_2089;
  assign _EVAL_3555 = _EVAL_2486 | _EVAL_1935;
  assign _EVAL_3520 = 9'h1b7 == _EVAL_1399 ? _EVAL_374 : _EVAL_1170;
  assign _EVAL_2862 = 9'h8b == _EVAL_1399;
  assign _EVAL_1822 = _EVAL_1693 | _EVAL_728;
  assign _EVAL_3814 = _EVAL_1603 | _EVAL_1261;
  assign _EVAL_2777 = 9'h103 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1568;
  assign _EVAL_3549 = 9'h22 == _EVAL_1399 ? 32'h0 : _EVAL_2480;
  assign _EVAL_1746 = 9'h19 == _EVAL_1399;
  assign _EVAL_329 = 9'h19a == _EVAL_1399 ? _EVAL_1856 : _EVAL_1769;
  assign _EVAL_3694 = 9'h71 == _EVAL_1399;
  assign _EVAL_2858 = 9'h12d == _EVAL_1399 ? _EVAL_1856 : _EVAL_3298;
  assign _EVAL_2992 = _EVAL_1362 | _EVAL_1390;
  assign _EVAL_2743 = 512'h1 << _EVAL_1399;
  assign _EVAL_2797 = 9'h69 == _EVAL_1399;
  assign _EVAL_1408 = 9'h1f5 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3233;
  assign _EVAL_244 = 9'hdf == _EVAL_1399 ? _EVAL_1856 : _EVAL_3465;
  assign _EVAL_439 = 9'h46 == _EVAL_1399;
  assign _EVAL_808 = _EVAL_234 ? _EVAL_1206 : _EVAL_3223;
  assign _EVAL_169 = 5'hb == _EVAL_958;
  assign _EVAL_1937 = 9'h1b5 == _EVAL_1399 ? _EVAL_374 : _EVAL_2558;
  assign _EVAL_2210 = 9'h37 == _EVAL_1399 ? 32'h0 : _EVAL_332;
  assign _EVAL_3600 = 9'h1f2 == _EVAL_1399 ? _EVAL_1856 : _EVAL_545;
  assign _EVAL_1221 = 9'h7d == _EVAL_1399 ? 32'h0 : _EVAL_608;
  assign _EVAL_3001 = _EVAL_3246 | _EVAL_951;
  assign _EVAL_2894 = 9'h98 == _EVAL_1399 ? 32'h0 : _EVAL_3542;
  assign _EVAL_2812 = 9'h115 == _EVAL_1399 ? _EVAL_374 : _EVAL_2816;
  assign _EVAL_1830 = _EVAL_3498 & _EVAL_473;
  assign _EVAL_1490 = 9'h131 == _EVAL_1399 ? _EVAL_374 : _EVAL_450;
  assign _EVAL_368 = _EVAL_3558[0];
  assign _EVAL_3829 = _EVAL_28[1];
  assign _EVAL_3661 = 9'h16f == _EVAL_1399 ? _EVAL_374 : _EVAL_2927;
  assign _EVAL_1804 = _EVAL_1752 & _EVAL_3485;
  assign _EVAL_1476 = 9'hc3 == _EVAL_1399;
  assign _EVAL_2895 = 9'h171 == _EVAL_1399 ? _EVAL_374 : _EVAL_2854;
  assign _EVAL_3531 = 9'h1be == _EVAL_1399 ? _EVAL_1856 : _EVAL_2533;
  assign _EVAL_2937 = 9'h1e1 == _EVAL_1399 ? _EVAL_1856 : _EVAL_56;
  assign _EVAL_1557 = _EVAL_1186 | _EVAL_2888;
  assign _EVAL_2021 = _EVAL_2992 | _EVAL_3423;
  assign _EVAL_2836 = _EVAL_1319 == 8'hff;
  assign _EVAL_859 = {6'h0,_EVAL_2978,_EVAL_2218,6'h0,_EVAL_2978,_EVAL_2218,6'h0,_EVAL_2978,_EVAL_2218};
  assign _EVAL_3470 = _EVAL_2883 | _EVAL_2593;
  assign _EVAL_2497 = 9'h14f == _EVAL_1399 ? _EVAL_1856 : _EVAL_785;
  assign _EVAL_2593 = _EVAL_2602 | _EVAL_2569;
  assign _EVAL_3722 = 9'h1fb == _EVAL_1399 ? _EVAL_1856 : _EVAL_2079;
  assign _EVAL_881 = 9'h7f == _EVAL_1399;
  assign _EVAL_3769 = 9'h180 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1790;
  assign _EVAL_3061 = 9'h3b == _EVAL_1399 ? 32'h0 : _EVAL_2755;
  assign _EVAL_2262 = _EVAL_2743[224];
  assign _EVAL_699 = _EVAL_499 | _EVAL_2881;
  assign _EVAL_1897 = _EVAL_83[15];
  assign _EVAL_2207 = 9'h88 == _EVAL_1399;
  assign _EVAL_949 = 9'h1ae == _EVAL_1399 ? _EVAL_374 : _EVAL_3403;
  assign _EVAL_3841 = _EVAL_468 & _EVAL_3485;
  assign _EVAL_3669 = 9'h35 == _EVAL_1399;
  assign _EVAL_2101 = _EVAL_1975 | _EVAL_3470;
  assign _EVAL_3537 = 9'h19e == _EVAL_1399 ? _EVAL_1856 : _EVAL_1659;
  assign _EVAL_2414 = _EVAL_2643 & _EVAL_1368;
  assign _EVAL_1066 = 9'h1ad == _EVAL_1399 ? _EVAL_1856 : _EVAL_2136;
  assign _EVAL_3132 = _EVAL_3663 | _EVAL_996;
  assign _EVAL_45 = _EVAL_1184 & _EVAL_3485;
  assign _EVAL_3783 = _EVAL_2955 | _EVAL_2573;
  assign _EVAL_2887 = _EVAL_1496 | _EVAL_65;
  assign _EVAL_1893 = _EVAL_3813 | _EVAL_2101;
  assign _EVAL_3035 = 9'h1e7 == _EVAL_1399 ? _EVAL_374 : _EVAL_2977;
  assign _EVAL_3366 = _EVAL_1238 | _EVAL_372;
  assign _EVAL_820 = 9'hc == _EVAL_1399 ? 32'h7b202473 : _EVAL_2001;
  assign _EVAL_1888 = _EVAL_1771 & _EVAL_2920;
  assign _EVAL_2616 = 9'hcc == _EVAL_1399 ? 32'h0 : _EVAL_2277;
  assign _EVAL_3427 = _EVAL_876 | _EVAL_753;
  assign _EVAL_2623 = 9'h181 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3769;
  assign _EVAL_1003 = 9'hf4 == _EVAL_1399 ? 32'h0 : _EVAL_2736;
  assign _EVAL_403 = _EVAL_1110 | _EVAL_3535;
  assign _EVAL_2499 = _EVAL_83[14];
  assign _EVAL_2051 = _EVAL_926 & _EVAL_234;
  assign _EVAL_3429 = _EVAL_870[2];
  assign _EVAL_996 = _EVAL_480 | _EVAL_154;
  assign _EVAL_3097 = 9'h1 == _EVAL_1399 ? 32'h380006f : 32'hc0006f;
  assign _EVAL_1206 = _EVAL_1437 ? 1'h0 : _EVAL_1152;
  assign _EVAL_3458 = _EVAL_3567 | _EVAL_1480;
  assign _EVAL_1368 = _EVAL_83[4];
  assign _EVAL_516 = 9'h198 == _EVAL_1399 ? _EVAL_1856 : _EVAL_969;
  assign _EVAL_514 = 9'h114 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2039;
  assign _EVAL_1925 = 9'ha2 == _EVAL_1399 ? 32'h0 : _EVAL_912;
  assign _EVAL_846 = 9'h162 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1258;
  assign _EVAL_3331 = _EVAL_965 | _EVAL_2732;
  assign _EVAL_2457 = 9'h99 == _EVAL_1399 ? 32'h0 : _EVAL_2894;
  assign _EVAL_1856 = _EVAL_306 == 10'h0;
  assign _EVAL_3800 = 9'h1b3 == _EVAL_1399 ? _EVAL_374 : _EVAL_669;
  assign _EVAL_2736 = 9'hf3 == _EVAL_1399 ? 32'h0 : _EVAL_1622;
  assign _EVAL_2770 = 9'h18f == _EVAL_1399 ? _EVAL_374 : _EVAL_2392;
  assign _EVAL_1275 = _EVAL_3795 & _EVAL_3196;
  assign _EVAL_1401 = {17'h7000,_EVAL_2138,_EVAL_957,7'h3};
  assign _EVAL_956 = 9'h1c1 == _EVAL_1399 ? _EVAL_374 : _EVAL_2063;
  assign _EVAL_766 = 9'h1ed == _EVAL_1399 ? _EVAL_374 : _EVAL_567;
  assign _EVAL_1026 = 9'h11 == _EVAL_1399 ? 32'h7b202473 : _EVAL_3017;
  assign _EVAL_1110 = debug_hartReset_0__EVAL_1;
  assign _EVAL_959 = _EVAL_2763 == 8'h0;
  assign _EVAL_1290 = 9'hb7 == _EVAL_1399 ? 32'h0 : _EVAL_2268;
  assign _EVAL_502 = _EVAL_83[0];
  assign _EVAL_1738 = 9'hd8 == _EVAL_1399 ? 32'h0 : _EVAL_3738;
  assign _EVAL_1159 = 9'h195 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3299;
  assign _EVAL_2911 = 9'h4c == _EVAL_1399;
  assign _EVAL_1341 = 9'h1b1 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2595;
  assign _EVAL_2724 = 9'h10 == _EVAL_1399 ? _EVAL_3670 : _EVAL_2120;
  assign _EVAL_3487 = _EVAL_3395 ? 1'h0 : _EVAL_3104;
  assign _EVAL_705 = 9'h63 == _EVAL_1399;
  assign _EVAL_3030 = _EVAL_204 | _EVAL_2145;
  assign _EVAL_306 = _EVAL_870 & 10'h200;
  assign _EVAL_130 = 9'h82 == _EVAL_1399;
  assign _EVAL_1597 = 9'h1af == _EVAL_1399 ? _EVAL_1856 : _EVAL_3745;
  assign _EVAL_2272 = _EVAL_710 & _EVAL_3666;
  assign _EVAL_2522 = _EVAL_2959 | _EVAL_481;
  assign _EVAL_2040 = 9'hd9 == _EVAL_1399;
  assign _EVAL_3403 = 9'h1ad == _EVAL_1399 ? _EVAL_374 : _EVAL_3493;
  assign _EVAL_1672 = 9'hfa == _EVAL_1399 ? 32'h0 : _EVAL_1994;
  assign _EVAL_2096 = 9'h137 == _EVAL_1399 ? _EVAL_374 : _EVAL_2306;
  assign _EVAL_763 = _EVAL_1493 | _EVAL_3235;
  assign _EVAL_317 = _EVAL_2929 | _EVAL_1237;
  assign _EVAL_1487 = 9'hd6 == _EVAL_1399;
  assign _EVAL_759 = _EVAL_1746 | _EVAL_2566;
  assign _EVAL_916 = 9'h128 == _EVAL_1399 ? _EVAL_1856 : _EVAL_180;
  assign _EVAL_2882 = 9'h7f == _EVAL_1399 ? 32'h0 : _EVAL_471;
  assign _EVAL_2809 = 9'h100 == _EVAL_1399 ? _EVAL_374 : _EVAL_1000;
  assign _EVAL_1020 = 9'had == _EVAL_1399;
  assign _EVAL_2627 = _EVAL_2040 | _EVAL_1121;
  assign _EVAL_692 = 9'h123 == _EVAL_1399 ? _EVAL_374 : _EVAL_2850;
  assign _EVAL_2031 = 9'h69 == _EVAL_1399 ? 32'h0 : _EVAL_789;
  assign _EVAL_3372 = 9'hda == _EVAL_1399 ? 32'h0 : _EVAL_2804;
  assign _EVAL_1993 = 9'hca == _EVAL_1399;
  assign _EVAL_2689 = 9'h1ba == _EVAL_1399 ? _EVAL_1856 : _EVAL_459;
  assign _EVAL_3409 = 9'h106 == _EVAL_1399 ? _EVAL_374 : _EVAL_1087;
  assign _EVAL_31 = {{2'd0}, _EVAL_3155};
  assign _EVAL_545 = 9'h1f1 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3189;
  assign _EVAL_1198 = _EVAL_3694 | _EVAL_3496;
  assign _EVAL_2251 = 9'h18b == _EVAL_1399 ? _EVAL_374 : _EVAL_3834;
  assign _EVAL_1258 = 9'h161 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1114;
  assign _EVAL_2308 = 9'h137 == _EVAL_1399 ? _EVAL_1856 : _EVAL_285;
  assign _EVAL_2932 = 9'hc8 == _EVAL_1399 ? 32'h0 : _EVAL_815;
  assign _EVAL_324 = 9'h18d == _EVAL_1399 ? _EVAL_374 : _EVAL_3459;
  assign _EVAL_2247 = 9'h15e == _EVAL_1399 ? _EVAL_374 : _EVAL_1036;
  assign _EVAL_1362 = _EVAL_863 | _EVAL_45;
  assign _EVAL_789 = 9'h68 == _EVAL_1399 ? 32'h0 : _EVAL_2588;
  assign _EVAL_3234 = 9'hc1 == _EVAL_1399;
  assign _EVAL_3005 = 9'h152 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2481;
  assign _EVAL_2360 = 9'h11d == _EVAL_1399 ? _EVAL_374 : _EVAL_3140;
  assign _EVAL_2076 = 9'h112 == _EVAL_1399 ? _EVAL_1856 : _EVAL_206;
  assign _EVAL_2057 = 9'h33 == _EVAL_1399 ? 32'h0 : _EVAL_809;
  assign _EVAL_713 = 9'h18e == _EVAL_1399 ? _EVAL_1856 : _EVAL_3169;
  assign _EVAL_1101 = 9'h1d2 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1953;
  assign _EVAL_1230 = _EVAL_3178 | _EVAL_1116;
  assign _EVAL_1873 = 9'hfa == _EVAL_1399;
  assign _EVAL_1687 = _EVAL_2771 | _EVAL_3039;
  assign _EVAL_2611 = 9'hdb == _EVAL_1399 ? _EVAL_3348 : _EVAL_3372;
  assign _EVAL_849 = 9'h3c == _EVAL_1399 ? 32'h0 : _EVAL_3061;
  assign _EVAL_65 = _EVAL_1426 | _EVAL_3366;
  assign _EVAL_1047 = _EVAL_3755 | _EVAL_2083;
  assign _EVAL_1564 = 9'h86 == _EVAL_1399;
  assign _EVAL_2871 = _EVAL_2472 | _EVAL_1095;
  assign _EVAL_3046 = 9'h15e == _EVAL_1399 ? _EVAL_1856 : _EVAL_3762;
  assign _EVAL_1374 = 9'h110 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1268;
  assign _EVAL_1991 = 9'h1e9 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2116;
  assign _EVAL_1138 = 9'h177 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1758;
  assign _EVAL_2488 = _EVAL_2743[221];
  assign _EVAL_3013 = 9'h102 == _EVAL_1399 ? _EVAL_374 : _EVAL_1104;
  assign _EVAL_3377 = 9'h83 == _EVAL_1399 ? 32'h0 : _EVAL_2125;
  assign _EVAL_1377 = 9'h127 == _EVAL_1399 ? _EVAL_374 : _EVAL_3709;
  assign _EVAL_1367 = _EVAL_1422 & _EVAL_1135;
  assign _EVAL_3069 = _EVAL_2207 | _EVAL_3776;
  assign _EVAL_3815 = _EVAL_1754 & _EVAL_2188;
  assign _EVAL_1496 = 9'h99 == _EVAL_1399;
  assign _EVAL_1365 = 9'ha == _EVAL_1399 ? 32'h147413 : _EVAL_2224;
  assign _EVAL_1921 = 9'h9e == _EVAL_1399;
  assign _EVAL_3146 = 9'h1ff == _EVAL_1399 ? _EVAL_374 : _EVAL_3093;
  assign _EVAL_1803 = 9'h95 == _EVAL_1399;
  assign _EVAL_1436 = 9'h191 == _EVAL_1399 ? _EVAL_374 : _EVAL_2737;
  assign _EVAL_3651 = 9'h22 == _EVAL_1399;
  assign _EVAL_2379 = _EVAL_1867 | _EVAL_1506;
  assign _EVAL_451 = _EVAL_1110 ? 1'h0 : _EVAL_2978;
  assign _EVAL_3650 = 9'hd1 == _EVAL_1399 ? 32'h0 : _EVAL_662;
  assign _EVAL_2986 = 9'h117 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1124;
  assign _EVAL_3326 = 9'h6e == _EVAL_1399 ? 32'h0 : _EVAL_3590;
  assign _EVAL_111 = 9'ha7 == _EVAL_1399 ? 32'h0 : _EVAL_182;
  assign _EVAL_592 = 9'h48 == _EVAL_1399 ? 32'h0 : _EVAL_2730;
  assign _EVAL_3027 = 5'hf == _EVAL_958;
  assign _EVAL_2653 = 9'h49 == _EVAL_1399 ? 32'h0 : _EVAL_592;
  assign _EVAL_1471 = _EVAL_382 & _EVAL_3761;
  assign _EVAL_3653 = 9'he1 == _EVAL_1399;
  assign _EVAL_3753 = 9'h156 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2398;
  assign _EVAL_752 = _EVAL_2246 ? _EVAL_2188 : _EVAL_2156;
  assign _EVAL_2097 = _EVAL_870[7];
  assign _EVAL_2847 = 9'hda == _EVAL_1399;
  assign _EVAL_3321 = 9'h10a == _EVAL_1399 ? _EVAL_374 : _EVAL_963;
  assign _EVAL_2788 = _EVAL_3841 | _EVAL_1804;
  assign _EVAL_110 = 9'h1ea == _EVAL_1399 ? _EVAL_374 : _EVAL_2697;
  assign _EVAL_2056 = _EVAL_2 & _EVAL_41;
  assign _EVAL_985 = _EVAL_3698 | _EVAL_497;
  assign _EVAL_2939 = 9'hbe == _EVAL_1399;
  assign _EVAL_1150 = 9'h17e == _EVAL_1399 ? _EVAL_374 : _EVAL_1243;
  assign _EVAL_272 = _EVAL_3236 | _EVAL_2761;
  assign _EVAL_735 = 9'h1c == _EVAL_1399 ? 32'h0 : _EVAL_1583;
  assign _EVAL_2571 = _EVAL_700 & _EVAL_3649;
  assign _EVAL_1007 = 9'h5a == _EVAL_1399 ? 32'h0 : _EVAL_943;
  assign _EVAL_2706 = 9'h1d9 == _EVAL_1399 ? _EVAL_374 : _EVAL_2095;
  assign _EVAL_3228 = 9'he7 == _EVAL_1399 ? 32'h0 : _EVAL_172;
  assign _EVAL_2120 = 9'hf == _EVAL_1399 ? _EVAL_3670 : _EVAL_1425;
  assign _EVAL_1177 = 9'h7d == _EVAL_1399;
  assign _EVAL_2674 = _EVAL_3129 | _EVAL_757;
  assign _EVAL_139 = _EVAL_200 & _EVAL_234;
  assign _EVAL_1941 = 9'h1f2 == _EVAL_1399 ? _EVAL_374 : _EVAL_2494;
  assign _EVAL_1395 = 9'h1bf == _EVAL_1399 ? _EVAL_374 : _EVAL_3295;
  assign _EVAL_837 = 9'h11a == _EVAL_1399 ? _EVAL_374 : _EVAL_2995;
  assign _EVAL_92 = 9'h16 == _EVAL_1399;
  assign _EVAL_930 = 9'h4b == _EVAL_1399 ? 32'h0 : _EVAL_2216;
  assign _EVAL_1957 = _EVAL_817 | _EVAL_3338;
  assign _EVAL_3404 = 9'h1a4 == _EVAL_1399 ? _EVAL_374 : _EVAL_1200;
  assign _EVAL_566 = 9'hb9 == _EVAL_1399 ? 32'h0 : _EVAL_2378;
  assign _EVAL_2110 = 9'h163 == _EVAL_1399 ? _EVAL_374 : _EVAL_1325;
  assign _EVAL_198 = 9'h157 == _EVAL_1399 ? _EVAL_374 : _EVAL_993;
  assign _EVAL_3064 = 9'h77 == _EVAL_1399 ? 32'h0 : _EVAL_1615;
  assign _EVAL_792 = _EVAL_2629 | _EVAL_1835;
  assign _EVAL_3411 = 9'h46 == _EVAL_1399 ? 32'h0 : _EVAL_2249;
  assign _EVAL_2419 = _EVAL_384 | _EVAL_3132;
  assign _EVAL_2437 = _EVAL_624 & _EVAL_3221;
  assign _EVAL_172 = 9'he6 == _EVAL_1399 ? 32'h0 : _EVAL_3021;
  assign _EVAL_1186 = 9'h90 == _EVAL_1399;
  assign _EVAL_2185 = _EVAL_3426 ? _EVAL_1135 : _EVAL_752;
  assign _EVAL_90 = _EVAL_619 | _EVAL_1528;
  assign _EVAL_1659 = 9'h19d == _EVAL_1399 ? _EVAL_1856 : _EVAL_906;
  assign _EVAL_347 = _EVAL_1240 | _EVAL_2256;
  assign _EVAL_3750 = _EVAL_2363[15:8];
  assign _EVAL_2052 = 9'h44 == _EVAL_1399 ? 32'h0 : _EVAL_964;
  assign _EVAL_3515 = _EVAL_3461 | _EVAL_2956;
  assign _EVAL_2128 = 9'h9 == _EVAL_1399 ? _EVAL_3670 : _EVAL_2831;
  assign _EVAL_3513 = 9'h103 == _EVAL_1399 ? _EVAL_374 : _EVAL_3013;
  assign _EVAL_2024 = 9'h15c == _EVAL_1399 ? _EVAL_374 : _EVAL_2286;
  assign _EVAL_1448 = _EVAL_28[2];
  assign _EVAL_3644 = 9'h38 == _EVAL_1399 ? 32'h0 : _EVAL_2210;
  assign _EVAL_3490 = 9'h76 == _EVAL_1399;
  assign _EVAL_1838 = 9'hd3 == _EVAL_1399;
  assign _EVAL_3472 = _EVAL_645 | _EVAL_2272;
  assign _EVAL_2885 = _EVAL_2373 | _EVAL_1911;
  assign _EVAL_3140 = 9'h11c == _EVAL_1399 ? _EVAL_374 : _EVAL_1823;
  assign _EVAL_571 = 9'h147 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3711;
  assign _EVAL_1821 = 9'h170 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1014;
  assign _EVAL_76 = 9'h115 == _EVAL_1399 ? _EVAL_1856 : _EVAL_514;
  assign _EVAL_1211 = _EVAL_870[5];
  assign _EVAL_558 = 9'h67 == _EVAL_1399;
  assign _EVAL_3508 = 9'h149 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3408;
  assign _EVAL_2804 = 9'hd9 == _EVAL_1399 ? 32'h0 : _EVAL_1738;
  assign _EVAL_2699 = 9'h152 == _EVAL_1399 ? _EVAL_374 : _EVAL_1012;
  assign _EVAL_601 = 9'h1dc == _EVAL_1399 ? _EVAL_374 : _EVAL_1658;
  assign _EVAL_2081 = _EVAL_2727 == 8'hff;
  assign _EVAL_3509 = _EVAL_2437 & _EVAL_3452;
  assign _EVAL_1590 = _EVAL_1082 & _EVAL_659;
  assign _EVAL_118 = 9'hfd == _EVAL_1399 ? 32'h0 : _EVAL_1350;
  assign _EVAL_402 = 9'h1c2 == _EVAL_1399 ? _EVAL_1856 : _EVAL_890;
  assign _EVAL_230 = _EVAL_3207[16];
  assign _EVAL_1450 = 9'h130 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2878;
  assign _EVAL_1319 = _EVAL_575[15:8];
  assign _EVAL_1807 = 9'h1d4 == _EVAL_1399 ? _EVAL_374 : _EVAL_2476;
  assign _EVAL_2063 = 9'h1c0 == _EVAL_1399 ? _EVAL_374 : _EVAL_1395;
  assign _EVAL_3568 = 9'h1ab == _EVAL_1399 ? _EVAL_1856 : _EVAL_2853;
  assign _EVAL_3244 = _EVAL_26[31:24];
  assign _EVAL_1883 = _EVAL_3750 == 8'hff;
  assign _EVAL_1231 = _EVAL_1993 | _EVAL_3096;
  assign _EVAL_2285 = 9'h1a == _EVAL_1399;
  assign _EVAL_1422 = _EVAL_2643 & _EVAL_2104;
  assign _EVAL_1725 = 9'h1c5 == _EVAL_1399 ? _EVAL_374 : _EVAL_2456;
  assign _EVAL_3212 = _EVAL_2964 | _EVAL_3530;
  assign _EVAL_3145 = 9'h88 == _EVAL_1399 ? 32'h0 : _EVAL_2223;
  assign _EVAL_3271 = 9'h112 == _EVAL_1399 ? _EVAL_374 : _EVAL_1478;
  assign _EVAL_1036 = 9'h15d == _EVAL_1399 ? _EVAL_374 : _EVAL_2024;
  assign _EVAL_3687 = 9'h1d6 == _EVAL_1399 ? _EVAL_374 : _EVAL_1982;
  assign _EVAL_2163 = _EVAL_3207[15:0];
  assign _EVAL_1332 = _EVAL_2279 | _EVAL_2366;
  assign _EVAL_2820 = 9'h108 == _EVAL_1399 ? _EVAL_374 : _EVAL_308;
  assign _EVAL_1658 = 9'h1db == _EVAL_1399 ? _EVAL_374 : _EVAL_1324;
  assign _EVAL_817 = 9'h84 == _EVAL_1399;
  assign _EVAL_401 = 9'h1c9 == _EVAL_1399 ? _EVAL_1856 : _EVAL_97;
  assign _EVAL_1834 = _EVAL_700 & _EVAL_2920;
  assign _EVAL_1360 = _EVAL_1182 | _EVAL_347;
  assign _EVAL_3219 = 9'h2 == _EVAL_1399 ? 32'h440006f : _EVAL_3097;
  assign _EVAL_229 = 9'h7 == _EVAL_1399 ? _EVAL_3670 : _EVAL_313;
  assign _EVAL_3774 = 9'ha5 == _EVAL_1399 ? 32'h0 : _EVAL_1019;
  assign _EVAL_2403 = _EVAL_3393 | _EVAL_2325;
  assign _EVAL_3259 = _EVAL_2237 | _EVAL_1646;
  assign _EVAL_3647 = 9'h199 == _EVAL_1399 ? _EVAL_374 : _EVAL_2945;
  assign _EVAL_16 = _EVAL_3066;
  assign _EVAL_1699 = _EVAL_28[3];
  assign _EVAL_685 = 9'h8a == _EVAL_1399;
  assign _EVAL_3539 = 9'h19a == _EVAL_1399 ? _EVAL_374 : _EVAL_3647;
  assign _EVAL_2881 = _EVAL_3490 | _EVAL_3838;
  assign _EVAL_2482 = 9'h78 == _EVAL_1399 ? 32'h0 : _EVAL_3064;
  assign _EVAL_2279 = 9'h4f == _EVAL_1399;
  assign _EVAL_3102 = _EVAL_11[31:24];
  assign _EVAL_3727 = 9'h133 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3576;
  assign _EVAL_942 = 9'haf == _EVAL_1399 ? 32'h0 : _EVAL_3288;
  assign _EVAL_1155 = _EVAL_3731 & _EVAL_3395;
  assign _EVAL_1127 = 9'h25 == _EVAL_1399;
  assign _EVAL_829 = _EVAL_3782 & _EVAL_2422;
  assign _EVAL_2445 = ~_EVAL_2978;
  assign _EVAL_3784 = _EVAL_1931 | _EVAL_851;
  assign _EVAL_1540 = _EVAL_2651 & _EVAL_234;
  assign _EVAL_2578 = 9'h187 == _EVAL_1399 ? _EVAL_374 : _EVAL_3506;
  assign _EVAL_1839 = 9'h8c == _EVAL_1399;
  assign _EVAL_3442 = 9'haf == _EVAL_1399;
  assign _EVAL_2886 = _EVAL_736 | _EVAL_3144;
  assign _EVAL_1723 = 9'he0 == _EVAL_1399 ? _EVAL_3682 : _EVAL_1697;
  assign _EVAL_2092 = 9'h5e == _EVAL_1399;
  assign _EVAL_2418 = 9'h1df == _EVAL_1399 ? _EVAL_1856 : _EVAL_219;
  assign _EVAL_3566 = 9'h51 == _EVAL_1399 ? 32'h0 : _EVAL_191;
  assign _EVAL_2774 = 9'hfb == _EVAL_1399;
  assign _EVAL_2641 = _EVAL_2532 | _EVAL_132;
  assign _EVAL_1977 = 9'h183 == _EVAL_1399 ? _EVAL_374 : _EVAL_931;
  assign _EVAL_127 = 9'h16a == _EVAL_1399 ? _EVAL_374 : _EVAL_1269;
  assign _EVAL_2254 = _EVAL_1339 & 12'h1;
  assign _EVAL_3239 = 9'h1f3 == _EVAL_1399 ? _EVAL_374 : _EVAL_1941;
  assign _EVAL_2538 = _EVAL_11[17:16];
  assign _EVAL_1693 = 9'hac == _EVAL_1399;
  assign _EVAL_2177 = 9'h1a9 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1517;
  assign _EVAL_2861 = _EVAL_2012 & _EVAL_181;
  assign _EVAL_1035 = 9'h15 == _EVAL_1399;
  assign _EVAL_1494 = 9'h192 == _EVAL_1399 ? _EVAL_1856 : _EVAL_788;
  assign _EVAL_3791 = _EVAL_3775 ? _EVAL_910 : 32'h0;
  assign _EVAL_1754 = _EVAL_1675 & _EVAL_1368;
  assign _EVAL_3663 = 9'h4a == _EVAL_1399;
  assign _EVAL_2255 = 9'h53 == _EVAL_1399 ? 32'h0 : _EVAL_2829;
  assign _EVAL_835 = 9'h1a0 == _EVAL_1399 ? _EVAL_374 : _EVAL_3421;
  assign _EVAL_1620 = _EVAL_29[2];
  assign _EVAL_719 = 9'h41 == _EVAL_1399 ? _EVAL_1856 : _EVAL_822;
  assign _EVAL_1307 = 9'h13f == _EVAL_1399 ? _EVAL_1856 : _EVAL_3689;
  assign _EVAL_1170 = 9'h1b6 == _EVAL_1399 ? _EVAL_374 : _EVAL_1937;
  assign _EVAL_2486 = 9'he6 == _EVAL_1399;
  assign _EVAL_526 = _EVAL_2731 | _EVAL_375;
  assign _EVAL_1160 = 9'h19f == _EVAL_1399 ? _EVAL_1856 : _EVAL_3537;
  assign _EVAL_219 = 9'h1de == _EVAL_1399 ? _EVAL_1856 : _EVAL_3736;
  assign _EVAL_2688 = 9'ha8 == _EVAL_1399;
  assign _EVAL_3103 = 9'h1b6 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3714;
  assign _EVAL_2326 = 9'hbc == _EVAL_1399 ? 32'h0 : _EVAL_1525;
  assign _EVAL_1098 = 9'h1b4 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1936;
  assign _EVAL_3676 = 9'h28 == _EVAL_1399 ? 32'h0 : _EVAL_3387;
  assign _EVAL_2851 = _EVAL_1734 | _EVAL_1599;
  assign _EVAL_459 = 9'h1b9 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1486;
  assign _EVAL_1271 = _EVAL_870[1];
  assign _EVAL_1669 = _EVAL_3595 | _EVAL_3259;
  assign _EVAL_131 = 9'h166 == _EVAL_1399 ? _EVAL_1856 : _EVAL_847;
  assign _EVAL_1081 = 9'h1a6 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2712;
  assign _EVAL_1420 = 9'ha == _EVAL_1399 ? _EVAL_3670 : _EVAL_2128;
  assign _EVAL_366 = _EVAL_2828 & _EVAL_234;
  assign _EVAL_2781 = 9'hdd == _EVAL_1399 ? _EVAL_1856 : _EVAL_3606;
  assign _EVAL_1547 = 9'h18 == _EVAL_1399 ? 32'h0 : _EVAL_1853;
  assign _EVAL_2395 = _EVAL_881 | _EVAL_3746;
  assign _EVAL_312 = 9'h71 == _EVAL_1399 ? 32'h0 : _EVAL_882;
  assign _EVAL_124 = _EVAL_506 | _EVAL_886;
  assign _EVAL_2174 = 9'h85 == _EVAL_1399;
  assign _EVAL_1720 = 9'h4e == _EVAL_1399;
  assign _EVAL_2687 = 9'h8b == _EVAL_1399 ? 32'h0 : _EVAL_3073;
  assign _EVAL_3530 = _EVAL_2113 | _EVAL_343;
  assign _EVAL_1257 = 9'h148 == _EVAL_1399 ? _EVAL_374 : _EVAL_1633;
  assign _EVAL_2115 = _EVAL_3388 | _EVAL_3069;
  assign _EVAL_382 = _EVAL_3795 & _EVAL_959;
  assign _EVAL_2791 = 9'hf6 == _EVAL_1399 ? 32'h0 : _EVAL_325;
  assign _EVAL_1567 = 9'h1c == _EVAL_1399;
  assign _EVAL_2700 = 9'heb == _EVAL_1399;
  assign _EVAL_2837 = 9'h1cb == _EVAL_1399 ? _EVAL_1856 : _EVAL_1742;
  assign _EVAL_1835 = _EVAL_1034 | _EVAL_1047;
  assign _EVAL_3776 = _EVAL_150 | _EVAL_3751;
  assign _EVAL_187 = 9'h1e4 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3171;
  assign _EVAL_49 = 9'he1 == _EVAL_1399 ? 32'h0 : _EVAL_1723;
  assign _EVAL_744 = 9'h1bc == _EVAL_1399 ? _EVAL_1856 : _EVAL_3323;
  assign _EVAL_3195 = 9'hc8 == _EVAL_1399;
  assign _EVAL_1429 = 9'h188 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3475;
  assign _EVAL_181 = ~_EVAL_2624;
  assign _EVAL_2695 = 9'h1c5 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3128;
  assign _EVAL_3281 = 9'h2e == _EVAL_1399;
  assign _EVAL_2504 = _EVAL_3558[6];
  assign _EVAL_771 = 9'h12a == _EVAL_1399 ? _EVAL_1856 : _EVAL_2220;
  assign _EVAL_3577 = _EVAL_1099 | _EVAL_3331;
  assign _EVAL_2306 = 9'h136 == _EVAL_1399 ? _EVAL_374 : _EVAL_327;
  assign _EVAL_2312 = 9'ha7 == _EVAL_1399;
  assign _EVAL_3169 = 9'h18d == _EVAL_1399 ? _EVAL_1856 : _EVAL_3217;
  assign _EVAL_1795 = 9'hec == _EVAL_1399 ? 32'h0 : _EVAL_2432;
  assign _EVAL_1220 = _EVAL_1476 | _EVAL_90;
  assign _EVAL_1276 = 9'h64 == _EVAL_1399 ? 32'h0 : _EVAL_258;
  assign _EVAL_1139 = 9'h5c == _EVAL_1399 ? 32'h0 : _EVAL_3200;
  assign _EVAL_2224 = 9'h9 == _EVAL_1399 ? 32'hfe0408e3 : _EVAL_2908;
  assign _EVAL_2712 = 9'h1a5 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2074;
  assign _EVAL_900 = 9'h169 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2073;
  assign _EVAL_95 = _EVAL_1448 ? 8'hff : 8'h0;
  assign _EVAL_608 = 9'h7c == _EVAL_1399 ? 32'h0 : _EVAL_123;
  assign _EVAL_3502 = 9'hce == _EVAL_1399;
  assign _EVAL_488 = 9'h1f == _EVAL_1399;
  assign _EVAL_1936 = 9'h1b3 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2162;
  assign _EVAL_1375 = 9'h6a == _EVAL_1399;
  assign _EVAL_832 = _EVAL_1487 | _EVAL_370;
  assign _EVAL_3094 = 9'h32 == _EVAL_1399;
  assign _EVAL_1399 = {_EVAL_3764,_EVAL_2097,_EVAL_3026,_EVAL_1211,_EVAL_2387,_EVAL_725,_EVAL_3429,_EVAL_1271,_EVAL_842};
  assign _EVAL_2378 = 9'hb8 == _EVAL_1399 ? 32'h0 : _EVAL_1290;
  assign _EVAL_921 = 9'he5 == _EVAL_1399;
  assign _EVAL_323 = 9'hbc == _EVAL_1399;
  assign _EVAL_2237 = 9'h30 == _EVAL_1399;
  assign _EVAL_339 = 9'h164 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1038;
  assign _EVAL_3641 = _EVAL_1841 | _EVAL_271;
  assign _EVAL_882 = 9'h70 == _EVAL_1399 ? 32'h0 : _EVAL_1285;
  assign _EVAL_1572 = 9'hea == _EVAL_1399;
  assign _EVAL_3436 = _EVAL_2988 | _EVAL_360;
  assign _EVAL_997 = _EVAL_3731 & _EVAL_2840;
  assign _EVAL_2324 = _EVAL_11[0];
  assign _EVAL_3825 = 9'he9 == _EVAL_1399;
  assign _EVAL_802 = _EVAL_1701 | _EVAL_697;
  assign _EVAL_1896 = _EVAL_968 | _EVAL_2522;
  assign _EVAL_2527 = 9'h8d == _EVAL_1399;
  assign _EVAL_2334 = 9'h188 == _EVAL_1399 ? _EVAL_374 : _EVAL_2578;
  assign _EVAL_1985 = 9'h12f == _EVAL_1399 ? _EVAL_374 : _EVAL_78;
  assign _EVAL_71 = 9'h15c == _EVAL_1399 ? _EVAL_1856 : _EVAL_3743;
  assign _EVAL_1512 = _EVAL_2092 | _EVAL_1230;
  assign _EVAL_3457 = 9'h6b == _EVAL_1399;
  assign _EVAL_327 = 9'h135 == _EVAL_1399 ? _EVAL_374 : _EVAL_432;
  assign _EVAL_760 = _EVAL_2970 | _EVAL_3290;
  assign _EVAL_2934 = 9'h141 == _EVAL_1399 ? _EVAL_374 : _EVAL_3059;
  assign _EVAL_799 = 9'h89 == _EVAL_1399 ? 32'h0 : _EVAL_3145;
  assign _EVAL_2233 = 9'h145 == _EVAL_1399 ? _EVAL_374 : _EVAL_541;
  assign _EVAL_3448 = _EVAL_2843 | _EVAL_833;
  assign _EVAL_1475 = _EVAL_2437 & _EVAL_638;
  assign _EVAL_2005 = _EVAL_1194 | _EVAL_3342;
  assign _EVAL_3551 = 9'h5c == _EVAL_1399;
  assign _EVAL_251 = 9'h173 == _EVAL_1399 ? _EVAL_374 : _EVAL_960;
  assign _EVAL_3328 = _EVAL_1433 | _EVAL_2524;
  assign _EVAL_3127 = _EVAL_3195 | _EVAL_792;
  assign _EVAL_1507 = 9'h120 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3325;
  assign _EVAL_2842 = 9'h3f == _EVAL_1399 ? 32'h0 : _EVAL_2384;
  assign _EVAL_1423 = _EVAL_3094 | _EVAL_1669;
  assign _EVAL_1104 = 9'h101 == _EVAL_1399 ? _EVAL_374 : _EVAL_2809;
  assign _EVAL_1147 = 9'h16b == _EVAL_1399 ? _EVAL_374 : _EVAL_127;
  assign _EVAL_2995 = 9'h119 == _EVAL_1399 ? _EVAL_374 : _EVAL_3739;
  assign _EVAL_378 = 9'h1cd == _EVAL_1399 ? _EVAL_1856 : _EVAL_2758;
  assign _EVAL_1049 = _EVAL_3782 & _EVAL_473;
  assign _EVAL_2771 = 9'h5b == _EVAL_1399;
  assign _EVAL_2915 = 9'he9 == _EVAL_1399 ? 32'h0 : _EVAL_3095;
  assign _EVAL_2619 = 9'ha8 == _EVAL_1399 ? 32'h0 : _EVAL_111;
  assign _EVAL_2870 = 9'h1ca == _EVAL_1399 ? _EVAL_374 : _EVAL_630;
  assign _EVAL_1167 = 9'hd2 == _EVAL_1399 ? 32'h0 : _EVAL_3650;
  assign _EVAL_374 = {6'h0,_EVAL_2978,_EVAL_2218,_EVAL_859};
  assign _EVAL_1736 = 9'hb5 == _EVAL_1399 ? 32'h0 : _EVAL_143;
  assign _EVAL_3408 = 9'h148 == _EVAL_1399 ? _EVAL_1856 : _EVAL_571;
  assign _EVAL_1935 = _EVAL_921 | _EVAL_2017;
  assign _EVAL_2807 = _EVAL_2411 & _EVAL_2188;
  assign _EVAL_1677 = 9'hc0 == _EVAL_1399 ? 32'h6c0006f : _EVAL_1312;
  assign _EVAL_2039 = 9'h113 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2076;
  assign _EVAL_406 = _EVAL_1631 & _EVAL_1841;
  assign _EVAL_941 = _EVAL_1838 | _EVAL_3009;
  assign _EVAL_2160 = 9'h41 == _EVAL_1399 ? 32'h0 : _EVAL_3359;
  assign _EVAL_762 = 9'h23 == _EVAL_1399;
  assign _EVAL_651 = _EVAL_2491 | _EVAL_3119;
  assign _EVAL_1682 = _EVAL_2363[9:0];
  assign _EVAL_730 = 9'h108 == _EVAL_1399 ? _EVAL_1856 : _EVAL_412;
  assign _EVAL_842 = _EVAL_870[0];
  assign _EVAL_512 = _EVAL_209 | _EVAL_1834;
  assign _EVAL_125 = 9'h149 == _EVAL_1399 ? _EVAL_374 : _EVAL_1257;
  assign _EVAL_485 = 9'h1d7 == _EVAL_1399 ? _EVAL_374 : _EVAL_3687;
  assign _EVAL_3614 = _EVAL_734 & _EVAL_3177;
  assign _EVAL_946 = 9'h30 == _EVAL_1399 ? 32'h0 : _EVAL_3276;
  assign _EVAL_527 = _EVAL_3027 ? _EVAL_3207 : _EVAL_3791;
  assign _EVAL_2343 = _EVAL_3047 | _EVAL_2683;
  assign _EVAL_2615 = 9'h1d2 == _EVAL_1399 ? _EVAL_374 : _EVAL_1196;
  assign _EVAL_1527 = 9'h93 == _EVAL_1399 ? 32'h0 : _EVAL_2544;
  assign _EVAL_236 = _EVAL_3011 | _EVAL_3511;
  assign _EVAL_697 = _EVAL_3135 | _EVAL_1789;
  assign _EVAL_1992 = 9'hcf == _EVAL_1399 ? 32'h0 : _EVAL_311;
  assign _EVAL_2220 = 9'h129 == _EVAL_1399 ? _EVAL_1856 : _EVAL_916;
  assign _EVAL_3736 = 9'h1dd == _EVAL_1399 ? _EVAL_1856 : _EVAL_857;
  assign _EVAL_3387 = 9'h27 == _EVAL_1399 ? 32'h0 : _EVAL_3067;
  assign _EVAL_2074 = 9'h1a4 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3832;
  assign _EVAL_2558 = 9'h1b4 == _EVAL_1399 ? _EVAL_374 : _EVAL_3800;
  assign _EVAL_2268 = 9'hb6 == _EVAL_1399 ? 32'h0 : _EVAL_1736;
  assign _EVAL_1132 = _EVAL_2862 | _EVAL_505;
  assign _EVAL_2501 = _EVAL_2688 | _EVAL_1553;
  assign _EVAL_2811 = 9'h145 == _EVAL_1399 ? _EVAL_1856 : _EVAL_711;
  assign _EVAL_1710 = _EVAL_3426 ? _EVAL_1576 : _EVAL_102;
  assign _EVAL_1311 = 9'h183 == _EVAL_1399 ? _EVAL_1856 : _EVAL_498;
  assign _EVAL_3832 = 9'h1a3 == _EVAL_1399 ? _EVAL_1856 : _EVAL_98;
  assign _EVAL_2412 = _EVAL_448 | _EVAL_1231;
  assign _EVAL_223 = 9'h4f == _EVAL_1399 ? 32'h0 : _EVAL_175;
  assign _EVAL_3839 = 9'h196 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1159;
  assign _EVAL_751 = 9'h8f == _EVAL_1399 ? 32'h0 : _EVAL_1244;
  assign _EVAL_649 = _EVAL_407 | _EVAL_1893;
  assign _EVAL_739 = 9'h125 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1891;
  assign _EVAL_611 = 9'h56 == _EVAL_1399 ? 32'h0 : _EVAL_3193;
  assign _EVAL_3496 = _EVAL_1989 | _EVAL_331;
  assign _EVAL_3329 = 9'h15f == _EVAL_1399 ? _EVAL_374 : _EVAL_2247;
  assign _EVAL_987 = _EVAL_3609 | _EVAL_3577;
  assign _EVAL_2246 = 5'h4 == _EVAL_958;
  assign _EVAL_2822 = _EVAL_29[3];
  assign _EVAL_1790 = 9'h17f == _EVAL_1399 ? _EVAL_1856 : _EVAL_721;
  assign _EVAL_1812 = 9'h106 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1544;
  assign _EVAL_2684 = 9'h101 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3068;
  assign _EVAL_3498 = _EVAL_1884 & _EVAL_1856;
  assign _EVAL_2789 = 9'h58 == _EVAL_1399 ? 32'h0 : _EVAL_1968;
  assign _EVAL_1513 = 9'hfb == _EVAL_1399 ? 32'h0 : _EVAL_1672;
  assign _EVAL_256 = 9'h164 == _EVAL_1399 ? _EVAL_374 : _EVAL_2110;
  assign _EVAL_1806 = 9'h14b == _EVAL_1399 ? _EVAL_374 : _EVAL_3157;
  assign _EVAL_3703 = 9'hc4 == _EVAL_1399 ? 32'h0 : _EVAL_54;
  assign _EVAL_184 = 9'h155 == _EVAL_1399 ? _EVAL_374 : _EVAL_2351;
  assign _EVAL_2390 = 9'h1a0 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1160;
  assign _EVAL_3634 = 9'h18 == _EVAL_1399;
  assign _EVAL_3325 = 9'h11f == _EVAL_1399 ? _EVAL_1856 : _EVAL_3456;
  assign _EVAL_1228 = _EVAL_2840 & _EVAL_3614;
  assign _EVAL_990 = 9'h1ce == _EVAL_1399 ? _EVAL_374 : _EVAL_1030;
  assign _EVAL_1561 = 9'h19b == _EVAL_1399 ? _EVAL_1856 : _EVAL_329;
  assign _EVAL_1905 = {1'h0,_EVAL_1358,1'h0,_EVAL_2012,8'h1};
  assign _EVAL_1869 = _EVAL_2018 & _EVAL_234;
  assign _EVAL_1734 = 9'hae == _EVAL_1399;
  assign _EVAL_2284 = 9'h1a2 == _EVAL_1399 ? _EVAL_374 : _EVAL_377;
  assign _EVAL_3739 = 9'h118 == _EVAL_1399 ? _EVAL_374 : _EVAL_1297;
  assign _EVAL_392 = _EVAL_2437 & _EVAL_1824;
  assign _EVAL_1633 = 9'h147 == _EVAL_1399 ? _EVAL_374 : _EVAL_1774;
  assign _EVAL_1939 = _EVAL_2347 & _EVAL_2188;
  assign _EVAL_3569 = 9'h10b == _EVAL_1399 ? _EVAL_1856 : _EVAL_1965;
  assign _EVAL_282 = {{10'd0}, _EVAL_1905};
  assign _EVAL_2314 = 9'h80 == _EVAL_1399 ? 32'h0 : _EVAL_2882;
  assign _EVAL_1052 = _EVAL_3209 | _EVAL_2379;
  assign _EVAL_2496 = 9'h2e == _EVAL_1399 ? 32'h0 : _EVAL_3220;
  assign _EVAL_3588 = _EVAL_464 & _EVAL_215;
  assign _EVAL_1900 = 9'h75 == _EVAL_1399 ? 32'h0 : _EVAL_249;
  assign _EVAL_2318 = 9'h12b == _EVAL_1399 ? _EVAL_1856 : _EVAL_771;
  assign _EVAL_3176 = 9'h16a == _EVAL_1399 ? _EVAL_1856 : _EVAL_900;
  assign _EVAL_499 = 9'h77 == _EVAL_1399;
  assign _EVAL_3542 = 9'h97 == _EVAL_1399 ? 32'h0 : _EVAL_1462;
  assign _EVAL_1646 = _EVAL_3816 | _EVAL_1274;
  assign _EVAL_2683 = _EVAL_323 | _EVAL_2721;
  assign _EVAL_3711 = 9'h146 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2811;
  assign _EVAL_2594 = _EVAL_1367 & _EVAL_2920;
  assign _EVAL_389 = 9'h1d3 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1101;
  assign _EVAL_492 = 9'h4 == _EVAL_1399 ? 32'h7b241073 : _EVAL_66;
  assign _EVAL_228 = 9'h1fb == _EVAL_1399 ? _EVAL_374 : _EVAL_2106;
  assign _EVAL_2741 = 9'h11 == _EVAL_1399 ? _EVAL_3670 : _EVAL_2724;
  assign _EVAL_1881 = _EVAL_2845 & _EVAL_234;
  assign _EVAL_37 = _EVAL_2;
  assign _EVAL_2400 = _EVAL_1467 & _EVAL_2819;
  assign _EVAL_1185 = _EVAL_2673 | _EVAL_304;
  assign _EVAL_2366 = _EVAL_1720 | _EVAL_3481;
  assign _EVAL_2451 = 9'h64 == _EVAL_1399;
  assign _EVAL_2077 = 9'h1bf == _EVAL_1399 ? _EVAL_1856 : _EVAL_3531;
  assign _EVAL_650 = _EVAL_3509 & _EVAL_1856;
  assign _EVAL_377 = 9'h1a1 == _EVAL_1399 ? _EVAL_374 : _EVAL_835;
  assign _EVAL_1166 = 9'hba == _EVAL_1399;
  assign _EVAL_2373 = 9'hef == _EVAL_1399;
  assign _EVAL_1545 = 9'hcd == _EVAL_1399 ? 32'h0 : _EVAL_2616;
  assign _EVAL_3672 = 9'hb6 == _EVAL_1399;
  assign _EVAL_1914 = _EVAL_3066 & _EVAL_3177;
  assign _EVAL_1183 = _EVAL_563 & _EVAL_2836;
  assign _EVAL_1383 = 9'ha3 == _EVAL_1399 ? 32'h0 : _EVAL_1925;
  assign _EVAL_436 = 9'hea == _EVAL_1399 ? 32'h0 : _EVAL_2915;
  assign _EVAL_599 = _EVAL_1815 | _EVAL_572;
  assign _EVAL_1846 = _EVAL_1675 & _EVAL_2104;
  assign _EVAL_2989 = 9'h1b1 == _EVAL_1399 ? _EVAL_374 : _EVAL_1096;
  assign _EVAL_2086 = 9'h10e == _EVAL_1399 ? _EVAL_374 : _EVAL_967;
  assign _EVAL_2317 = _EVAL_1110 | _EVAL_1914;
  assign _EVAL_765 = 9'h25 == _EVAL_1399 ? 32'h0 : _EVAL_1366;
  assign _EVAL_174 = 9'h96 == _EVAL_1399;
  assign _EVAL_3518 = {1'h0,_EVAL_3610};
  assign _EVAL_1731 = 9'h14d == _EVAL_1399 ? _EVAL_374 : _EVAL_1613;
  assign _EVAL_484 = 9'h193 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1494;
  assign _EVAL_1972 = 9'hb4 == _EVAL_1399;
  assign _EVAL_2850 = 9'h122 == _EVAL_1399 ? _EVAL_374 : _EVAL_891;
  assign _EVAL_1099 = 9'hf8 == _EVAL_1399;
  assign _EVAL_3087 = 9'h9e == _EVAL_1399 ? 32'h0 : _EVAL_3320;
  assign _EVAL_2565 = 9'h14b == _EVAL_1399 ? _EVAL_1856 : _EVAL_3612;
  assign _EVAL_1151 = _EVAL_3474 == 8'hff;
  assign _EVAL_3160 = _EVAL_1176 ? _EVAL_2188 : _EVAL_420;
  assign _EVAL_3742 = 9'h50 == _EVAL_1399;
  assign _EVAL_575 = {_EVAL_3770,_EVAL_530,_EVAL_2280,_EVAL_991};
  assign _EVAL_1767 = 9'h173 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1445;
  assign _EVAL_1324 = 9'h1da == _EVAL_1399 ? _EVAL_374 : _EVAL_2706;
  assign _EVAL_3090 = 9'h45 == _EVAL_1399;
  assign _EVAL_1004 = 9'hde == _EVAL_1399 ? _EVAL_1576 : _EVAL_972;
  assign _EVAL_995 = _EVAL_1184 ? _EVAL_11 : 32'h0;
  assign _EVAL_1556 = 9'h23 == _EVAL_1399 ? 32'h0 : _EVAL_3549;
  assign _EVAL_1523 = _EVAL_650 & _EVAL_2819;
  assign _EVAL_1928 = _EVAL_1035 | _EVAL_2642;
  assign _EVAL_2959 = 9'h51 == _EVAL_1399;
  assign _EVAL_206 = 9'h111 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1374;
  assign _EVAL_3593 = 9'h9d == _EVAL_1399;
  assign _EVAL_325 = 9'hf5 == _EVAL_1399 ? 32'h0 : _EVAL_1003;
  assign _EVAL_3246 = 9'hb8 == _EVAL_1399;
  assign _EVAL_934 = 9'haa == _EVAL_1399;
  assign _EVAL_3251 = 9'h142 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2410;
  assign _EVAL_154 = _EVAL_3003 | _EVAL_1706;
  assign _EVAL_2643 = _EVAL_2056 & _EVAL_3155;
  assign _EVAL_1425 = 9'he == _EVAL_1399 ? _EVAL_3670 : _EVAL_1149;
  assign _EVAL_2920 = _EVAL_551 != 8'h0;
  assign _EVAL_1213 = 9'hd == _EVAL_1399 ? 32'h10002223 : _EVAL_820;
  assign _EVAL_3576 = 9'h132 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1357;
  assign _EVAL_952 = _EVAL_700 & _EVAL_1303;
  assign _EVAL_2598 = _EVAL_1375 | _EVAL_2698;
  assign _EVAL_225 = 9'h1ea == _EVAL_1399 ? _EVAL_1856 : _EVAL_1991;
  assign _EVAL_1902 = 9'h185 == _EVAL_1399 ? _EVAL_374 : _EVAL_3500;
  assign _EVAL_2138 = _EVAL_3207[22:20];
  assign _EVAL_2190 = _EVAL_683 | _EVAL_272;
  assign _EVAL_3652 = _EVAL_1123 | _EVAL_654;
  assign _EVAL_2506 = 9'he2 == _EVAL_1399 ? 32'h0 : _EVAL_49;
  assign _EVAL_3299 = 9'h194 == _EVAL_1399 ? _EVAL_1856 : _EVAL_484;
  assign _EVAL_3586 = 9'h171 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1821;
  assign _EVAL_3591 = 9'h150 == _EVAL_1399 ? _EVAL_374 : _EVAL_841;
  assign _EVAL_3738 = 9'hd7 == _EVAL_1399 ? 32'h0 : _EVAL_790;
  assign _EVAL_3464 = 9'h174 == _EVAL_1399 ? _EVAL_374 : _EVAL_251;
  assign _EVAL_2274 = _EVAL_1176 ? {{9'd0}, _EVAL_147} : _EVAL_3349;
  assign _EVAL_3039 = _EVAL_696 | _EVAL_2291;
  assign _EVAL_2583 = _EVAL_1771 & _EVAL_1380;
  assign _EVAL_1460 = _EVAL_209 & _EVAL_234;
  assign _EVAL_2368 = 9'h6 == _EVAL_1399 ? 32'h10802023 : _EVAL_1942;
  assign _EVAL_686 = 9'h166 == _EVAL_1399 ? _EVAL_374 : _EVAL_1724;
  assign _EVAL_951 = _EVAL_607 | _EVAL_3339;
  assign _EVAL_1182 = 9'h6d == _EVAL_1399;
  assign _EVAL_3698 = 9'h62 == _EVAL_1399;
  assign _EVAL_3459 = 9'h18c == _EVAL_1399 ? _EVAL_374 : _EVAL_2251;
  assign _EVAL_442 = 9'hd3 == _EVAL_1399 ? 32'h0 : _EVAL_1167;
  assign _EVAL_1224 = 9'h1e7 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1040;
  assign _EVAL_2090 = 9'h140 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1307;
  assign _EVAL_2422 = _EVAL_2662 == 8'hff;
  assign _EVAL_3763 = _EVAL_1051 ? _EVAL_2188 : _EVAL_3100;
  assign _EVAL_2476 = 9'h1d3 == _EVAL_1399 ? _EVAL_374 : _EVAL_2615;
  assign _EVAL_3428 = 9'hc9 == _EVAL_1399 ? 32'h0 : _EVAL_2932;
  assign _EVAL_1087 = 9'h105 == _EVAL_1399 ? _EVAL_374 : _EVAL_393;
  assign _EVAL_3795 = _EVAL_1184 & _EVAL_234;
  assign _EVAL_1979 = 9'h5f == _EVAL_1399;
  assign _EVAL_2888 = _EVAL_3134 | _EVAL_3252;
  assign _EVAL_3388 = 9'h89 == _EVAL_1399;
  assign _EVAL_2216 = 9'h4a == _EVAL_1399 ? 32'h0 : _EVAL_2653;
  assign _EVAL_320 = 9'he3 == _EVAL_1399;
  assign _EVAL_3682 = {_EVAL_555,_EVAL_266,_EVAL_2757,_EVAL_2720};
  assign _EVAL_1057 = 9'h1d9 == _EVAL_1399 ? _EVAL_1856 : _EVAL_606;
  assign _EVAL_2769 = 9'h126 == _EVAL_1399 ? _EVAL_1856 : _EVAL_739;
  assign _EVAL_2845 = _EVAL_563 & _EVAL_3101;
  assign _EVAL_768 = _EVAL_1979 | _EVAL_1512;
  assign _EVAL_654 = _EVAL_3480 | _EVAL_3723;
  assign _EVAL_1243 = 9'h17d == _EVAL_1399 ? _EVAL_374 : _EVAL_2979;
  assign _EVAL_1037 = _EVAL_724 & _EVAL_234;
  assign _EVAL_2628 = _EVAL_575[10:8];
  assign _EVAL_3279 = 9'h1d0 == _EVAL_1399 ? _EVAL_374 : _EVAL_1571;
  assign _EVAL_710 = _EVAL_724 | _EVAL_2594;
  assign _EVAL_3583 = 9'h72 == _EVAL_1399 ? 32'h0 : _EVAL_312;
  assign _EVAL_2111 = 9'hcd == _EVAL_1399;
  assign _EVAL_1732 = 9'h19b == _EVAL_1399 ? _EVAL_374 : _EVAL_3539;
  assign _EVAL_1975 = 9'h3d == _EVAL_1399;
  assign _EVAL_1589 = _EVAL_563 & _EVAL_2081;
  assign _EVAL_2569 = _EVAL_866 | _EVAL_2219;
  assign _EVAL_754 = _EVAL_1177 | _EVAL_3652;
  assign _EVAL_721 = 9'h17e == _EVAL_1399 ? _EVAL_1856 : _EVAL_2383;
  assign _EVAL_2402 = 9'h59 == _EVAL_1399;
  assign _EVAL_275 = _EVAL_470 & _EVAL_2400;
  assign _EVAL_1641 = 9'he4 == _EVAL_1399 ? 32'h0 : _EVAL_538;
  assign _EVAL_474 = _EVAL_642 & _EVAL_2422;
  assign _EVAL_3830 = 9'h158 == _EVAL_1399 ? _EVAL_374 : _EVAL_198;
  assign _EVAL_2162 = 9'h1b2 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1341;
  assign _EVAL_890 = 9'h1c1 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2704;
  assign _EVAL_1 = _EVAL_14;
  assign _EVAL_2730 = 9'h47 == _EVAL_1399 ? 32'h0 : _EVAL_3411;
  assign _EVAL_3221 = ~_EVAL_2004;
  assign _EVAL_3823 = 9'h12e == _EVAL_1399 ? _EVAL_1856 : _EVAL_2858;
  assign _EVAL_3816 = 9'h2f == _EVAL_1399;
  assign _EVAL_3824 = _EVAL_2988 & _EVAL_234;
  assign _EVAL_2136 = 9'h1ac == _EVAL_1399 ? _EVAL_1856 : _EVAL_3568;
  assign _EVAL_1114 = 9'h160 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2519;
  assign _EVAL_700 = _EVAL_2414 & _EVAL_2188;
  assign _EVAL_3116 = _EVAL_1699 ? 8'hff : 8'h0;
  assign _EVAL_1859 = _EVAL_488 | _EVAL_2994;
  assign _EVAL_2951 = _EVAL_3772 | _EVAL_2354;
  assign _EVAL_551 = _EVAL_575[7:0];
  assign _EVAL_2996 = _EVAL_1752 & _EVAL_234;
  assign _EVAL_3500 = 9'h184 == _EVAL_1399 ? _EVAL_374 : _EVAL_1977;
  assign _EVAL_1982 = 9'h1d5 == _EVAL_1399 ? _EVAL_374 : _EVAL_1807;
  assign _EVAL_2775 = 9'hb0 == _EVAL_1399 ? 32'h0 : _EVAL_942;
  assign _EVAL_2749 = _EVAL_2628 == 3'h7;
  assign _EVAL_83 = 32'h1 << _EVAL_958;
  assign _EVAL_3524 = _EVAL_2911 | _EVAL_2419;
  assign _EVAL_2961 = _EVAL_997 & _EVAL_3761;
  assign _EVAL_2261 = _EVAL_11[15:8];
  assign _EVAL_3613 = 9'h60 == _EVAL_1399;
  assign _EVAL_2095 = 9'h1d8 == _EVAL_1399 ? _EVAL_374 : _EVAL_485;
  assign _EVAL_748 = _EVAL_3558[4];
  assign _EVAL_3182 = _EVAL_1675 & _EVAL_502;
  assign _EVAL_1226 = 9'h1f3 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3600;
  assign _EVAL_2392 = 9'h18e == _EVAL_1399 ? _EVAL_374 : _EVAL_324;
  assign _EVAL_3280 = 9'h1c3 == _EVAL_1399 ? _EVAL_1856 : _EVAL_402;
  assign _EVAL_3606 = 9'hdc == _EVAL_1399 ? _EVAL_1856 : _EVAL_2080;
  assign _EVAL_836 = _EVAL_2437 & _EVAL_2262;
  assign _EVAL_98 = 9'h1a2 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3668;
  assign _EVAL_965 = 9'hf7 == _EVAL_1399;
  assign _EVAL_353 = 9'h197 == _EVAL_1399 ? _EVAL_374 : _EVAL_2222;
  assign _EVAL_3804 = 9'h179 == _EVAL_1399 ? _EVAL_374 : _EVAL_2295;
  assign _EVAL_1824 = _EVAL_2743[64];
  assign _EVAL_152 = 9'h84 == _EVAL_1399 ? 32'h0 : _EVAL_3377;
  assign _EVAL_3254 = 9'hff == _EVAL_1399;
  assign _EVAL_3426 = 5'h1 == _EVAL_958;
  assign _EVAL_1014 = 9'h16f == _EVAL_1399 ? _EVAL_1856 : _EVAL_94;
  assign _EVAL_1755 = 9'h17b == _EVAL_1399 ? _EVAL_374 : _EVAL_1578;
  assign _EVAL_2821 = 9'hbd == _EVAL_1399 ? 32'h0 : _EVAL_2326;
  assign _EVAL_2744 = 9'h185 == _EVAL_1399 ? _EVAL_1856 : _EVAL_121;
  assign _EVAL_1274 = _EVAL_3281 | _EVAL_124;
  assign _EVAL_809 = 9'h32 == _EVAL_1399 ? 32'h0 : _EVAL_722;
  assign _EVAL_115 = 9'h78 == _EVAL_1399;
  assign _EVAL_27 = _EVAL_33;
  assign _EVAL_3456 = 9'h11e == _EVAL_1399 ? _EVAL_1856 : _EVAL_795;
  assign _EVAL_2595 = 9'h1b0 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1597;
  assign _EVAL_2742 = _EVAL_130 | _EVAL_3783;
  assign _EVAL_1942 = 9'h5 == _EVAL_1399 ? 32'hf1402473 : _EVAL_492;
  assign _EVAL_727 = 9'h20 == _EVAL_1399 ? 32'h0 : _EVAL_2463;
  assign _EVAL_1771 = _EVAL_1181 & _EVAL_1135;
  assign _EVAL_2610 = 9'h18a == _EVAL_1399 ? _EVAL_1856 : _EVAL_636;
  assign _EVAL_3447 = 9'h1e5 == _EVAL_1399 ? _EVAL_1856 : _EVAL_187;
  assign _EVAL_1467 = _EVAL_1475 & _EVAL_1856;
  assign _EVAL_2746 = _EVAL_2714 & _EVAL_234;
  assign _EVAL_1891 = 9'h124 == _EVAL_1399 ? _EVAL_1856 : _EVAL_205;
  assign _EVAL_3236 = 9'ha1 == _EVAL_1399;
  assign _EVAL_669 = 9'h1b2 == _EVAL_1399 ? _EVAL_374 : _EVAL_2989;
  assign _EVAL_2659 = 9'h193 == _EVAL_1399 ? _EVAL_374 : _EVAL_2508;
  assign _EVAL_753 = _EVAL_1127 | _EVAL_236;
  assign _EVAL_876 = 9'h26 == _EVAL_1399;
  assign _EVAL_866 = 9'h3a == _EVAL_1399;
  assign _EVAL_2878 = 9'h12f == _EVAL_1399 ? _EVAL_1856 : _EVAL_3823;
  assign _EVAL_3071 = 9'h61 == _EVAL_1399 ? 32'h0 : _EVAL_1934;
  assign _EVAL_35 = _EVAL_20;
  assign _EVAL_372 = _EVAL_174 | _EVAL_1728;
  assign _EVAL_2624 = _EVAL_11[10:8];
  assign _EVAL_2367 = 9'h1f9 == _EVAL_1399 ? _EVAL_374 : _EVAL_1328;
  assign _EVAL_3187 = 9'h133 == _EVAL_1399 ? _EVAL_374 : _EVAL_2002;
  assign _EVAL_1853 = 9'h17 == _EVAL_1399 ? 32'h0 : _EVAL_1343;
  assign _EVAL_891 = 9'h121 == _EVAL_1399 ? _EVAL_374 : _EVAL_546;
  assign _EVAL_895 = 9'ha6 == _EVAL_1399;
  assign _EVAL_972 = 9'hdd == _EVAL_1399 ? _EVAL_3031 : _EVAL_486;
  assign _EVAL_3235 = _EVAL_2178 | _EVAL_3230;
  assign _EVAL_2145 = _EVAL_1921 | _EVAL_2709;
  assign _EVAL_2125 = 9'h82 == _EVAL_1399 ? 32'h0 : _EVAL_3604;
  assign _EVAL_2731 = 9'hd1 == _EVAL_1399;
  assign _EVAL_3809 = _EVAL_2265 | _EVAL_1896;
  assign _EVAL_784 = _EVAL_1839 | _EVAL_1132;
  assign _EVAL_72 = 9'h12 == _EVAL_1399 ? 32'h7b200073 : _EVAL_1026;
  assign _EVAL_2816 = 9'h114 == _EVAL_1399 ? _EVAL_374 : _EVAL_1653;
  assign _EVAL_3612 = 9'h14a == _EVAL_1399 ? _EVAL_1856 : _EVAL_3508;
  assign _EVAL_1478 = 9'h111 == _EVAL_1399 ? _EVAL_374 : _EVAL_908;
  assign _EVAL_662 = 9'hd0 == _EVAL_1399 ? 32'h0 : _EVAL_1992;
  assign _EVAL_1569 = _EVAL_2847 | _EVAL_2627;
  assign _EVAL_3200 = 9'h5b == _EVAL_1399 ? 32'h0 : _EVAL_1007;
  assign _EVAL_308 = 9'h107 == _EVAL_1399 ? _EVAL_374 : _EVAL_3409;
  assign _EVAL_3723 = _EVAL_363 | _EVAL_651;
  assign _EVAL_2256 = _EVAL_3457 | _EVAL_2598;
  assign _EVAL_1933 = 9'h7a == _EVAL_1399 ? 32'h0 : _EVAL_2471;
  assign _EVAL_1437 = _EVAL_1471 | _EVAL_2961;
  assign _EVAL_2008 = 9'he4 == _EVAL_1399;
  assign _EVAL_567 = 9'h1ec == _EVAL_1399 ? _EVAL_374 : _EVAL_1516;
  assign _EVAL_2635 = 9'h68 == _EVAL_1399;
  assign _EVAL_3143 = _EVAL_11[23:16];
  assign _EVAL_3495 = _EVAL_169 ? _EVAL_547 : _EVAL_1435;
  assign _EVAL_3519 = _EVAL_1771 & _EVAL_1303;
  assign _EVAL_1842 = {7'h1c,_EVAL_957,5'h0,_EVAL_2138,5'h0,7'h23};
  assign _EVAL_3276 = 9'h2f == _EVAL_1399 ? 32'h0 : _EVAL_2496;
  assign _EVAL_3469 = 9'h12d == _EVAL_1399 ? _EVAL_374 : _EVAL_2928;
  assign _EVAL_23 = _EVAL_40;
  assign _EVAL_3316 = 9'ha9 == _EVAL_1399 ? 32'h0 : _EVAL_2619;
  assign _EVAL_3369 = _EVAL_2828 | _EVAL_1888;
  assign _EVAL_3417 = _EVAL_3588 & _EVAL_234;
  assign _EVAL_2974 = 9'h39 == _EVAL_1399;
  assign _EVAL_94 = 9'h16e == _EVAL_1399 ? _EVAL_1856 : _EVAL_3545;
  assign _EVAL_2758 = 9'h1cc == _EVAL_1399 ? _EVAL_1856 : _EVAL_2837;
  assign _EVAL_506 = 9'h2d == _EVAL_1399;
  assign _EVAL_1023 = 9'h93 == _EVAL_1399;
  assign _EVAL_3506 = 9'h186 == _EVAL_1399 ? _EVAL_374 : _EVAL_1902;
  assign _EVAL_2411 = _EVAL_1675 & _EVAL_1897;
  assign _EVAL_3067 = 9'h26 == _EVAL_1399 ? 32'h0 : _EVAL_765;
  assign _EVAL_2921 = 9'h154 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3379;
  assign _EVAL_117 = _EVAL_421 & _EVAL_2604;
  assign _EVAL_2899 = 9'h13d == _EVAL_1399 ? _EVAL_1856 : _EVAL_1747;
  assign _EVAL_3425 = ~_EVAL_18;
  assign _EVAL_2432 = 9'heb == _EVAL_1399 ? 32'h0 : _EVAL_436;
  assign _EVAL_960 = 9'h172 == _EVAL_1399 ? _EVAL_374 : _EVAL_2895;
  assign _EVAL_3762 = 9'h15d == _EVAL_1399 ? _EVAL_1856 : _EVAL_71;
  assign _EVAL_2725 = 9'h1b == _EVAL_1399;
  assign _EVAL_470 = _EVAL_1987 == 2'h2;
  assign _EVAL_2686 = 9'h1e2 == _EVAL_1399 ? _EVAL_374 : _EVAL_2217;
  assign _EVAL_1357 = 9'h131 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1450;
  assign _EVAL_1769 = 9'h199 == _EVAL_1399 ? _EVAL_1856 : _EVAL_516;
  assign _EVAL_3203 = _EVAL_17 & _EVAL_25;
  assign _EVAL_1675 = _EVAL_2056 & _EVAL_2302;
  assign _EVAL_1860 = _EVAL_558 | _EVAL_3212;
  assign _EVAL_3115 = 9'h134 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3727;
  assign _EVAL_2440 = 9'h1aa == _EVAL_1399 ? _EVAL_374 : _EVAL_1799;
  assign _EVAL_2648 = 9'h119 == _EVAL_1399 ? _EVAL_1856 : _EVAL_415;
  assign _EVAL_2398 = 9'h155 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2921;
  assign _EVAL_2994 = _EVAL_982 | _EVAL_760;
  assign _EVAL_156 = 9'hc4 == _EVAL_1399;
  assign _EVAL_642 = _EVAL_836 & _EVAL_1856;
  assign _EVAL_1774 = 9'h146 == _EVAL_1399 ? _EVAL_374 : _EVAL_2233;
  assign _EVAL_993 = 9'h156 == _EVAL_1399 ? _EVAL_374 : _EVAL_184;
  assign _EVAL_1578 = 9'h17a == _EVAL_1399 ? _EVAL_374 : _EVAL_3804;
  assign _EVAL_1149 = 9'hd == _EVAL_1399 ? _EVAL_3670 : _EVAL_1069;
  assign _EVAL_2359 = 9'h47 == _EVAL_1399;
  assign _EVAL_1495 = 9'h129 == _EVAL_1399 ? _EVAL_374 : _EVAL_3194;
  assign _EVAL_3264 = _EVAL_3782 & _EVAL_1883;
  assign _EVAL_3283 = 9'hb2 == _EVAL_1399;
  assign _EVAL_1841 = _EVAL_3247 & _EVAL_2819;
  assign _EVAL_2196 = 9'h174 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1767;
  assign _EVAL_2459 = 9'h6c == _EVAL_1399 ? 32'h0 : _EVAL_1639;
  assign _EVAL_332 = 9'h36 == _EVAL_1399 ? 32'h0 : _EVAL_2194;
  assign _EVAL_2217 = 9'h1e1 == _EVAL_1399 ? _EVAL_374 : _EVAL_3088;
  assign _EVAL_1697 = 9'hdf == _EVAL_1399 ? 32'h100073 : _EVAL_1004;
  assign _EVAL_2810 = 9'h18f == _EVAL_1399 ? _EVAL_1856 : _EVAL_713;
  assign _EVAL_3275 = 9'hf == _EVAL_1399 ? 32'hf1402473 : _EVAL_2591;
  assign _EVAL_3003 = 9'h48 == _EVAL_1399;
  assign _EVAL_943 = 9'h59 == _EVAL_1399 ? 32'h0 : _EVAL_2789;
  assign _EVAL_2908 = 9'h8 == _EVAL_1399 ? 32'h347413 : _EVAL_2452;
  assign _EVAL_2339 = _EVAL_705 | _EVAL_985;
  assign _EVAL_2761 = _EVAL_1163 | _EVAL_3030;
  assign _EVAL_3633 = _EVAL_1166 | _EVAL_2453;
  assign _EVAL_1140 = 9'h1e3 == _EVAL_1399 ? _EVAL_374 : _EVAL_2686;
  assign _EVAL_2573 = _EVAL_1773 | _EVAL_2395;
  assign _EVAL_3073 = 9'h8a == _EVAL_1399 ? 32'h0 : _EVAL_799;
  assign _EVAL_1051 = 5'he == _EVAL_958;
  assign _EVAL_147 = {1'h1,_EVAL_1592};
  assign _EVAL_2970 = 9'h1d == _EVAL_1399;
  assign _EVAL_3826 = 9'h139 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1314;
  assign _EVAL_2194 = 9'h35 == _EVAL_1399 ? 32'h0 : _EVAL_1370;
  assign _EVAL_2756 = _EVAL_2111 | _EVAL_2581;
  assign _EVAL_725 = _EVAL_870[3];
  assign _EVAL_1461 = 9'h1ed == _EVAL_1399 ? _EVAL_1856 : _EVAL_1508;
  assign _EVAL_3511 = _EVAL_762 | _EVAL_1654;
  assign _EVAL_3799 = _EVAL_3613 | _EVAL_768;
  assign _EVAL_363 = 9'h7a == _EVAL_1399;
  assign _EVAL_2705 = 9'h1d5 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1880;
  assign _EVAL_313 = 9'h6 == _EVAL_1399 ? _EVAL_3670 : _EVAL_2552;
  assign _EVAL_2841 = _EVAL_2333 | _EVAL_3555;
  assign _EVAL_265 = _EVAL_1023 | _EVAL_317;
  assign _EVAL_3123 = 9'h10c == _EVAL_1399 ? _EVAL_374 : _EVAL_2144;
  assign _EVAL_2358 = _EVAL_879 | _EVAL_2841;
  assign _EVAL_3310 = _EVAL_1089 | _EVAL_2501;
  assign _EVAL_2763 = _EVAL_995[31:24];
  assign _EVAL_3675 = 9'h1f0 == _EVAL_1399 ? _EVAL_374 : _EVAL_2417;
  assign _EVAL_3567 = 9'hfc == _EVAL_1399;
  assign _EVAL_2838 = 9'hf3 == _EVAL_1399;
  assign _EVAL_2336 = _EVAL_2445 & _EVAL_1018;
  assign _EVAL_121 = 9'h184 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1311;
  assign _EVAL_3038 = _EVAL_3203 & _EVAL_19;
  assign _EVAL_2347 = _EVAL_1675 & _EVAL_2499;
  assign _EVAL_614 = 9'h180 == _EVAL_1399 ? _EVAL_374 : _EVAL_1875;
  assign _EVAL_1486 = 9'h1b8 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3159;
  assign _EVAL_2104 = _EVAL_83[1];
  assign _EVAL_868 = 9'hd2 == _EVAL_1399;
  assign _EVAL_3724 = 9'h122 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3227;
  assign _EVAL_858 = 9'h14e == _EVAL_1399 ? _EVAL_374 : _EVAL_1731;
  assign _EVAL_984 = 9'h9c == _EVAL_1399;
  assign _EVAL_3023 = 9'h4 == _EVAL_1399 ? _EVAL_3670 : _EVAL_1334;
  assign _EVAL_3782 = _EVAL_2650 & _EVAL_1856;
  assign _EVAL_1978 = _EVAL_61 & 16'h3;
  assign _EVAL_3834 = 9'h18a == _EVAL_1399 ? _EVAL_374 : _EVAL_3695;
  assign _EVAL_3298 = 9'h12c == _EVAL_1399 ? _EVAL_1856 : _EVAL_2318;
  assign _EVAL_861 = _EVAL_3825 | _EVAL_2358;
  assign _EVAL_55 = 9'h91 == _EVAL_1399 ? 32'h0 : _EVAL_2173;
  assign _EVAL_572 = _EVAL_2845 | _EVAL_2583;
  assign _EVAL_833 = _EVAL_1097 | _EVAL_1859;
  assign _EVAL_1343 = 9'h16 == _EVAL_1399 ? 32'h0 : _EVAL_1591;
  assign _EVAL_1516 = 9'h1eb == _EVAL_1399 ? _EVAL_374 : _EVAL_110;
  assign _EVAL_1145 = _EVAL_2714 | _EVAL_952;
  assign _EVAL_1069 = 9'hc == _EVAL_1399 ? _EVAL_3670 : _EVAL_1021;
  assign _EVAL_1706 = _EVAL_2359 | _EVAL_2958;
  assign _EVAL_1046 = 9'h17a == _EVAL_1399 ? _EVAL_1856 : _EVAL_689;
  assign _EVAL_2650 = _EVAL_2437 & _EVAL_2488;
  assign _EVAL_498 = 9'h182 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2623;
  assign _EVAL_3106 = _EVAL_3588 & _EVAL_3485;
  assign debug_hartReset_0__EVAL = _EVAL_38;
  assign _EVAL_2735 = 9'h11f == _EVAL_1399 ? _EVAL_374 : _EVAL_707;
  assign _EVAL_790 = 9'hd6 == _EVAL_1399 ? 32'h0 : _EVAL_605;
  assign _EVAL_2655 = _EVAL_3337 == 7'h8;
  assign _EVAL_2089 = 9'h1dd == _EVAL_1399 ? _EVAL_374 : _EVAL_601;
  assign _EVAL_3755 = 9'hc5 == _EVAL_1399;
  assign _EVAL_547 = {{31'd0}, _EVAL_2157};
  assign _EVAL_54 = 9'hc3 == _EVAL_1399 ? 32'h0 : _EVAL_109;
  assign _EVAL_3155 = _EVAL_0 == 3'h4;
  assign _EVAL_3731 = _EVAL_2716 | _EVAL_3472;
  assign _EVAL_1544 = 9'h105 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2703;
  assign _EVAL_3052 = 9'hac == _EVAL_1399 ? 32'h0 : _EVAL_409;
  assign _EVAL_3836 = _EVAL_83[8];
  assign _EVAL_3043 = _EVAL_551 == 8'hff;
  assign _EVAL_2831 = 9'h8 == _EVAL_1399 ? _EVAL_3670 : _EVAL_229;
  assign _EVAL_2015 = 9'hed == _EVAL_1399 ? 32'h0 : _EVAL_1795;
  assign _EVAL_209 = _EVAL_3815 & _EVAL_3043;
  assign _EVAL_628 = 9'h1a7 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1081;
  assign _EVAL_3420 = _EVAL_386 ? _EVAL_1135 : _EVAL_2185;
  assign _EVAL_2290 = 9'h61 == _EVAL_1399;
  assign _EVAL_1268 = 9'h10f == _EVAL_1399 ? _EVAL_1856 : _EVAL_3238;
  assign _EVAL_1270 = 9'h177 == _EVAL_1399 ? _EVAL_374 : _EVAL_3754;
  assign _EVAL_3270 = 9'h19d == _EVAL_1399 ? _EVAL_374 : _EVAL_2780;
  assign _EVAL_3598 = 9'hca == _EVAL_1399 ? 32'h0 : _EVAL_3428;
  assign _EVAL_3220 = 9'h2d == _EVAL_1399 ? 32'h0 : _EVAL_3657;
  assign _EVAL_509 = 9'h57 == _EVAL_1399;
  assign _EVAL_2704 = 9'h1c0 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2077;
  assign _EVAL_3709 = 9'h126 == _EVAL_1399 ? _EVAL_374 : _EVAL_1154;
  assign _EVAL_419 = 9'h9b == _EVAL_1399 ? 32'h0 : _EVAL_1419;
  assign _EVAL_3485 = ~_EVAL_234;
  assign _EVAL_1598 = 9'h1ba == _EVAL_1399 ? _EVAL_374 : _EVAL_257;
  assign _EVAL_2755 = 9'h3a == _EVAL_1399 ? 32'h0 : _EVAL_3309;
  assign _EVAL_3379 = 9'h153 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3005;
  assign _EVAL_2480 = 9'h21 == _EVAL_1399 ? 32'h0 : _EVAL_727;
  assign _EVAL_702 = 9'h95 == _EVAL_1399 ? 32'h0 : _EVAL_2818;
  assign _EVAL_1880 = 9'h1d4 == _EVAL_1399 ? _EVAL_1856 : _EVAL_389;
  assign _EVAL_2006 = 9'h1bc == _EVAL_1399 ? _EVAL_374 : _EVAL_3265;
  assign _EVAL_2864 = _EVAL_2363[31:24];
  assign _EVAL_1321 = 9'h175 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2196;
  assign _EVAL_3493 = 9'h1ac == _EVAL_1399 ? _EVAL_374 : _EVAL_3589;
  assign _EVAL_304 = _EVAL_1335 ? 1'h0 : _EVAL_451;
  assign _EVAL_2794 = 9'h1c2 == _EVAL_1399 ? _EVAL_374 : _EVAL_956;
  assign _EVAL_3113 = _EVAL_26[23:16];
  assign _EVAL_1217 = _EVAL_575 == 32'hffffffff;
  assign _EVAL_3838 = _EVAL_2091 | _EVAL_3328;
  assign _EVAL_1012 = 9'h151 == _EVAL_1399 ? _EVAL_374 : _EVAL_3591;
  assign _EVAL_1650 = 9'h33 == _EVAL_1399;
  assign _EVAL_2073 = 9'h168 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3557;
  assign _EVAL_3356 = 9'h2c == _EVAL_1399;
  assign _EVAL_1407 = 9'h157 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3753;
  assign _EVAL_2280 = _EVAL_3806 ? 8'hff : 8'h0;
  assign _EVAL_634 = 9'h175 == _EVAL_1399 ? _EVAL_374 : _EVAL_3464;
  assign _EVAL_785 = 9'h14e == _EVAL_1399 ? _EVAL_1856 : _EVAL_458;
  assign _EVAL_3193 = 9'h55 == _EVAL_1399 ? 32'h0 : _EVAL_613;
  assign _EVAL_619 = 9'hc2 == _EVAL_1399;
  assign _EVAL_3481 = _EVAL_617 | _EVAL_3524;
  assign _EVAL_9 = _EVAL_3788 ? _EVAL_3146 : 32'h0;
  assign _EVAL_659 = _EVAL_2163 <= 16'h101f;
  assign _EVAL_1174 = 9'h27 == _EVAL_1399;
  assign _EVAL_3745 = 9'h1ae == _EVAL_1399 ? _EVAL_1856 : _EVAL_1066;
  assign _EVAL_3059 = 9'h140 == _EVAL_1399 ? _EVAL_374 : _EVAL_2750;
  assign _EVAL_1152 = _EVAL_1275 | _EVAL_1155;
  assign _EVAL_2075 = _EVAL_1523 ? 1'h0 : _EVAL_2218;
  assign _EVAL_1758 = 9'h176 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1321;
  assign _EVAL_3237 = _EVAL_2725 | _EVAL_1538;
  assign _EVAL_3262 = 9'h72 == _EVAL_1399;
  assign _EVAL_3009 = _EVAL_868 | _EVAL_526;
  assign _EVAL_906 = 9'h19c == _EVAL_1399 ? _EVAL_1856 : _EVAL_1561;
  assign _EVAL_153 = 9'h13b == _EVAL_1399 ? _EVAL_1856 : _EVAL_3717;
  assign _EVAL_3002 = 9'h1fc == _EVAL_1399 ? _EVAL_374 : _EVAL_228;
  assign _EVAL_365 = 9'h91 == _EVAL_1399;
  assign _EVAL_869 = 9'h139 == _EVAL_1399 ? _EVAL_374 : _EVAL_434;
  assign _EVAL_724 = _EVAL_1273 & _EVAL_3043;
  assign _EVAL_2560 = 9'h1d7 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1071;
  assign _EVAL_689 = 9'h179 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2636;
  assign _EVAL_1653 = 9'h113 == _EVAL_1399 ? _EVAL_374 : _EVAL_3271;
  assign _EVAL_3751 = _EVAL_1564 | _EVAL_3710;
  assign _EVAL_2604 = _EVAL_3395 ? 1'h0 : _EVAL_1228;
  assign _EVAL_2463 = 9'h1f == _EVAL_1399 ? 32'h0 : _EVAL_2429;
  assign _EVAL_493 = 9'h2a == _EVAL_1399;
  assign _EVAL_638 = _EVAL_2743[67];
  assign _EVAL_1304 = 9'hb3 == _EVAL_1399;
  assign _EVAL_1285 = 9'h6f == _EVAL_1399 ? 32'h0 : _EVAL_3326;
  assign _EVAL_1823 = 9'h11b == _EVAL_1399 ? _EVAL_374 : _EVAL_837;
  assign _EVAL_1400 = _EVAL_3498 & _EVAL_1151;
  assign _EVAL_1041 = 9'h13d == _EVAL_1399 ? _EVAL_374 : _EVAL_723;
  assign _EVAL_3359 = 9'h40 == _EVAL_1399 ? 32'h0 : _EVAL_2842;
  assign _EVAL_1953 = 9'h1d1 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1044;
  assign _EVAL_88 = _EVAL_167[0];
  assign _EVAL_2801 = 9'h1c7 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1518;
  assign _EVAL_1218 = _EVAL_3677[17:0];
  assign _EVAL_3671 = 9'h167 == _EVAL_1399 ? _EVAL_374 : _EVAL_686;
  assign _EVAL_1773 = 9'h80 == _EVAL_1399;
  assign _EVAL_258 = 9'h63 == _EVAL_1399 ? 32'h0 : _EVAL_3499;
  assign _EVAL_2193 = 9'h1f5 == _EVAL_1399 ? _EVAL_374 : _EVAL_1514;
  assign _EVAL_1761 = _EVAL_3782 & _EVAL_1151;
  assign _EVAL_1934 = 9'h60 == _EVAL_1399 ? 32'h0 : _EVAL_3250;
  assign _EVAL_2854 = 9'h170 == _EVAL_1399 ? _EVAL_374 : _EVAL_3661;
  assign _EVAL_78 = 9'h12e == _EVAL_1399 ? _EVAL_374 : _EVAL_3469;
  assign _EVAL_3482 = _EVAL_734 ? 1'h0 : 1'h1;
  assign _EVAL_1096 = 9'h1b0 == _EVAL_1399 ? _EVAL_374 : _EVAL_3476;
  assign _EVAL_481 = _EVAL_3742 | _EVAL_1332;
  assign _EVAL_2121 = _EVAL_93 | _EVAL_1713;
  assign _EVAL_215 = _EVAL_612 == 2'h3;
  assign _EVAL_1040 = 9'h1e6 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3447;
  assign _EVAL_1426 = 9'h98 == _EVAL_1399;
  assign _EVAL_93 = 9'h34 == _EVAL_1399;
  assign _EVAL_3717 = 9'h13a == _EVAL_1399 ? _EVAL_1856 : _EVAL_3826;
  assign _EVAL_3085 = _EVAL_28[0];
  assign _EVAL_1983 = _EVAL_2005 | _EVAL_2168;
  assign _EVAL_1832 = 9'hd4 == _EVAL_1399 ? 32'h0 : _EVAL_442;
  assign _EVAL_546 = 9'h120 == _EVAL_1399 ? _EVAL_374 : _EVAL_2735;
  assign _EVAL_554 = 9'hf4 == _EVAL_1399;
  assign _EVAL_2709 = _EVAL_3593 | _EVAL_214;
  assign _EVAL_2819 = _EVAL_1682 == 10'h3ff;
  assign _EVAL_3250 = 9'h5f == _EVAL_1399 ? 32'h0 : _EVAL_2078;
  assign _EVAL_1872 = _EVAL_3254 | _EVAL_2014;
  assign _EVAL_2481 = 9'h151 == _EVAL_1399 ? _EVAL_1856 : _EVAL_622;
  assign _EVAL_1351 = 9'h8c == _EVAL_1399 ? 32'h0 : _EVAL_2687;
  assign _EVAL_1779 = 9'h1c3 == _EVAL_1399 ? _EVAL_374 : _EVAL_2794;
  assign _EVAL_2491 = 9'h79 == _EVAL_1399;
  assign _EVAL_1335 = _EVAL_217 & _EVAL_2819;
  assign _EVAL_133 = 9'h65 == _EVAL_1399 ? 32'h0 : _EVAL_1276;
  assign _EVAL_3152 = _EVAL_2163 & 16'h1f;
  assign _EVAL_2750 = 9'h13f == _EVAL_1399 ? _EVAL_374 : _EVAL_909;
  assign _EVAL_2083 = _EVAL_156 | _EVAL_1220;
  assign _EVAL_3101 = _EVAL_2264 == 8'hff;
  assign _EVAL_3100 = _EVAL_3027 ? _EVAL_2188 : _EVAL_279;
  assign _EVAL_1681 = _EVAL_234 ? 1'h0 : _EVAL_2896;
  assign _EVAL_1599 = _EVAL_1020 | _EVAL_1822;
  assign _EVAL_2472 = 9'hcf == _EVAL_1399;
  assign _EVAL_1297 = 9'h117 == _EVAL_1399 ? _EVAL_374 : _EVAL_3025;
  assign _EVAL_3806 = _EVAL_29[1];
  assign _EVAL_2590 = _EVAL_674 | _EVAL_1031;
  assign _EVAL_1200 = 9'h1a3 == _EVAL_1399 ? _EVAL_374 : _EVAL_2284;
  assign _EVAL_2091 = 9'h75 == _EVAL_1399;
  assign _EVAL_384 = 9'h4b == _EVAL_1399;
  assign _EVAL_2333 = 9'he7 == _EVAL_1399;
  assign _EVAL_3475 = 9'h187 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3596;
  assign _EVAL_1133 = 9'h16d == _EVAL_1399 ? _EVAL_374 : _EVAL_653;
  assign _EVAL_249 = 9'h74 == _EVAL_1399 ? 32'h0 : _EVAL_1849;
  assign _EVAL_1328 = 9'h1f8 == _EVAL_1399 ? _EVAL_374 : _EVAL_1685;
  assign _EVAL_1082 = _EVAL_2163 >= 16'h1000;
  assign _EVAL_3233 = 9'h1f4 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1226;
  assign _EVAL_421 = _EVAL_1987 == 2'h1;
  assign _EVAL_2913 = 9'h86 == _EVAL_1399 ? 32'h0 : _EVAL_2299;
  assign _EVAL_123 = 9'h7b == _EVAL_1399 ? 32'h0 : _EVAL_1933;
  assign _EVAL_711 = 9'h144 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3183;
  assign _EVAL_3159 = 9'h1b7 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3103;
  assign _EVAL_205 = 9'h123 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3724;
  assign _EVAL_728 = _EVAL_3343 | _EVAL_3020;
  assign _EVAL_3004 = 9'h13 == _EVAL_1399 ? 32'h10002623 : _EVAL_72;
  assign _EVAL_1994 = 9'hf9 == _EVAL_1399 ? 32'h0 : _EVAL_268;
  assign _EVAL_1380 = _EVAL_2264 != 8'h0;
  assign _EVAL_1219 = 9'h2a == _EVAL_1399 ? 32'h0 : _EVAL_1469;
  assign _EVAL_569 = 9'h16c == _EVAL_1399 ? _EVAL_1856 : _EVAL_620;
  assign _EVAL_3177 = ~_EVAL_3105;
  assign _EVAL_653 = 9'h16c == _EVAL_1399 ? _EVAL_374 : _EVAL_1147;
  assign _EVAL_2581 = _EVAL_202 | _EVAL_2412;
  assign _EVAL_2054 = 9'h15a == _EVAL_1399 ? _EVAL_1856 : _EVAL_2589;
  assign _EVAL_431 = 9'h17b == _EVAL_1399 ? _EVAL_1856 : _EVAL_1046;
  assign _EVAL_613 = 9'h54 == _EVAL_1399 ? 32'h0 : _EVAL_2255;
  assign _EVAL_2116 = 9'h1e8 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1224;
  assign _EVAL_2988 = _EVAL_1273 & _EVAL_2081;
  assign _EVAL_2524 = _EVAL_233 | _EVAL_2166;
  assign _EVAL_2965 = _EVAL_2103 | _EVAL_2674;
  assign _EVAL_2780 = 9'h19c == _EVAL_1399 ? _EVAL_374 : _EVAL_1732;
  assign _EVAL_683 = 9'ha2 == _EVAL_1399;
  assign _EVAL_867 = _EVAL_2707 | _EVAL_1798;
  assign _EVAL_2157 = _EVAL_910 != 32'h0;
  assign debug_hartReset_0__EVAL_2 = _EVAL_7;
  assign _EVAL_1303 = _EVAL_1319 != 8'h0;
  assign _EVAL_464 = _EVAL_2786 & _EVAL_2655;
  assign _EVAL_969 = 9'h197 == _EVAL_1399 ? _EVAL_1856 : _EVAL_3839;
  assign _EVAL_769 = 9'h8e == _EVAL_1399;
  assign _EVAL_3047 = 9'hbd == _EVAL_1399;
  assign _EVAL_3154 = 9'h190 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2810;
  assign _EVAL_2727 = _EVAL_575[23:16];
  assign _EVAL_1615 = 9'h76 == _EVAL_1399 ? 32'h0 : _EVAL_1900;
  assign _EVAL_1747 = 9'h13c == _EVAL_1399 ? _EVAL_1856 : _EVAL_153;
  assign _EVAL_2149 = _EVAL_493 | _EVAL_802;
  assign _EVAL_2188 = _EVAL_3337 == 7'h0;
  assign _EVAL_617 = 9'h4d == _EVAL_1399;
  assign _EVAL_311 = 9'hce == _EVAL_1399 ? 32'h0 : _EVAL_1545;
  assign _EVAL_3393 = _EVAL_2590 | _EVAL_3436;
  assign _EVAL_886 = _EVAL_3356 | _EVAL_2340;
  assign _EVAL_879 = 9'he8 == _EVAL_1399;
  assign debug_hartReset_0__EVAL_0 = _EVAL;
  assign _EVAL_1339 = {{11'd0}, _EVAL_2324};
  assign _EVAL_17 = 1'h1;
  assign _EVAL_143 = 9'hb4 == _EVAL_1399 ? 32'h0 : _EVAL_3688;
  assign _EVAL_2178 = 9'h55 == _EVAL_1399;
  assign _EVAL_2294 = 9'h11b == _EVAL_1399 ? _EVAL_1856 : _EVAL_3076;
  assign _EVAL_2453 = _EVAL_2855 | _EVAL_3001;
  assign _EVAL_3748 = 9'hfe == _EVAL_1399 ? 32'h0 : _EVAL_118;
  assign _EVAL_1184 = _EVAL_2807 & _EVAL_1217;
  assign _EVAL_126 = 9'h1f8 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1136;
  assign _EVAL_734 = _EVAL_1721 | _EVAL_1590;
  assign _EVAL_1376 = _EVAL_3498 & _EVAL_1883;
  assign _EVAL_3670 = _EVAL_306 == 10'h200;
  assign _EVAL_1433 = 9'h74 == _EVAL_1399;
  assign _EVAL_3122 = _EVAL_3837 | _EVAL_265;
  assign _EVAL_1576 = {_EVAL_3050,_EVAL_3777,_EVAL_1894,_EVAL_3138};
  assign _EVAL_1312 = 9'hbf == _EVAL_1399 ? 32'h0 : _EVAL_2517;
  assign _EVAL_3288 = 9'hae == _EVAL_1399 ? 32'h0 : _EVAL_540;
  assign _EVAL_1532 = 9'h5d == _EVAL_1399 ? 32'h0 : _EVAL_1139;
  assign _EVAL_982 = 9'h1e == _EVAL_1399;
  assign _EVAL_1034 = 9'hc6 == _EVAL_1399;
  assign _EVAL_1606 = _EVAL_895 | _EVAL_333;
  assign _EVAL_2175 = 9'h1e2 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2937;
  assign _EVAL_3088 = 9'h1e0 == _EVAL_1399 ? _EVAL_374 : _EVAL_2143;
  assign _EVAL_3045 = 9'h12 == _EVAL_1399 ? _EVAL_3670 : _EVAL_2741;
  assign _EVAL_3144 = _EVAL_2041 | _EVAL_2190;
  assign _EVAL_58 = 9'h194 == _EVAL_1399 ? _EVAL_374 : _EVAL_2659;
  assign _EVAL_3157 = 9'h14a == _EVAL_1399 ? _EVAL_374 : _EVAL_125;
  assign _EVAL_1314 = 9'h138 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2308;
  assign _EVAL_736 = 9'ha4 == _EVAL_1399;
  assign _EVAL_344 = 9'h1ee == _EVAL_1399 ? _EVAL_374 : _EVAL_766;
  assign _EVAL_1030 = 9'h1cd == _EVAL_1399 ? _EVAL_374 : _EVAL_2584;
  assign _EVAL_1044 = 9'h1d0 == _EVAL_1399 ? _EVAL_1856 : _EVAL_171;
  assign _EVAL_3385 = _EVAL_3558[1];
  assign _EVAL_2890 = 9'h1d == _EVAL_1399 ? 32'h0 : _EVAL_735;
  assign _EVAL_200 = _EVAL_1273 & _EVAL_3101;
  assign _EVAL_2452 = 9'h7 == _EVAL_1399 ? 32'h40044403 : _EVAL_2368;
  assign _EVAL_150 = 9'h87 == _EVAL_1399;
  assign _EVAL_2508 = 9'h192 == _EVAL_1399 ? _EVAL_374 : _EVAL_1436;
  assign _EVAL_2955 = 9'h81 == _EVAL_1399;
  assign _EVAL_2264 = _EVAL_575[31:24];
  assign _EVAL_3637 = 9'hb2 == _EVAL_1399 ? 32'h0 : _EVAL_1593;
  assign _EVAL_1911 = _EVAL_2455 | _EVAL_1052;
  assign _EVAL_3558 = _EVAL_21[8:2];
  assign _EVAL_1728 = _EVAL_1803 | _EVAL_3122;
  assign _EVAL_386 = 5'h0 == _EVAL_958;
  assign _EVAL_3320 = 9'h9d == _EVAL_1399 ? 32'h0 : _EVAL_2512;
  assign _EVAL_1701 = 9'h29 == _EVAL_1399;
  assign _EVAL_793 = 5'ha == _EVAL_958;
  assign _EVAL_2235 = 9'hd0 == _EVAL_1399;
  assign _EVAL_505 = _EVAL_685 | _EVAL_2115;
  assign _EVAL_2332 = 9'h1f6 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1408;
  assign _EVAL_2494 = 9'h1f1 == _EVAL_1399 ? _EVAL_374 : _EVAL_3675;
  assign _EVAL_707 = 9'h11e == _EVAL_1399 ? _EVAL_374 : _EVAL_2360;
  assign _EVAL_630 = 9'h1c9 == _EVAL_1399 ? _EVAL_374 : _EVAL_212;
  assign _EVAL_2166 = _EVAL_3262 | _EVAL_1198;
  assign _EVAL_3714 = 9'h1b5 == _EVAL_1399 ? _EVAL_1856 : _EVAL_1098;
  assign _EVAL_3171 = 9'h1e3 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2175;
  assign _EVAL_1568 = 9'h102 == _EVAL_1399 ? _EVAL_1856 : _EVAL_2684;
  assign _EVAL_2156 = _EVAL_3662 ? _EVAL_2655 : _EVAL_3160;
  assign _EVAL_1721 = ~_EVAL_1562;
  assign _EVAL_1685 = 9'h1f7 == _EVAL_1399 ? _EVAL_374 : _EVAL_3526;
  assign _EVAL_530 = _EVAL_1620 ? 8'hff : 8'h0;
  assign _EVAL_3231 = 9'h181 == _EVAL_1399 ? _EVAL_374 : _EVAL_614;
  assign _EVAL_2893 = 9'h1fc == _EVAL_1399 ? _EVAL_1856 : _EVAL_3722;
  assign _EVAL_645 = _EVAL_3369 & _EVAL_88;
  assign _EVAL_2325 = _EVAL_200 | _EVAL_3268;
  assign _EVAL_1050 = _EVAL_234 ? 1'h0 : _EVAL_117;
  assign _EVAL_2958 = _EVAL_439 | _EVAL_1665;
  assign _EVAL_343 = _EVAL_2451 | _EVAL_2339;
  assign _EVAL_2479 = _EVAL_1008 | _EVAL_510;
  assign _EVAL_1039 = _EVAL_583 | _EVAL_941;
  assign _EVAL_1347 = _EVAL_234 ? 1'h0 : _EVAL_2691;
  assign _EVAL_797 = 9'hf1 == _EVAL_1399;
  assign _EVAL_2299 = 9'h85 == _EVAL_1399 ? 32'h0 : _EVAL_152;
  assign _EVAL_248 = 9'hfe == _EVAL_1399;
  assign _EVAL_1095 = _EVAL_3502 | _EVAL_2756;
  assign _EVAL_2399 = 9'h124 == _EVAL_1399 ? _EVAL_374 : _EVAL_692;
  assign _EVAL_1410 = _EVAL_386 ? _EVAL_3031 : _EVAL_1710;
  assign _EVAL_1611 = _EVAL_2838 | _EVAL_3814;
  assign _EVAL_207 = 9'h1b8 == _EVAL_1399 ? _EVAL_374 : _EVAL_3520;
  assign _EVAL_1135 = _EVAL_3337 == 7'h20;
  assign _EVAL_3788 = 9'h1ff == _EVAL_1399 ? _EVAL_1856 : _EVAL_3148;
  assign _EVAL_3119 = _EVAL_115 | _EVAL_699;
  assign _EVAL_2103 = 9'h37 == _EVAL_1399;
  assign _EVAL_1472 = 9'h38 == _EVAL_1399;
  assign _EVAL_214 = _EVAL_984 | _EVAL_2479;
  assign _EVAL_1884 = _EVAL_2437 & _EVAL_1945;
  assign _EVAL_2458 = _EVAL_995[23:0];
  assign _EVAL_3604 = 9'h81 == _EVAL_1399 ? 32'h0 : _EVAL_2314;
  assign _EVAL_3302 = 9'h1fd == _EVAL_1399 ? _EVAL_374 : _EVAL_3002;
  assign _EVAL_696 = 9'h5a == _EVAL_1399;
  assign _EVAL_217 = _EVAL_3418 & _EVAL_1856;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_67 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_167 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_266 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_351 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_555 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_819 = _RAND_5[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_1778 = _RAND_6[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_1805 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_1894 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_1987 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_2012 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_2218 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_2720 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_2757 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_2905 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_2978 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_2987 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_3000 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_3050 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_3066 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_3105 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_3138 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_3348 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_3402 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_3433 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_3777 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  if (_EVAL_3065) begin
    _EVAL_3066 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL) begin
    if (_EVAL_3425) begin
      _EVAL_67 <= 8'h0;
    end else if (_EVAL_3795) begin
      _EVAL_67 <= _EVAL_2763;
    end
    if (_EVAL_3425) begin
      _EVAL_167 <= 16'h0;
    end else if (_EVAL_3417) begin
      _EVAL_167 <= _EVAL_1978;
    end
    if (_EVAL_3425) begin
      _EVAL_266 <= 8'h0;
    end else if (_EVAL_474) begin
      _EVAL_266 <= _EVAL_3113;
    end else if (_EVAL_1540) begin
      if (_EVAL_2651) begin
        _EVAL_266 <= _EVAL_3143;
      end
    end
    if (_EVAL_3425) begin
      _EVAL_351 <= 8'h0;
    end else if (_EVAL_1049) begin
      _EVAL_351 <= _EVAL_3244;
    end else if (_EVAL_1881) begin
      if (_EVAL_2845) begin
        _EVAL_351 <= _EVAL_3102;
      end
    end
    if (_EVAL_3425) begin
      _EVAL_555 <= 8'h0;
    end else if (_EVAL_1871) begin
      _EVAL_555 <= _EVAL_3244;
    end else if (_EVAL_1869) begin
      if (_EVAL_2018) begin
        _EVAL_555 <= _EVAL_3102;
      end
    end
    if (_EVAL_3425) begin
      _EVAL_819 <= 24'h0;
    end else if (_EVAL_3795) begin
      _EVAL_819 <= _EVAL_2458;
    end
    if (_EVAL_3425) begin
      _EVAL_1778 <= 12'h0;
    end else if (_EVAL_2996) begin
      _EVAL_1778 <= _EVAL_2254;
    end
    if (_EVAL_3425) begin
      _EVAL_1805 <= 8'h0;
    end else if (_EVAL_3264) begin
      _EVAL_1805 <= _EVAL_2711;
    end else if (_EVAL_2183) begin
      if (_EVAL_1183) begin
        _EVAL_1805 <= _EVAL_2261;
      end
    end
    if (_EVAL_3425) begin
      _EVAL_1894 <= 8'h0;
    end else if (_EVAL_1376) begin
      _EVAL_1894 <= _EVAL_2711;
    end else if (_EVAL_2051) begin
      if (_EVAL_926) begin
        _EVAL_1894 <= _EVAL_2261;
      end
    end
    if (_EVAL_3425) begin
      _EVAL_1987 <= 2'h0;
    end else if (_EVAL_234) begin
      if (_EVAL_1437) begin
        _EVAL_1987 <= 2'h1;
      end
    end else if (_EVAL_421) begin
      if (_EVAL_3395) begin
        _EVAL_1987 <= 2'h0;
      end else if (_EVAL_1228) begin
        _EVAL_1987 <= 2'h0;
      end else begin
        _EVAL_1987 <= 2'h2;
      end
    end else if (_EVAL_470) begin
      if (_EVAL_2400) begin
        _EVAL_1987 <= 2'h0;
      end else if (_EVAL_406) begin
        _EVAL_1987 <= 2'h0;
      end
    end
    if (_EVAL_3425) begin
      _EVAL_2012 <= 3'h0;
    end else if (_EVAL_2021) begin
      _EVAL_2012 <= 3'h1;
    end else if (_EVAL_1347) begin
      _EVAL_2012 <= 3'h3;
    end else if (_EVAL_808) begin
      _EVAL_2012 <= 3'h2;
    end else if (_EVAL_1050) begin
      _EVAL_2012 <= 3'h4;
    end else if (_EVAL_1215) begin
      _EVAL_2012 <= _EVAL_2861;
    end
    if (_EVAL_3425) begin
      _EVAL_2218 <= 1'h0;
    end else begin
      _EVAL_2218 <= _EVAL_3700;
    end
    if (_EVAL_3425) begin
      _EVAL_2720 <= 8'h0;
    end else if (_EVAL_1191) begin
      _EVAL_2720 <= _EVAL_2420;
    end else if (_EVAL_1460) begin
      if (_EVAL_209) begin
        _EVAL_2720 <= _EVAL_3390;
      end
    end
    if (_EVAL_3425) begin
      _EVAL_2757 <= 8'h0;
    end else if (_EVAL_2029) begin
      _EVAL_2757 <= _EVAL_2711;
    end else if (_EVAL_2746) begin
      if (_EVAL_2714) begin
        _EVAL_2757 <= _EVAL_2261;
      end
    end
    if (_EVAL_3425) begin
      _EVAL_2905 <= 8'h0;
    end else if (_EVAL_829) begin
      _EVAL_2905 <= _EVAL_3113;
    end else if (_EVAL_549) begin
      if (_EVAL_1589) begin
        _EVAL_2905 <= _EVAL_3143;
      end
    end
    if (_EVAL_3425) begin
      _EVAL_2978 <= 1'h0;
    end else begin
      _EVAL_2978 <= _EVAL_1185;
    end
    if (_EVAL_3425) begin
      _EVAL_2987 <= 1'h0;
    end else begin
      _EVAL_2987 <= _EVAL_403;
    end
    if (_EVAL_1681) begin
      if (_EVAL_616) begin
        _EVAL_3000 <= 32'h13;
      end else begin
        _EVAL_3000 <= 32'h100073;
      end
    end
    if (_EVAL_3425) begin
      _EVAL_3050 <= 8'h0;
    end else if (_EVAL_1830) begin
      _EVAL_3050 <= _EVAL_3244;
    end else if (_EVAL_139) begin
      if (_EVAL_200) begin
        _EVAL_3050 <= _EVAL_3102;
      end
    end
    if (_EVAL_3425) begin
      _EVAL_3105 <= 1'h0;
    end else if (_EVAL_1110) begin
      _EVAL_3105 <= 1'h0;
    end else begin
      _EVAL_3105 <= _EVAL_3641;
    end
    if (_EVAL_3425) begin
      _EVAL_3138 <= 8'h0;
    end else if (_EVAL_1400) begin
      _EVAL_3138 <= _EVAL_2420;
    end else if (_EVAL_1037) begin
      if (_EVAL_724) begin
        _EVAL_3138 <= _EVAL_3390;
      end
    end
    if (_EVAL_1681) begin
      if (_EVAL_1562) begin
        if (_EVAL_230) begin
          _EVAL_3348 <= _EVAL_1401;
        end else begin
          _EVAL_3348 <= _EVAL_1842;
        end
      end else begin
        _EVAL_3348 <= 32'h13;
      end
    end
    if (_EVAL_38) begin
      _EVAL_3402 <= 1'h0;
    end else if (_EVAL_3425) begin
      _EVAL_3402 <= 1'h0;
    end else if (_EVAL_3203) begin
      _EVAL_3402 <= _EVAL_12;
    end
    if (_EVAL_3425) begin
      _EVAL_3433 <= 8'h0;
    end else if (_EVAL_1761) begin
      _EVAL_3433 <= _EVAL_2420;
    end else if (_EVAL_366) begin
      if (_EVAL_2828) begin
        _EVAL_3433 <= _EVAL_3390;
      end
    end
    if (_EVAL_3425) begin
      _EVAL_3777 <= 8'h0;
    end else if (_EVAL_3701) begin
      _EVAL_3777 <= _EVAL_3113;
    end else if (_EVAL_3824) begin
      if (_EVAL_2988) begin
        _EVAL_3777 <= _EVAL_3143;
      end
    end
  end
  always @(posedge _EVAL or posedge _EVAL_3065) begin
    if (_EVAL_3065) begin
      _EVAL_3066 <= 1'h0;
    end else if (_EVAL_3425) begin
      _EVAL_3066 <= 1'h0;
    end else begin
      _EVAL_3066 <= _EVAL_113;
    end
  end
endmodule
