//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_25_assert(
  input  [2:0]  _EVAL,
  input  [30:0] _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [2:0]  _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [1:0]  _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [3:0]  _EVAL_17,
  input         _EVAL_18
);
  wire  _EVAL_19;
  wire [4:0] _EVAL_20;
  wire  _EVAL_21;
  wire [3:0] _EVAL_22;
  wire [4:0] _EVAL_23;
  wire [5:0] _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire [7:0] _EVAL_39;
  wire  _EVAL_41;
  wire [4:0] _EVAL_42;
  wire [3:0] _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  reg  _EVAL_46;
  reg [31:0] _RAND_0;
  wire [4:0] _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire [3:0] _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_72;
  wire [1:0] _EVAL_73;
  wire [4:0] _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire [1:0] _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire [12:0] _EVAL_89;
  wire [32:0] _EVAL_90;
  reg [2:0] _EVAL_91;
  reg [31:0] _RAND_1;
  wire  _EVAL_93;
  wire  _EVAL_94;
  reg [31:0] _EVAL_95;
  reg [31:0] _RAND_2;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire [12:0] _EVAL_102;
  wire [3:0] _EVAL_103;
  wire [7:0] _EVAL_104;
  wire  _EVAL_105;
  wire [4:0] _EVAL_106;
  wire [31:0] _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  reg [1:0] _EVAL_117;
  reg [31:0] _RAND_3;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire [3:0] _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire [31:0] _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire [4:0] _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  reg  _EVAL_149;
  reg [31:0] _RAND_4;
  wire [3:0] _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_159;
  wire [1:0] _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  reg [3:0] _EVAL_169;
  reg [31:0] _RAND_5;
  reg [2:0] _EVAL_170;
  reg [31:0] _RAND_6;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  reg [2:0] _EVAL_185;
  reg [31:0] _RAND_7;
  wire  _EVAL_186;
  wire [4:0] _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  reg [3:0] _EVAL_190;
  reg [31:0] _RAND_8;
  wire [30:0] _EVAL_191;
  wire  _EVAL_192;
  wire [7:0] _EVAL_193;
  reg [2:0] _EVAL_194;
  reg [31:0] _RAND_9;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire [4:0] _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire [1:0] _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire [4:0] _EVAL_214;
  wire  _EVAL_215;
  reg [3:0] _EVAL_216;
  reg [31:0] _RAND_10;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire [31:0] _EVAL_219;
  wire  _EVAL_220;
  wire [4:0] _EVAL_221;
  wire [5:0] _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire [30:0] _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire [3:0] _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  reg [30:0] _EVAL_247;
  reg [31:0] _RAND_11;
  wire [31:0] _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  reg [2:0] _EVAL_251;
  reg [31:0] _RAND_12;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  reg [3:0] _EVAL_256;
  reg [31:0] _RAND_13;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire [3:0] _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire [5:0] _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  reg [4:0] _EVAL_272;
  reg [31:0] _RAND_14;
  wire [7:0] _EVAL_273;
  wire  _EVAL_274;
  wire [3:0] _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire [3:0] _EVAL_279;
  wire  _EVAL_280;
  wire [4:0] _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  reg [2:0] _EVAL_285;
  reg [31:0] _RAND_15;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_289;
  wire [30:0] _EVAL_290;
  wire [5:0] _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  reg [2:0] _EVAL_295;
  reg [31:0] _RAND_16;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_252 = _EVAL_37 | _EVAL_1;
  assign _EVAL_105 = _EVAL_83 == 2'h1;
  assign _EVAL_161 = 2'h1 << _EVAL_85;
  assign _EVAL_48 = _EVAL_10 & _EVAL_67;
  assign _EVAL_278 = _EVAL_141 | _EVAL_1;
  assign _EVAL_77 = ~_EVAL_36;
  assign _EVAL_174 = _EVAL_103 == 4'h0;
  assign _EVAL_162 = _EVAL_56 | _EVAL_1;
  assign _EVAL_186 = ~_EVAL_101;
  assign _EVAL_78 = _EVAL_10 & _EVAL_98;
  assign _EVAL_99 = _EVAL_246 & _EVAL_274;
  assign _EVAL_63 = _EVAL_289 & _EVAL_120;
  assign _EVAL_54 = _EVAL_5 == 3'h7;
  assign _EVAL_277 = _EVAL_217 | _EVAL_79;
  assign _EVAL_235 = _EVAL_136 | _EVAL_1;
  assign _EVAL_47 = _EVAL_272 >> _EVAL_12;
  assign _EVAL_233 = _EVAL_8 <= 3'h6;
  assign _EVAL_181 = _EVAL_210 | _EVAL_1;
  assign _EVAL_89 = 13'h3f << _EVAL_8;
  assign _EVAL_208 = _EVAL_179 | _EVAL_230;
  assign _EVAL_72 = _EVAL_31 & _EVAL_120;
  assign _EVAL_215 = ~_EVAL_270;
  assign _EVAL_144 = _EVAL_83 == 2'h0;
  assign _EVAL_177 = _EVAL_61 | _EVAL_1;
  assign _EVAL_56 = _EVAL_7 <= 3'h4;
  assign _EVAL_132 = _EVAL_13 != 2'h2;
  assign _EVAL_182 = ~_EVAL_165;
  assign _EVAL_204 = _EVAL_23 != 5'h0;
  assign _EVAL_238 = _EVAL_0 == _EVAL_247;
  assign _EVAL_236 = _EVAL_217 | _EVAL_231;
  assign _EVAL_52 = _EVAL_3 == _EVAL_295;
  assign _EVAL_33 = _EVAL_232 == 31'h0;
  assign _EVAL_96 = _EVAL_8 == _EVAL_170;
  assign _EVAL_41 = ~_EVAL_234;
  assign _EVAL_129 = _EVAL_13 == 2'h0;
  assign _EVAL_283 = ~_EVAL_119;
  assign _EVAL_232 = _EVAL_0 & _EVAL_191;
  assign _EVAL_192 = _EVAL_5 == 3'h0;
  assign _EVAL_22 = _EVAL_74[3:0];
  assign _EVAL_196 = _EVAL_130 | _EVAL_1;
  assign _EVAL_118 = _EVAL_53 & _EVAL_41;
  assign _EVAL_254 = ~_EVAL_57;
  assign _EVAL_290 = _EVAL_0 ^ 31'h40000000;
  assign _EVAL_38 = ~_EVAL_278;
  assign _EVAL_279 = _EVAL_17 & _EVAL_122;
  assign _EVAL_44 = ~_EVAL_120;
  assign _EVAL_79 = _EVAL_125 & _EVAL_63;
  assign _EVAL_23 = _EVAL_273[4:0];
  assign _EVAL_253 = _EVAL_166 | _EVAL_1;
  assign _EVAL_219 = _EVAL_90[31:0];
  assign _EVAL_116 = _EVAL_5 == 3'h3;
  assign _EVAL_115 = _EVAL_88 | _EVAL_1;
  assign _EVAL_66 = ~_EVAL_181;
  assign _EVAL_126 = _EVAL_11 & _EVAL_60;
  assign _EVAL_159 = _EVAL_195 | _EVAL_65;
  assign _EVAL_61 = _EVAL_142 | _EVAL_18;
  assign _EVAL_39 = _EVAL_118 ? _EVAL_193 : 8'h0;
  assign _EVAL_234 = _EVAL == 3'h6;
  assign _EVAL_101 = _EVAL_258 | _EVAL_1;
  assign _EVAL_195 = ~_EVAL_172;
  assign _EVAL_193 = 8'h1 << _EVAL_2;
  assign _EVAL_291 = _EVAL_102[5:0];
  assign _EVAL_228 = ~_EVAL_197;
  assign _EVAL_29 = _EVAL_105 | _EVAL_144;
  assign _EVAL_262 = _EVAL_218 | _EVAL_1;
  assign _EVAL_263 = ~_EVAL_222;
  assign _EVAL_237 = _EVAL_15 == _EVAL_149;
  assign _EVAL_135 = _EVAL_7 == 3'h0;
  assign _EVAL_100 = _EVAL_289 & _EVAL_44;
  assign _EVAL_87 = ~_EVAL_18;
  assign _EVAL_119 = _EVAL_52 | _EVAL_1;
  assign _EVAL_258 = _EVAL_13 <= 2'h2;
  assign _EVAL_155 = _EVAL_87 | _EVAL_1;
  assign _EVAL_70 = _EVAL_110 & _EVAL_289;
  assign _EVAL_273 = _EVAL_99 ? _EVAL_104 : 8'h0;
  assign _EVAL_203 = _EVAL_5[2];
  assign _EVAL_242 = _EVAL_2 == _EVAL_285;
  assign _EVAL_211 = _EVAL_161 | 2'h1;
  assign _EVAL_120 = _EVAL_0[0];
  assign _EVAL_85 = _EVAL_8[0];
  assign _EVAL_213 = _EVAL_233 & _EVAL_124;
  assign _EVAL_59 = _EVAL_51 | _EVAL_1;
  assign _EVAL_224 = _EVAL_33 | _EVAL_1;
  assign _EVAL_84 = ~_EVAL_27;
  assign _EVAL_74 = _EVAL_256 - 4'h1;
  assign _EVAL_103 = ~_EVAL_17;
  assign _EVAL_167 = ~_EVAL_245;
  assign _EVAL_173 = _EVAL_11 & _EVAL_234;
  assign _EVAL_122 = ~_EVAL_150;
  assign _EVAL_223 = _EVAL == _EVAL_91;
  assign _EVAL_102 = 13'h3f << _EVAL_3;
  assign _EVAL_187 = _EVAL_216 - 4'h1;
  assign _EVAL_42 = _EVAL_169 - 4'h1;
  assign _EVAL_134 = _EVAL_157 | _EVAL_58;
  assign _EVAL_113 = _EVAL_5 == 3'h4;
  assign _EVAL_191 = {{25'd0}, _EVAL_263};
  assign _EVAL_250 = ~_EVAL_175;
  assign _EVAL_201 = _EVAL_190 - 4'h1;
  assign _EVAL_156 = _EVAL <= 3'h6;
  assign _EVAL_260 = ~_EVAL_220;
  assign _EVAL_176 = ~_EVAL_69;
  assign _EVAL_293 = ~_EVAL_252;
  assign _EVAL_64 = _EVAL_209 | _EVAL_1;
  assign _EVAL_292 = _EVAL_10 & _EVAL_54;
  assign _EVAL_276 = _EVAL_246 & _EVAL_45;
  assign _EVAL_75 = _EVAL_95 < plusarg_reader_out;
  assign _EVAL_280 = _EVAL_246 | _EVAL_243;
  assign _EVAL_82 = _EVAL_10 & _EVAL_121;
  assign _EVAL_217 = _EVAL_157 | _EVAL_70;
  assign _EVAL_225 = _EVAL_5 == 3'h6;
  assign _EVAL_20 = _EVAL_106 >> _EVAL_2;
  assign _EVAL_80 = _EVAL_208 | _EVAL_168;
  assign _EVAL_214 = _EVAL_282 & _EVAL_221;
  assign _EVAL_145 = _EVAL_39[4:0];
  assign _EVAL_68 = _EVAL_5 == 3'h1;
  assign _EVAL_184 = _EVAL_10 & _EVAL_116;
  assign _EVAL_123 = _EVAL_10 & _EVAL_225;
  assign _EVAL_261 = _EVAL_238 | _EVAL_1;
  assign _EVAL_65 = plusarg_reader_out == 32'h0;
  assign _EVAL_165 = _EVAL_35 | _EVAL_1;
  assign _EVAL_207 = ~_EVAL_177;
  assign _EVAL_265 = _EVAL_134 | _EVAL_81;
  assign _EVAL_245 = _EVAL_142 | _EVAL_1;
  assign _EVAL_175 = _EVAL_47[0];
  assign _EVAL_257 = _EVAL_7 <= 3'h2;
  assign _EVAL_267 = _EVAL == 3'h4;
  assign _EVAL_282 = _EVAL_272 | _EVAL_23;
  assign _EVAL_248 = _EVAL_107;
  assign _EVAL_172 = _EVAL_272 != 5'h0;
  assign _EVAL_209 = _EVAL_5 == _EVAL_251;
  assign _EVAL_50 = _EVAL == 3'h0;
  assign _EVAL_143 = _EVAL_243 & _EVAL_151;
  assign _EVAL_35 = ~_EVAL_16;
  assign _EVAL_55 = _EVAL_263[5:2];
  assign _EVAL_127 = _EVAL_157 | _EVAL_1;
  assign _EVAL_197 = _EVAL_199 | _EVAL_1;
  assign _EVAL_210 = _EVAL_14 == _EVAL_46;
  assign _EVAL_151 = _EVAL_169 == 4'h0;
  assign _EVAL_166 = _EVAL_159 | _EVAL_75;
  assign _EVAL_205 = ~_EVAL_146;
  assign _EVAL_124 = $signed(_EVAL_248) == 32'sh0;
  assign _EVAL_24 = ~_EVAL_291;
  assign _EVAL_229 = _EVAL_223 | _EVAL_1;
  assign _EVAL_154 = ~_EVAL_224;
  assign _EVAL_73 = _EVAL_12[2:1];
  assign _EVAL_286 = _EVAL_10 & _EVAL_192;
  assign _EVAL_147 = _EVAL_198 | _EVAL_21;
  assign _EVAL_163 = ~_EVAL_109;
  assign _EVAL_240 = ~_EVAL_229;
  assign _EVAL_128 = _EVAL[0];
  assign _EVAL_157 = _EVAL_8 >= 3'h2;
  assign _EVAL_121 = _EVAL_5 == 3'h5;
  assign _EVAL_241 = _EVAL_187[3:0];
  assign _EVAL_37 = _EVAL_29 | _EVAL_249;
  assign _EVAL_51 = _EVAL_7 <= 3'h1;
  assign _EVAL_106 = _EVAL_23 | _EVAL_272;
  assign _EVAL_255 = ~_EVAL_151;
  assign _EVAL_249 = _EVAL_2 == 3'h4;
  assign _EVAL_150 = {_EVAL_277,_EVAL_236,_EVAL_265,_EVAL_139};
  assign _EVAL_148 = ~_EVAL_200;
  assign _EVAL_179 = _EVAL_73 == 2'h1;
  assign _EVAL_62 = _EVAL_96 | _EVAL_1;
  assign _EVAL_58 = _EVAL_110 & _EVAL_31;
  assign _EVAL_81 = _EVAL_125 & _EVAL_72;
  assign _EVAL_137 = {1'b0,$signed(_EVAL_290)};
  assign _EVAL_26 = ~_EVAL_152;
  assign _EVAL_98 = _EVAL_5 == 3'h2;
  assign _EVAL_244 = ~_EVAL_138;
  assign _EVAL_183 = ~_EVAL_203;
  assign _EVAL_139 = _EVAL_134 | _EVAL_49;
  assign _EVAL_222 = _EVAL_89[5:0];
  assign _EVAL_69 = _EVAL_237 | _EVAL_1;
  assign _EVAL_202 = ~_EVAL_62;
  assign _EVAL_57 = _EVAL_80 | _EVAL_1;
  assign _EVAL_153 = _EVAL == 3'h2;
  assign _EVAL_28 = ~_EVAL_253;
  assign _EVAL_125 = _EVAL_211[0];
  assign _EVAL_133 = _EVAL_10 & _EVAL_68;
  assign _EVAL_138 = _EVAL_174 | _EVAL_1;
  assign _EVAL_53 = _EVAL_243 & _EVAL_271;
  assign _EVAL_86 = _EVAL_11 & _EVAL_19;
  assign _EVAL_270 = _EVAL_250 | _EVAL_1;
  assign _EVAL_94 = ~_EVAL_264;
  assign _EVAL_246 = _EVAL_6 & _EVAL_10;
  assign _EVAL_140 = _EVAL_7 != 3'h0;
  assign _EVAL_271 = _EVAL_190 == 4'h0;
  assign _EVAL_142 = ~_EVAL_14;
  assign _EVAL_93 = ~_EVAL_111;
  assign _EVAL_21 = ~_EVAL_204;
  assign _EVAL_231 = _EVAL_125 & _EVAL_100;
  assign _EVAL_141 = _EVAL_17 == _EVAL_150;
  assign _EVAL_32 = _EVAL_11 & _EVAL_50;
  assign _EVAL_111 = _EVAL_108 | _EVAL_1;
  assign _EVAL_67 = ~_EVAL_45;
  assign _EVAL_31 = ~_EVAL_289;
  assign _EVAL_188 = ~_EVAL_261;
  assign _EVAL_164 = ~_EVAL_127;
  assign _EVAL_275 = _EVAL_201[3:0];
  assign _EVAL_152 = _EVAL_257 | _EVAL_1;
  assign _EVAL_114 = ~_EVAL_162;
  assign _EVAL_83 = _EVAL_2[2:1];
  assign _EVAL_269 = _EVAL_11 & _EVAL_255;
  assign _EVAL_230 = _EVAL_73 == 2'h0;
  assign _EVAL_45 = _EVAL_216 == 4'h0;
  assign _EVAL_36 = _EVAL_213 | _EVAL_1;
  assign _EVAL_136 = _EVAL_279 == 4'h0;
  assign _EVAL_220 = _EVAL_147 | _EVAL_1;
  assign _EVAL_274 = _EVAL_256 == 4'h0;
  assign _EVAL_108 = _EVAL_7 <= 3'h3;
  assign _EVAL_287 = _EVAL_10 & _EVAL_113;
  assign _EVAL_221 = ~_EVAL_145;
  assign _EVAL_27 = _EVAL_129 | _EVAL_1;
  assign _EVAL_97 = ~_EVAL_196;
  assign _EVAL_206 = ~_EVAL_212;
  assign _EVAL_90 = _EVAL_95 + 32'h1;
  assign _EVAL_199 = _EVAL_20[0];
  assign _EVAL_107 = $signed(_EVAL_137) & -32'sh2000;
  assign _EVAL_112 = ~_EVAL_59;
  assign _EVAL_180 = ~_EVAL_115;
  assign _EVAL_294 = ~_EVAL_262;
  assign _EVAL_25 = ~_EVAL_131;
  assign _EVAL_168 = _EVAL_12 == 3'h4;
  assign _EVAL_239 = _EVAL_11 & _EVAL_267;
  assign _EVAL_200 = _EVAL_284 | _EVAL_1;
  assign _EVAL_49 = _EVAL_125 & _EVAL_189;
  assign _EVAL_266 = ~_EVAL_155;
  assign _EVAL_130 = _EVAL_3 >= 3'h2;
  assign _EVAL_189 = _EVAL_31 & _EVAL_44;
  assign _EVAL_43 = _EVAL_42[3:0];
  assign _EVAL_146 = _EVAL_140 | _EVAL_1;
  assign _EVAL_131 = _EVAL_156 | _EVAL_1;
  assign _EVAL_109 = _EVAL_132 | _EVAL_1;
  assign _EVAL_110 = _EVAL_211[1];
  assign _EVAL_284 = _EVAL_13 == _EVAL_117;
  assign _EVAL_34 = _EVAL_11 & _EVAL_153;
  assign _EVAL_243 = _EVAL_9 & _EVAL_11;
  assign _EVAL_88 = _EVAL_12 == _EVAL_194;
  assign _EVAL_268 = ~_EVAL_235;
  assign _EVAL_198 = _EVAL_23 != _EVAL_145;
  assign _EVAL_19 = _EVAL == 3'h5;
  assign _EVAL_212 = _EVAL_242 | _EVAL_1;
  assign _EVAL_227 = ~_EVAL_1;
  assign _EVAL_259 = _EVAL_24[5:2];
  assign _EVAL_218 = _EVAL_7 == _EVAL_185;
  assign _EVAL_264 = _EVAL_135 | _EVAL_1;
  assign _EVAL_178 = ~_EVAL_64;
  assign _EVAL_104 = 8'h1 << _EVAL_12;
  assign _EVAL_289 = _EVAL_0[1];
  assign _EVAL_60 = _EVAL == 3'h1;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_46 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_91 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_95 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_117 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_149 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_169 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_170 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_185 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_190 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_194 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_216 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_247 = _RAND_11[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_251 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_256 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_272 = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_285 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_295 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_4) begin
    if (_EVAL_143) begin
      _EVAL_46 <= _EVAL_14;
    end
    if (_EVAL_143) begin
      _EVAL_91 <= _EVAL;
    end
    if (_EVAL_1) begin
      _EVAL_95 <= 32'h0;
    end else if (_EVAL_280) begin
      _EVAL_95 <= 32'h0;
    end else begin
      _EVAL_95 <= _EVAL_219;
    end
    if (_EVAL_143) begin
      _EVAL_117 <= _EVAL_13;
    end
    if (_EVAL_143) begin
      _EVAL_149 <= _EVAL_15;
    end
    if (_EVAL_1) begin
      _EVAL_169 <= 4'h0;
    end else if (_EVAL_243) begin
      if (_EVAL_151) begin
        if (_EVAL_128) begin
          _EVAL_169 <= _EVAL_259;
        end else begin
          _EVAL_169 <= 4'h0;
        end
      end else begin
        _EVAL_169 <= _EVAL_43;
      end
    end
    if (_EVAL_276) begin
      _EVAL_170 <= _EVAL_8;
    end
    if (_EVAL_276) begin
      _EVAL_185 <= _EVAL_7;
    end
    if (_EVAL_1) begin
      _EVAL_190 <= 4'h0;
    end else if (_EVAL_243) begin
      if (_EVAL_271) begin
        if (_EVAL_128) begin
          _EVAL_190 <= _EVAL_259;
        end else begin
          _EVAL_190 <= 4'h0;
        end
      end else begin
        _EVAL_190 <= _EVAL_275;
      end
    end
    if (_EVAL_276) begin
      _EVAL_194 <= _EVAL_12;
    end
    if (_EVAL_1) begin
      _EVAL_216 <= 4'h0;
    end else if (_EVAL_246) begin
      if (_EVAL_45) begin
        if (_EVAL_183) begin
          _EVAL_216 <= _EVAL_55;
        end else begin
          _EVAL_216 <= 4'h0;
        end
      end else begin
        _EVAL_216 <= _EVAL_241;
      end
    end
    if (_EVAL_276) begin
      _EVAL_247 <= _EVAL_0;
    end
    if (_EVAL_276) begin
      _EVAL_251 <= _EVAL_5;
    end
    if (_EVAL_1) begin
      _EVAL_256 <= 4'h0;
    end else if (_EVAL_246) begin
      if (_EVAL_274) begin
        if (_EVAL_183) begin
          _EVAL_256 <= _EVAL_55;
        end else begin
          _EVAL_256 <= 4'h0;
        end
      end else begin
        _EVAL_256 <= _EVAL_22;
      end
    end
    if (_EVAL_1) begin
      _EVAL_272 <= 5'h0;
    end else begin
      _EVAL_272 <= _EVAL_214;
    end
    if (_EVAL_143) begin
      _EVAL_285 <= _EVAL_2;
    end
    if (_EVAL_143) begin
      _EVAL_295 <= _EVAL_3;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d2fcae8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f731a641)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b848bd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b45e7ecd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d3e8929)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e05b7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f4bb00b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(881615a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3057aa6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5368afcb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56fd5752)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2658ee53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5504eb2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8818e591)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(643a8060)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d0b319a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bffdaca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17e3ee7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2797d7a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79808ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45ffb970)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa6623e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9921198)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1596d71e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0159ecf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdbc5cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(947e8384)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3183cec0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(456a8953)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d15d71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91277150)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fcf5c44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e9e6fc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_66) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a5170f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(feace9d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccdf4eee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7c27495)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f8ad5eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9ae872c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cf3a629)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bb5bb12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0ce27d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(697593cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f0e8c3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6197d9e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_66) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bc196e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49a5db30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed114575)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e1d648a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_294) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6eed72f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8a380b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_294) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa571a8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fae2013)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d11108a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce15ec2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56fb871d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80625db7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12f120)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b883bdff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b892417e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(956592c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d34aaab9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(820af394)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(600bd221)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7bf5969)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48f86f2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ab63fca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9f23fbc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6aac8835)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cd7d0c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bef25851)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9bfbef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a5d4de1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8260212a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8daed546)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19a5616c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29289122)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86546731)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70690027)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e8ae8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(679676c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d83b4d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5ca522c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f787914c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3769b33d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(377bdbda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13822e39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e386f58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(689f50d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc30db05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f00616ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e0adf3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a61e280c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
