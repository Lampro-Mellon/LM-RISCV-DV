//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_125_assert(
  input          _EVAL,
  input  [2:0]   _EVAL_0,
  input          _EVAL_1,
  input          _EVAL_2,
  input          _EVAL_3,
  input  [3:0]   _EVAL_4,
  input  [1:0]   _EVAL_5,
  input  [2:0]   _EVAL_6,
  input          _EVAL_7,
  input          _EVAL_8,
  input          _EVAL_9,
  input          _EVAL_10,
  input          _EVAL_11,
  input  [127:0] _EVAL_12,
  input          _EVAL_13,
  input  [1:0]   _EVAL_14
);
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  reg  _EVAL_27;
  reg [31:0] _RAND_0;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  reg  _EVAL_39;
  reg [31:0] _RAND_1;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire [1:0] _EVAL_45;
  wire  _EVAL_46;
  reg [2:0] _EVAL_47;
  reg [31:0] _RAND_2;
  wire [1:0] _EVAL_48;
  wire  _EVAL_49;
  wire [1:0] _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire [32:0] _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  reg [127:0] _EVAL_61;
  reg [127:0] _RAND_3;
  wire  _EVAL_63;
  reg  _EVAL_64;
  reg [31:0] _RAND_4;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  reg  _EVAL_71;
  reg [31:0] _RAND_5;
  wire  _EVAL_72;
  reg  _EVAL_73;
  reg [31:0] _RAND_6;
  wire  _EVAL_74;
  wire [127:0] _EVAL_75;
  reg  _EVAL_76;
  reg [31:0] _RAND_7;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire [128:0] _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  reg [31:0] _EVAL_85;
  reg [31:0] _RAND_8;
  wire [1:0] _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  reg [2:0] _EVAL_90;
  reg [31:0] _RAND_9;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire [128:0] _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire [1:0] _EVAL_98;
  wire  _EVAL_99;
  wire [128:0] _EVAL_100;
  wire  _EVAL_101;
  wire [1:0] _EVAL_102;
  wire  _EVAL_103;
  wire [31:0] _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  reg  _EVAL_119;
  reg [31:0] _RAND_10;
  reg [1:0] _EVAL_120;
  reg [31:0] _RAND_11;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  reg [1:0] _EVAL_124;
  reg [31:0] _RAND_12;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire [3:0] _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  reg  _EVAL_169;
  reg [31:0] _RAND_13;
  wire  _EVAL_170;
  wire [1:0] _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_179 = _EVAL_142 | _EVAL_92;
  assign _EVAL_35 = _EVAL_8 & _EVAL_141;
  assign _EVAL_102 = _EVAL_73 - 1'h1;
  assign _EVAL_31 = _EVAL_45[0];
  assign _EVAL_53 = _EVAL_5 == _EVAL_124;
  assign _EVAL_37 = _EVAL_143 | _EVAL_92;
  assign _EVAL_129 = ~_EVAL_92;
  assign _EVAL_15 = _EVAL_98[0];
  assign _EVAL_165 = ~_EVAL_95;
  assign _EVAL_148 = _EVAL_164 | _EVAL_92;
  assign _EVAL_161 = _EVAL_80 | _EVAL_92;
  assign _EVAL_130 = _EVAL_89 & _EVAL_133;
  assign _EVAL_141 = _EVAL_6 == 3'h7;
  assign _EVAL_172 = _EVAL_4 == 4'hf;
  assign _EVAL_147 = _EVAL_72 | _EVAL_92;
  assign _EVAL_139 = _EVAL_15 | _EVAL_169;
  assign _EVAL_48 = _EVAL_119 - 1'h1;
  assign _EVAL_115 = ~_EVAL_73;
  assign _EVAL_25 = _EVAL_8 & _EVAL_16;
  assign _EVAL_121 = ~_EVAL_28;
  assign _EVAL_142 = ~_EVAL_13;
  assign _EVAL_88 = _EVAL_7 & _EVAL_59;
  assign _EVAL_24 = _EVAL_175 | _EVAL_92;
  assign _EVAL_104 = _EVAL_57[31:0];
  assign _EVAL_59 = ~_EVAL_133;
  assign _EVAL_178 = _EVAL_6 == 3'h4;
  assign _EVAL_30 = ~_EVAL_43;
  assign _EVAL_97 = _EVAL_159 | _EVAL_92;
  assign _EVAL_52 = _EVAL_14 <= 2'h2;
  assign _EVAL_145 = _EVAL_8 & _EVAL_178;
  assign _EVAL_81 = _EVAL_100;
  assign _EVAL_92 = _EVAL_1;
  assign _EVAL_44 = _EVAL_69 | _EVAL_107;
  assign _EVAL_103 = _EVAL_7 & _EVAL_19;
  assign _EVAL_158 = _EVAL_8 & _EVAL_55;
  assign _EVAL_177 = _EVAL_160 | _EVAL_92;
  assign _EVAL_114 = _EVAL_8 & _EVAL_146;
  assign _EVAL_168 = _EVAL_7 & _EVAL_132;
  assign _EVAL_111 = _EVAL_22 | _EVAL_92;
  assign _EVAL_173 = _EVAL_6 == 3'h1;
  assign _EVAL_67 = _EVAL_50[0];
  assign _EVAL_176 = _EVAL_75 == 128'h0;
  assign _EVAL_122 = _EVAL_7 & _EVAL_101;
  assign _EVAL_63 = _EVAL_8 & _EVAL_56;
  assign _EVAL_50 = _EVAL_135 ? _EVAL_171 : 2'h0;
  assign _EVAL_79 = _EVAL_86[0];
  assign _EVAL_74 = _EVAL_53 | _EVAL_92;
  assign _EVAL_171 = 2'h1 << _EVAL_13;
  assign _EVAL_70 = ~_EVAL_153;
  assign _EVAL_43 = _EVAL_20 | _EVAL_92;
  assign _EVAL_36 = ~_EVAL_67;
  assign _EVAL_17 = _EVAL_0 == 3'h6;
  assign _EVAL_136 = _EVAL_172 | _EVAL_92;
  assign _EVAL_41 = _EVAL_0 == 3'h1;
  assign _EVAL_57 = _EVAL_85 + 32'h1;
  assign _EVAL_125 = ~_EVAL_163;
  assign _EVAL_100 = $signed(_EVAL_93) & -129'sh100000000000000000000000000000000;
  assign _EVAL_137 = _EVAL_139 >> _EVAL_13;
  assign _EVAL_54 = _EVAL_5 >= 2'h2;
  assign _EVAL_166 = ~_EVAL_4;
  assign _EVAL_164 = _EVAL_44 | _EVAL_23;
  assign _EVAL_55 = _EVAL_6 == 3'h2;
  assign _EVAL_69 = ~_EVAL_169;
  assign _EVAL_91 = ~_EVAL_74;
  assign _EVAL_117 = _EVAL_169 | _EVAL_15;
  assign _EVAL_72 = _EVAL_12 == _EVAL_61;
  assign _EVAL_95 = _EVAL_137 | _EVAL_92;
  assign _EVAL_144 = _EVAL_0 <= 3'h6;
  assign _EVAL_170 = _EVAL_7 & _EVAL_17;
  assign _EVAL_29 = _EVAL_8 & _EVAL_113;
  assign _EVAL_116 = _EVAL_54 | _EVAL_92;
  assign _EVAL_157 = ~_EVAL_33;
  assign _EVAL_127 = _EVAL_105 | _EVAL_92;
  assign _EVAL_49 = ~_EVAL_161;
  assign _EVAL_146 = _EVAL_6 == 3'h0;
  assign _EVAL_94 = _EVAL_42 | _EVAL_92;
  assign _EVAL_26 = _EVAL_131 | _EVAL_92;
  assign _EVAL_101 = _EVAL_0 == 3'h2;
  assign _EVAL_159 = _EVAL_6 == _EVAL_47;
  assign _EVAL_135 = _EVAL_40 & _EVAL_38;
  assign _EVAL_38 = ~_EVAL_17;
  assign _EVAL_160 = _EVAL_11 == _EVAL_27;
  assign _EVAL_154 = _EVAL_176 | _EVAL_92;
  assign _EVAL_34 = _EVAL_8 & _EVAL_65;
  assign _EVAL_19 = _EVAL_0 == 3'h5;
  assign _EVAL_89 = _EVAL & _EVAL_7;
  assign _EVAL_80 = _EVAL_14 == _EVAL_120;
  assign _EVAL_22 = $signed(_EVAL_81) == 129'sh0;
  assign _EVAL_66 = ~_EVAL_46;
  assign _EVAL_110 = ~_EVAL_136;
  assign _EVAL_131 = _EVAL_2 == _EVAL_64;
  assign _EVAL_162 = ~_EVAL_154;
  assign _EVAL_132 = _EVAL_0 == 3'h0;
  assign _EVAL_33 = _EVAL_69 | _EVAL_92;
  assign _EVAL_18 = _EVAL_102[0];
  assign _EVAL_105 = ~_EVAL_10;
  assign _EVAL_155 = _EVAL_84 & _EVAL_152;
  assign _EVAL_108 = _EVAL_7 & _EVAL_78;
  assign _EVAL_99 = ~_EVAL_150;
  assign _EVAL_112 = ~_EVAL_96;
  assign _EVAL_87 = ~_EVAL_97;
  assign _EVAL_163 = _EVAL_140 | _EVAL_92;
  assign _EVAL_77 = ~_EVAL_37;
  assign _EVAL_128 = ~_EVAL_179;
  assign _EVAL_16 = _EVAL_6 == 3'h3;
  assign _EVAL_84 = _EVAL_3 & _EVAL_8;
  assign _EVAL_58 = _EVAL_48[0];
  assign _EVAL_118 = ~_EVAL_71;
  assign _EVAL_152 = ~_EVAL_119;
  assign _EVAL_156 = _EVAL_8 & _EVAL_173;
  assign _EVAL_83 = ~_EVAL_147;
  assign _EVAL_82 = ~_EVAL_127;
  assign _EVAL_21 = _EVAL_2 < 1'h1;
  assign _EVAL_109 = ~_EVAL_111;
  assign _EVAL_150 = _EVAL_106 | _EVAL_92;
  assign _EVAL_133 = ~_EVAL_76;
  assign _EVAL_149 = _EVAL_84 | _EVAL_89;
  assign _EVAL_32 = ~_EVAL_177;
  assign _EVAL_93 = {1'b0,$signed(_EVAL_12)};
  assign _EVAL_106 = _EVAL_166 == 4'h0;
  assign _EVAL_45 = _EVAL_76 - 1'h1;
  assign _EVAL_175 = _EVAL_13 == _EVAL_39;
  assign _EVAL_98 = _EVAL_155 ? 2'h1 : 2'h0;
  assign _EVAL_56 = ~_EVAL_115;
  assign _EVAL_96 = _EVAL_51 | _EVAL_92;
  assign _EVAL_113 = _EVAL_6 == 3'h6;
  assign _EVAL_78 = _EVAL_0 == 3'h4;
  assign _EVAL_20 = ~_EVAL_11;
  assign _EVAL_140 = _EVAL_0 == _EVAL_90;
  assign _EVAL_126 = _EVAL_84 & _EVAL_115;
  assign _EVAL_28 = _EVAL_144 | _EVAL_92;
  assign _EVAL_46 = _EVAL_21 | _EVAL_92;
  assign _EVAL_23 = _EVAL_85 < plusarg_reader_out;
  assign _EVAL_153 = _EVAL_52 | _EVAL_92;
  assign _EVAL_174 = ~_EVAL_26;
  assign _EVAL_40 = _EVAL_89 & _EVAL_118;
  assign _EVAL_75 = _EVAL_12 & 128'h3;
  assign _EVAL_60 = ~_EVAL_94;
  assign _EVAL_143 = _EVAL_14 != 2'h2;
  assign _EVAL_167 = ~_EVAL_148;
  assign _EVAL_123 = ~_EVAL_116;
  assign _EVAL_68 = _EVAL_7 & _EVAL_41;
  assign _EVAL_107 = plusarg_reader_out == 32'h0;
  assign _EVAL_86 = _EVAL_71 - 1'h1;
  assign _EVAL_42 = _EVAL_14 == 2'h0;
  assign _EVAL_51 = _EVAL_20 | _EVAL_10;
  assign _EVAL_65 = _EVAL_6 == 3'h5;
  assign _EVAL_138 = ~_EVAL_24;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_27 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_39 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_47 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {4{`RANDOM}};
  _EVAL_61 = _RAND_3[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_64 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_71 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_73 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_76 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_85 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_90 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_119 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_120 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_124 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_169 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  if (_EVAL_1) begin
    _EVAL_71 = 1'h0;
  end
  if (_EVAL_1) begin
    _EVAL_73 = 1'h0;
  end
  if (_EVAL_1) begin
    _EVAL_76 = 1'h0;
  end
  if (_EVAL_1) begin
    _EVAL_85 = 32'h0;
  end
  if (_EVAL_1) begin
    _EVAL_119 = 1'h0;
  end
  if (_EVAL_1) begin
    _EVAL_169 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_9) begin
    if (_EVAL_130) begin
      _EVAL_27 <= _EVAL_11;
    end
    if (_EVAL_130) begin
      _EVAL_39 <= _EVAL_13;
    end
    if (_EVAL_126) begin
      _EVAL_47 <= _EVAL_6;
    end
    if (_EVAL_126) begin
      _EVAL_61 <= _EVAL_12;
    end
    if (_EVAL_130) begin
      _EVAL_64 <= _EVAL_2;
    end
    if (_EVAL_130) begin
      _EVAL_90 <= _EVAL_0;
    end
    if (_EVAL_130) begin
      _EVAL_120 <= _EVAL_14;
    end
    if (_EVAL_130) begin
      _EVAL_124 <= _EVAL_5;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5a81e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_66) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7bb6960)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5355497f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c235be2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dbf053e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88d83a88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fee0369)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c34f92b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e46f215f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cdc4642)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d6e2081)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4775be1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4d4c038)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af314b42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eab52114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15ce0d44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be10a63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(524413da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6d84cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4343277)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c248592f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62f38a60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eeaa93bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e3f9763)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56e72a8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32f9eca1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b0869c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(427ef5ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f4c81c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7913d73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdcd54b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(722da240)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e387ad4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1315c67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faee49e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bc0ac66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93539acc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f57c7bea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56c8f0e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2262996)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b78916a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd7a5ca6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d9538f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(763d2a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_66) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cda668dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(726c8dcb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ccf3b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14667850)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e722e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c58712d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_66) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf2b0580)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38ebbf05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fc74b63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_66) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42697acb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9848e74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad418d13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dbbed6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(618034f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4d9ca85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5c6bdb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fe42ce9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3245f2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(377acc4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6e6e4f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge _EVAL_9 or posedge _EVAL_1) begin
    if (_EVAL_1) begin
      _EVAL_71 <= 1'h0;
    end else if (_EVAL_89) begin
      if (_EVAL_118) begin
        _EVAL_71 <= 1'h0;
      end else begin
        _EVAL_71 <= _EVAL_79;
      end
    end
  end
  always @(posedge _EVAL_9 or posedge _EVAL_1) begin
    if (_EVAL_1) begin
      _EVAL_73 <= 1'h0;
    end else if (_EVAL_84) begin
      if (_EVAL_115) begin
        _EVAL_73 <= 1'h0;
      end else begin
        _EVAL_73 <= _EVAL_18;
      end
    end
  end
  always @(posedge _EVAL_9 or posedge _EVAL_1) begin
    if (_EVAL_1) begin
      _EVAL_76 <= 1'h0;
    end else if (_EVAL_89) begin
      if (_EVAL_133) begin
        _EVAL_76 <= 1'h0;
      end else begin
        _EVAL_76 <= _EVAL_31;
      end
    end
  end
  always @(posedge _EVAL_9 or posedge _EVAL_1) begin
    if (_EVAL_1) begin
      _EVAL_85 <= 32'h0;
    end else if (_EVAL_149) begin
      _EVAL_85 <= 32'h0;
    end else begin
      _EVAL_85 <= _EVAL_104;
    end
  end
  always @(posedge _EVAL_9 or posedge _EVAL_1) begin
    if (_EVAL_1) begin
      _EVAL_119 <= 1'h0;
    end else if (_EVAL_84) begin
      if (_EVAL_152) begin
        _EVAL_119 <= 1'h0;
      end else begin
        _EVAL_119 <= _EVAL_58;
      end
    end
  end
  always @(posedge _EVAL_9 or posedge _EVAL_1) begin
    if (_EVAL_1) begin
      _EVAL_169 <= 1'h0;
    end else begin
      _EVAL_169 <= _EVAL_117 & _EVAL_36;
    end
  end

endmodule
