//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_148(
  output        _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [11:0] _EVAL_4,
  output        _EVAL_5,
  output        _EVAL_6,
  output        _EVAL_7,
  output [2:0]  _EVAL_8,
  output [31:0] _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  output        _EVAL_12,
  input  [31:0] _EVAL_13,
  input         _EVAL_14,
  input  [3:0]  _EVAL_15,
  output        _EVAL_16,
  input  [3:0]  _EVAL_17,
  input  [2:0]  _EVAL_18,
  input  [31:0] _EVAL_19,
  input         _EVAL_20,
  output [31:0] _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  output [1:0]  _EVAL_24,
  input  [2:0]  _EVAL_25,
  output [2:0]  _EVAL_26,
  input  [8:0]  _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  output [1:0]  _EVAL_30,
  input         _EVAL_31,
  input  [2:0]  _EVAL_32,
  input         _EVAL_33,
  output        _EVAL_34,
  input  [1:0]  _EVAL_35,
  output [2:0]  _EVAL_36
);
  wire  AsyncQueueSink__EVAL;
  wire  AsyncQueueSink__EVAL_0;
  wire  AsyncQueueSink__EVAL_1;
  wire  AsyncQueueSink__EVAL_2;
  wire  AsyncQueueSink__EVAL_3;
  wire  AsyncQueueSink__EVAL_4;
  wire  AsyncQueueSink__EVAL_5;
  wire  AsyncQueueSink__EVAL_6;
  wire  AsyncQueueSink__EVAL_7;
  wire  AsyncQueueSink__EVAL_8;
  wire [9:0] AsyncQueueSink__EVAL_9;
  wire  AsyncQueueSink__EVAL_10;
  wire  dmactiveSync__EVAL;
  wire  dmactiveSync__EVAL_0;
  wire  dmactiveSync__EVAL_1;
  wire  dmactiveSync__EVAL_2;
  wire [1:0] dmiXing__EVAL;
  wire [2:0] dmiXing__EVAL_0;
  wire  dmiXing__EVAL_1;
  wire  dmiXing__EVAL_2;
  wire  dmiXing__EVAL_3;
  wire [31:0] dmiXing__EVAL_4;
  wire [2:0] dmiXing__EVAL_5;
  wire [3:0] dmiXing__EVAL_6;
  wire  dmiXing__EVAL_7;
  wire [2:0] dmiXing__EVAL_8;
  wire  dmiXing__EVAL_9;
  wire  dmiXing__EVAL_10;
  wire [1:0] dmiXing__EVAL_11;
  wire [2:0] dmiXing__EVAL_12;
  wire  dmiXing__EVAL_13;
  wire  dmiXing__EVAL_14;
  wire  dmiXing__EVAL_15;
  wire  dmiXing__EVAL_16;
  wire [8:0] dmiXing__EVAL_17;
  wire [1:0] dmiXing__EVAL_18;
  wire [8:0] dmiXing__EVAL_19;
  wire  dmiXing__EVAL_20;
  wire [31:0] dmiXing__EVAL_21;
  wire  dmiXing__EVAL_22;
  wire  dmiXing__EVAL_23;
  wire [31:0] dmiXing__EVAL_24;
  wire [2:0] dmiXing__EVAL_25;
  wire  dmiXing__EVAL_26;
  wire [31:0] dmiXing__EVAL_27;
  wire [3:0] dmiXing__EVAL_28;
  wire  dmInner__EVAL;
  wire [2:0] dmInner__EVAL_0;
  wire [1:0] dmInner__EVAL_1;
  wire  dmInner__EVAL_2;
  wire [9:0] dmInner__EVAL_3;
  wire [2:0] dmInner__EVAL_4;
  wire [2:0] dmInner__EVAL_5;
  wire  dmInner__EVAL_6;
  wire  dmInner__EVAL_7;
  wire  dmInner__EVAL_8;
  wire [31:0] dmInner__EVAL_9;
  wire [31:0] dmInner__EVAL_10;
  wire [31:0] dmInner__EVAL_11;
  wire  dmInner__EVAL_12;
  wire [2:0] dmInner__EVAL_13;
  wire [1:0] dmInner__EVAL_14;
  wire [2:0] dmInner__EVAL_15;
  wire  dmInner__EVAL_16;
  wire  dmInner__EVAL_17;
  wire  dmInner__EVAL_18;
  wire  dmInner__EVAL_19;
  wire  dmInner__EVAL_20;
  wire [8:0] dmInner__EVAL_21;
  wire  dmInner__EVAL_22;
  wire [1:0] dmInner__EVAL_23;
  wire [2:0] dmInner__EVAL_24;
  wire  dmInner__EVAL_25;
  wire [31:0] dmInner__EVAL_26;
  wire  dmInner__EVAL_27;
  wire [3:0] dmInner__EVAL_28;
  wire [3:0] dmInner__EVAL_29;
  wire  dmInner__EVAL_30;
  wire [2:0] dmInner__EVAL_31;
  wire  dmInner__EVAL_32;
  wire  dmInner__EVAL_33;
  wire  dmInner__EVAL_34;
  wire  dmInner__EVAL_35;
  wire [11:0] dmInner__EVAL_36;
  wire  dmInner__EVAL_37;
  wire  dmInner__EVAL_38;
  wire [2:0] dmInner__EVAL_39;
  wire [1:0] dmInner__EVAL_40;
  wire  dmInner__EVAL_41;
  _EVAL_147 AsyncQueueSink (
    ._EVAL(AsyncQueueSink__EVAL),
    ._EVAL_0(AsyncQueueSink__EVAL_0),
    ._EVAL_1(AsyncQueueSink__EVAL_1),
    ._EVAL_2(AsyncQueueSink__EVAL_2),
    ._EVAL_3(AsyncQueueSink__EVAL_3),
    ._EVAL_4(AsyncQueueSink__EVAL_4),
    ._EVAL_5(AsyncQueueSink__EVAL_5),
    ._EVAL_6(AsyncQueueSink__EVAL_6),
    ._EVAL_7(AsyncQueueSink__EVAL_7),
    ._EVAL_8(AsyncQueueSink__EVAL_8),
    ._EVAL_9(AsyncQueueSink__EVAL_9),
    ._EVAL_10(AsyncQueueSink__EVAL_10)
  );
  _EVAL_140 dmactiveSync (
    ._EVAL(dmactiveSync__EVAL),
    ._EVAL_0(dmactiveSync__EVAL_0),
    ._EVAL_1(dmactiveSync__EVAL_1),
    ._EVAL_2(dmactiveSync__EVAL_2)
  );
  _EVAL_145 dmiXing (
    ._EVAL(dmiXing__EVAL),
    ._EVAL_0(dmiXing__EVAL_0),
    ._EVAL_1(dmiXing__EVAL_1),
    ._EVAL_2(dmiXing__EVAL_2),
    ._EVAL_3(dmiXing__EVAL_3),
    ._EVAL_4(dmiXing__EVAL_4),
    ._EVAL_5(dmiXing__EVAL_5),
    ._EVAL_6(dmiXing__EVAL_6),
    ._EVAL_7(dmiXing__EVAL_7),
    ._EVAL_8(dmiXing__EVAL_8),
    ._EVAL_9(dmiXing__EVAL_9),
    ._EVAL_10(dmiXing__EVAL_10),
    ._EVAL_11(dmiXing__EVAL_11),
    ._EVAL_12(dmiXing__EVAL_12),
    ._EVAL_13(dmiXing__EVAL_13),
    ._EVAL_14(dmiXing__EVAL_14),
    ._EVAL_15(dmiXing__EVAL_15),
    ._EVAL_16(dmiXing__EVAL_16),
    ._EVAL_17(dmiXing__EVAL_17),
    ._EVAL_18(dmiXing__EVAL_18),
    ._EVAL_19(dmiXing__EVAL_19),
    ._EVAL_20(dmiXing__EVAL_20),
    ._EVAL_21(dmiXing__EVAL_21),
    ._EVAL_22(dmiXing__EVAL_22),
    ._EVAL_23(dmiXing__EVAL_23),
    ._EVAL_24(dmiXing__EVAL_24),
    ._EVAL_25(dmiXing__EVAL_25),
    ._EVAL_26(dmiXing__EVAL_26),
    ._EVAL_27(dmiXing__EVAL_27),
    ._EVAL_28(dmiXing__EVAL_28)
  );
  _EVAL_141 dmInner (
    ._EVAL(dmInner__EVAL),
    ._EVAL_0(dmInner__EVAL_0),
    ._EVAL_1(dmInner__EVAL_1),
    ._EVAL_2(dmInner__EVAL_2),
    ._EVAL_3(dmInner__EVAL_3),
    ._EVAL_4(dmInner__EVAL_4),
    ._EVAL_5(dmInner__EVAL_5),
    ._EVAL_6(dmInner__EVAL_6),
    ._EVAL_7(dmInner__EVAL_7),
    ._EVAL_8(dmInner__EVAL_8),
    ._EVAL_9(dmInner__EVAL_9),
    ._EVAL_10(dmInner__EVAL_10),
    ._EVAL_11(dmInner__EVAL_11),
    ._EVAL_12(dmInner__EVAL_12),
    ._EVAL_13(dmInner__EVAL_13),
    ._EVAL_14(dmInner__EVAL_14),
    ._EVAL_15(dmInner__EVAL_15),
    ._EVAL_16(dmInner__EVAL_16),
    ._EVAL_17(dmInner__EVAL_17),
    ._EVAL_18(dmInner__EVAL_18),
    ._EVAL_19(dmInner__EVAL_19),
    ._EVAL_20(dmInner__EVAL_20),
    ._EVAL_21(dmInner__EVAL_21),
    ._EVAL_22(dmInner__EVAL_22),
    ._EVAL_23(dmInner__EVAL_23),
    ._EVAL_24(dmInner__EVAL_24),
    ._EVAL_25(dmInner__EVAL_25),
    ._EVAL_26(dmInner__EVAL_26),
    ._EVAL_27(dmInner__EVAL_27),
    ._EVAL_28(dmInner__EVAL_28),
    ._EVAL_29(dmInner__EVAL_29),
    ._EVAL_30(dmInner__EVAL_30),
    ._EVAL_31(dmInner__EVAL_31),
    ._EVAL_32(dmInner__EVAL_32),
    ._EVAL_33(dmInner__EVAL_33),
    ._EVAL_34(dmInner__EVAL_34),
    ._EVAL_35(dmInner__EVAL_35),
    ._EVAL_36(dmInner__EVAL_36),
    ._EVAL_37(dmInner__EVAL_37),
    ._EVAL_38(dmInner__EVAL_38),
    ._EVAL_39(dmInner__EVAL_39),
    ._EVAL_40(dmInner__EVAL_40),
    ._EVAL_41(dmInner__EVAL_41)
  );
  assign dmInner__EVAL_26 = _EVAL_13;
  assign dmInner__EVAL_18 = dmactiveSync__EVAL_1;
  assign dmiXing__EVAL_3 = _EVAL_33;
  assign _EVAL_30 = dmInner__EVAL_1;
  assign dmInner__EVAL_15 = dmiXing__EVAL_12;
  assign dmiXing__EVAL_19 = _EVAL_27;
  assign dmiXing__EVAL_13 = dmInner__EVAL_6;
  assign dmInner__EVAL_2 = dmiXing__EVAL_10;
  assign _EVAL_12 = dmInner__EVAL_35;
  assign dmiXing__EVAL_15 = dmInner__EVAL_27;
  assign _EVAL_6 = dmInner__EVAL_8;
  assign dmInner__EVAL_41 = dmiXing__EVAL_16;
  assign dmInner__EVAL_14 = _EVAL_35;
  assign _EVAL_16 = dmiXing__EVAL_7;
  assign dmactiveSync__EVAL = _EVAL_33;
  assign dmInner__EVAL_19 = AsyncQueueSink__EVAL_8;
  assign dmInner__EVAL_20 = _EVAL_20;
  assign dmInner__EVAL_3 = AsyncQueueSink__EVAL_9;
  assign dmInner__EVAL_32 = _EVAL_23;
  assign dmInner__EVAL_38 = _EVAL_33;
  assign dmInner__EVAL_11 = dmiXing__EVAL_4;
  assign dmInner__EVAL_7 = _EVAL_11;
  assign _EVAL_7 = dmiXing__EVAL_20;
  assign AsyncQueueSink__EVAL_1 = _EVAL_28;
  assign dmInner__EVAL_0 = dmiXing__EVAL_25;
  assign _EVAL_21 = dmiXing__EVAL_27;
  assign dmInner__EVAL_36 = _EVAL_4;
  assign dmInner__EVAL = _EVAL_2;
  assign dmInner__EVAL_33 = dmiXing__EVAL_1;
  assign dmInner__EVAL_30 = dmiXing__EVAL_23;
  assign dmiXing__EVAL_22 = _EVAL_2;
  assign _EVAL = dmiXing__EVAL_9;
  assign dmInner__EVAL_39 = _EVAL_10;
  assign dmiXing__EVAL_14 = dmInner__EVAL_37;
  assign dmiXing__EVAL_21 = _EVAL_19;
  assign dmiXing__EVAL_6 = _EVAL_15;
  assign dmiXing__EVAL_5 = dmInner__EVAL_31;
  assign dmInner__EVAL_28 = _EVAL_17;
  assign dmiXing__EVAL_26 = _EVAL_22;
  assign dmInner__EVAL_22 = AsyncQueueSink__EVAL;
  assign dmInner__EVAL_5 = _EVAL_25;
  assign _EVAL_26 = dmiXing__EVAL_0;
  assign dmiXing__EVAL_24 = dmInner__EVAL_10;
  assign dmInner__EVAL_13 = _EVAL_32;
  assign _EVAL_8 = dmInner__EVAL_24;
  assign _EVAL_9 = dmInner__EVAL_9;
  assign dmInner__EVAL_29 = dmiXing__EVAL_28;
  assign AsyncQueueSink__EVAL_3 = _EVAL_0;
  assign AsyncQueueSink__EVAL_7 = _EVAL_3;
  assign dmactiveSync__EVAL_2 = _EVAL_14;
  assign dmInner__EVAL_12 = AsyncQueueSink__EVAL_0;
  assign _EVAL_34 = AsyncQueueSink__EVAL_10;
  assign _EVAL_36 = dmInner__EVAL_4;
  assign AsyncQueueSink__EVAL_6 = _EVAL_2;
  assign AsyncQueueSink__EVAL_4 = _EVAL_33;
  assign dmInner__EVAL_25 = AsyncQueueSink__EVAL_5;
  assign dmiXing__EVAL_8 = _EVAL_18;
  assign dmInner__EVAL_34 = _EVAL_31;
  assign _EVAL_24 = dmiXing__EVAL_11;
  assign _EVAL_5 = dmInner__EVAL_16;
  assign dmInner__EVAL_21 = dmiXing__EVAL_17;
  assign AsyncQueueSink__EVAL_2 = _EVAL_29;
  assign dmactiveSync__EVAL_0 = _EVAL_2;
  assign dmInner__EVAL_40 = dmiXing__EVAL;
  assign dmiXing__EVAL_18 = dmInner__EVAL_23;
  assign dmiXing__EVAL_2 = _EVAL_1;
endmodule
