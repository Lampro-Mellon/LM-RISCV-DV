//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_34_assert(
  input         _EVAL,
  input  [3:0]  _EVAL_0,
  input  [3:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [3:0]  _EVAL_10,
  input         _EVAL_11,
  input  [1:0]  _EVAL_12,
  input  [31:0] _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17
);
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire [32:0] _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire [7:0] _EVAL_34;
  wire [3:0] _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  reg  _EVAL_42;
  reg [31:0] _RAND_0;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire [31:0] _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  reg [5:0] _EVAL_59;
  reg [31:0] _RAND_1;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire [32:0] _EVAL_63;
  reg  _EVAL_64;
  reg [31:0] _RAND_2;
  reg [1:0] _EVAL_65;
  reg [31:0] _RAND_3;
  wire [32:0] _EVAL_66;
  wire  _EVAL_67;
  wire [32:0] _EVAL_68;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire [7:0] _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  reg  _EVAL_86;
  reg [31:0] _RAND_4;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_91;
  wire [32:0] _EVAL_92;
  wire [1:0] _EVAL_93;
  wire [31:0] _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire [3:0] _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire [5:0] _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  reg [31:0] _EVAL_141;
  reg [31:0] _RAND_5;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire [32:0] _EVAL_149;
  wire  _EVAL_150;
  wire [31:0] _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire [3:0] _EVAL_155;
  wire [32:0] _EVAL_157;
  wire  _EVAL_158;
  wire [32:0] _EVAL_159;
  wire [5:0] _EVAL_160;
  wire [32:0] _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire [6:0] _EVAL_165;
  wire [32:0] _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire [31:0] _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  reg [3:0] _EVAL_177;
  reg [31:0] _RAND_6;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire [5:0] _EVAL_180;
  wire [5:0] _EVAL_181;
  reg [2:0] _EVAL_182;
  reg [31:0] _RAND_7;
  wire  _EVAL_183;
  wire [7:0] _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire [6:0] _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire [1:0] _EVAL_201;
  wire [32:0] _EVAL_202;
  wire [32:0] _EVAL_203;
  wire [1:0] _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire [5:0] _EVAL_207;
  wire  _EVAL_208;
  wire [31:0] _EVAL_209;
  wire [32:0] _EVAL_210;
  wire [22:0] _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  reg [2:0] _EVAL_215;
  reg [31:0] _RAND_8;
  wire [32:0] _EVAL_216;
  wire [6:0] _EVAL_217;
  wire  _EVAL_218;
  reg [5:0] _EVAL_219;
  reg [31:0] _RAND_9;
  wire [32:0] _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire [32:0] _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  reg [5:0] _EVAL_234;
  reg [31:0] _RAND_10;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire [32:0] _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire [6:0] _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  reg [5:0] _EVAL_256;
  reg [31:0] _RAND_11;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire [32:0] _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire [31:0] _EVAL_269;
  wire  _EVAL_270;
  wire [1:0] _EVAL_271;
  wire [1:0] _EVAL_272;
  wire [31:0] _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  reg [31:0] _EVAL_280;
  reg [31:0] _RAND_12;
  wire  _EVAL_281;
  wire [22:0] _EVAL_282;
  wire  _EVAL_283;
  reg  _EVAL_284;
  reg [31:0] _RAND_13;
  wire [31:0] _EVAL_285;
  reg [3:0] _EVAL_286;
  reg [31:0] _RAND_14;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_291;
  wire  _EVAL_292;
  reg [2:0] _EVAL_293;
  reg [31:0] _RAND_15;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire [32:0] _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_305;
  wire [5:0] _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire [3:0] _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire [7:0] _EVAL_316;
  wire  _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_212 = _EVAL_45 | _EVAL_3;
  assign _EVAL_135 = _EVAL_5 & _EVAL_301;
  assign _EVAL_82 = ~_EVAL_79;
  assign _EVAL_311 = _EVAL_119 & _EVAL_218;
  assign _EVAL_228 = _EVAL_5 & _EVAL_136;
  assign _EVAL_93 = _EVAL_204 | 2'h1;
  assign _EVAL_314 = _EVAL_2 == 3'h5;
  assign _EVAL_83 = _EVAL_124 | _EVAL_3;
  assign _EVAL_287 = _EVAL_18 | _EVAL_3;
  assign _EVAL_180 = _EVAL_217[5:0];
  assign _EVAL_245 = _EVAL_283 | _EVAL_3;
  assign _EVAL_118 = _EVAL_243 | _EVAL_107;
  assign _EVAL_217 = _EVAL_59 - 6'h1;
  assign _EVAL_220 = _EVAL_66;
  assign _EVAL_25 = _EVAL_303 | _EVAL_3;
  assign _EVAL_152 = _EVAL_272[0];
  assign _EVAL_144 = _EVAL_27 & _EVAL_242;
  assign _EVAL_41 = ~_EVAL_123;
  assign _EVAL_159 = $signed(_EVAL_300) & -33'sh1000000;
  assign _EVAL_230 = ~_EVAL_294;
  assign _EVAL_222 = _EVAL_259 | _EVAL_144;
  assign _EVAL_125 = _EVAL_9 == 3'h0;
  assign _EVAL_131 = ~_EVAL_3;
  assign _EVAL_92 = _EVAL_159;
  assign _EVAL_55 = _EVAL_175 & _EVAL_99;
  assign _EVAL_119 = _EVAL_13[1];
  assign _EVAL_90 = _EVAL_313 & _EVAL_254;
  assign _EVAL_39 = _EVAL_221 & _EVAL_139;
  assign _EVAL_242 = $signed(_EVAL_166) == 33'sh0;
  assign _EVAL_179 = _EVAL_93[0];
  assign _EVAL_68 = {1'b0,$signed(_EVAL_46)};
  assign _EVAL_127 = _EVAL_34[7:2];
  assign _EVAL_270 = _EVAL_105 == 4'h0;
  assign _EVAL_254 = $signed(_EVAL_224) == 33'sh0;
  assign _EVAL_160 = _EVAL_81[7:2];
  assign _EVAL_23 = ~_EVAL_212;
  assign _EVAL_95 = _EVAL_168 | _EVAL_197;
  assign _EVAL_36 = _EVAL_12 <= 2'h2;
  assign _EVAL_153 = _EVAL_42 >> _EVAL_14;
  assign _EVAL_195 = _EVAL_125 | _EVAL_3;
  assign _EVAL_251 = _EVAL_201[0];
  assign _EVAL_145 = ~_EVAL_112;
  assign _EVAL_238 = ~_EVAL_14;
  assign _EVAL_52 = _EVAL_119 & _EVAL_239;
  assign _EVAL_239 = _EVAL_13[0];
  assign _EVAL_264 = _EVAL_2[0];
  assign _EVAL_37 = _EVAL_10 >= 4'h2;
  assign _EVAL_30 = $signed(_EVAL_92) == 33'sh0;
  assign _EVAL_75 = _EVAL_5 & _EVAL_274;
  assign _EVAL_184 = _EVAL_282[7:0];
  assign _EVAL_73 = ~_EVAL_312;
  assign _EVAL_278 = _EVAL_235 | _EVAL_84;
  assign _EVAL_175 = _EVAL_42 | _EVAL_251;
  assign _EVAL_218 = ~_EVAL_239;
  assign _EVAL_173 = $signed(_EVAL_21) == 33'sh0;
  assign _EVAL_295 = _EVAL_100 | _EVAL_90;
  assign _EVAL_189 = _EVAL_219 - 6'h1;
  assign _EVAL_300 = {1'b0,$signed(_EVAL_285)};
  assign _EVAL_302 = ~_EVAL_158;
  assign _EVAL_285 = _EVAL_13 ^ 32'h2000000;
  assign _EVAL_32 = _EVAL_292 | _EVAL_3;
  assign _EVAL_306 = _EVAL_165[5:0];
  assign _EVAL_190 = ~_EVAL_281;
  assign _EVAL_233 = _EVAL_12 == 2'h0;
  assign _EVAL_44 = ~_EVAL_208;
  assign _EVAL_166 = _EVAL_203;
  assign _EVAL_123 = _EVAL_238 | _EVAL_3;
  assign _EVAL_139 = _EVAL_234 == 6'h0;
  assign _EVAL_281 = _EVAL_270 | _EVAL_3;
  assign _EVAL_47 = _EVAL_129 & _EVAL_176;
  assign _EVAL_27 = _EVAL_0 <= 4'h6;
  assign _EVAL_130 = ~_EVAL_310;
  assign _EVAL_176 = _EVAL_59 == 6'h0;
  assign _EVAL_161 = $signed(_EVAL_63) & -33'sh1000;
  assign _EVAL_26 = ~_EVAL_88;
  assign _EVAL_246 = _EVAL_256 == 6'h0;
  assign _EVAL_203 = $signed(_EVAL_266) & -33'sh2000;
  assign _EVAL_274 = _EVAL_4 == 3'h0;
  assign _EVAL_299 = ~_EVAL_255;
  assign _EVAL_148 = _EVAL_296 | _EVAL_197;
  assign _EVAL_307 = _EVAL_0 <= 4'h2;
  assign _EVAL_196 = ~_EVAL_289;
  assign _EVAL_40 = _EVAL_2 == 3'h1;
  assign _EVAL_165 = _EVAL_256 - 6'h1;
  assign _EVAL_34 = ~_EVAL_184;
  assign _EVAL_167 = _EVAL_4 == _EVAL_182;
  assign _EVAL_147 = ~_EVAL_121;
  assign _EVAL_56 = _EVAL_179 & _EVAL_52;
  assign _EVAL_122 = _EVAL_235 | _EVAL_140;
  assign _EVAL_275 = _EVAL_221 & _EVAL_267;
  assign _EVAL_114 = ~_EVAL_317;
  assign _EVAL_205 = _EVAL_11 & _EVAL_87;
  assign _EVAL_181 = _EVAL_189[5:0];
  assign _EVAL_185 = _EVAL_57 | _EVAL_3;
  assign _EVAL_45 = _EVAL_2 == _EVAL_215;
  assign _EVAL_193 = _EVAL_305 | _EVAL_3;
  assign _EVAL_279 = _EVAL_12 == _EVAL_65;
  assign _EVAL_291 = _EVAL_11 & _EVAL_24;
  assign _EVAL_288 = _EVAL_232 | _EVAL_174;
  assign _EVAL_128 = _EVAL_5 & _EVAL_74;
  assign _EVAL_158 = _EVAL_298 | _EVAL_3;
  assign _EVAL_292 = _EVAL_9 <= 3'h1;
  assign _EVAL_46 = _EVAL_13 ^ 32'h80000000;
  assign _EVAL_163 = _EVAL_17 == _EVAL_64;
  assign _EVAL_310 = _EVAL_102 | _EVAL_3;
  assign _EVAL_97 = ~_EVAL_137;
  assign _EVAL_255 = _EVAL_188 | _EVAL_3;
  assign _EVAL_200 = _EVAL_315 | _EVAL_56;
  assign _EVAL_109 = _EVAL_36 | _EVAL_3;
  assign _EVAL_277 = _EVAL_0 >= 4'h2;
  assign _EVAL_211 = 23'hff << _EVAL_0;
  assign _EVAL_84 = _EVAL_179 & _EVAL_241;
  assign _EVAL_149 = {1'b0,$signed(_EVAL_13)};
  assign _EVAL_315 = _EVAL_277 | _EVAL_258;
  assign _EVAL_223 = ~_EVAL_25;
  assign _EVAL_241 = _EVAL_240 & _EVAL_218;
  assign _EVAL_305 = _EVAL_9 <= 3'h2;
  assign _EVAL_260 = _EVAL_57 | _EVAL_15;
  assign _EVAL_201 = _EVAL_39 ? _EVAL_271 : 2'h0;
  assign _EVAL_258 = _EVAL_133 & _EVAL_119;
  assign _EVAL_243 = ~_EVAL_42;
  assign _EVAL_67 = ~_EVAL_225;
  assign _EVAL_318 = _EVAL_280 < plusarg_reader_out;
  assign _EVAL_266 = {1'b0,$signed(_EVAL_94)};
  assign _EVAL_87 = _EVAL_2 == 3'h2;
  assign _EVAL_169 = ~_EVAL_195;
  assign _EVAL_20 = _EVAL_213 | _EVAL_265;
  assign _EVAL_240 = ~_EVAL_119;
  assign _EVAL_194 = ~_EVAL_245;
  assign _EVAL_31 = _EVAL_4 == 3'h6;
  assign _EVAL_112 = _EVAL_2 == 3'h6;
  assign _EVAL_308 = _EVAL_20 | _EVAL_3;
  assign _EVAL_262 = ~_EVAL_319;
  assign _EVAL_294 = _EVAL_4[2];
  assign _EVAL_183 = ~_EVAL_198;
  assign _EVAL_94 = _EVAL_13 ^ 32'h40000000;
  assign _EVAL_85 = ~_EVAL_70;
  assign _EVAL_283 = _EVAL == _EVAL_284;
  assign _EVAL_235 = _EVAL_277 | _EVAL_120;
  assign _EVAL_88 = _EVAL_37 | _EVAL_3;
  assign _EVAL_28 = _EVAL_2 <= 3'h6;
  assign _EVAL_186 = ~_EVAL_113;
  assign _EVAL_312 = _EVAL_279 | _EVAL_3;
  assign _EVAL_96 = _EVAL_9 == _EVAL_293;
  assign _EVAL_77 = _EVAL_4 == 3'h1;
  assign _EVAL_150 = _EVAL_5 & _EVAL_89;
  assign _EVAL_115 = _EVAL_11 & _EVAL_112;
  assign _EVAL_168 = _EVAL_173 | _EVAL_30;
  assign _EVAL_72 = _EVAL_4 == 3'h7;
  assign _EVAL_105 = _EVAL_1 & _EVAL_155;
  assign _EVAL_206 = _EVAL_118 | _EVAL_318;
  assign _EVAL_225 = _EVAL_49 | _EVAL_3;
  assign _EVAL_296 = _EVAL_254 | _EVAL_30;
  assign _EVAL_282 = 23'hff << _EVAL_10;
  assign _EVAL_100 = _EVAL_307 & _EVAL_95;
  assign _EVAL_29 = ~_EVAL_32;
  assign _EVAL_209 = _EVAL_210[31:0];
  assign _EVAL_138 = ~_EVAL_261;
  assign _EVAL_250 = _EVAL_234 - 6'h1;
  assign _EVAL_157 = {1'b0,$signed(_EVAL_269)};
  assign _EVAL_202 = $signed(_EVAL_149) & -33'sh5000;
  assign _EVAL_143 = _EVAL_233 | _EVAL_3;
  assign _EVAL_103 = _EVAL_12 != 2'h2;
  assign _EVAL_33 = _EVAL_117 | _EVAL_3;
  assign _EVAL_208 = _EVAL_38 | _EVAL_3;
  assign _EVAL_74 = _EVAL_4 == 3'h3;
  assign _EVAL_61 = _EVAL_0[0];
  assign _EVAL_140 = _EVAL_179 & _EVAL_268;
  assign _EVAL_133 = _EVAL_93[1];
  assign _EVAL_191 = ~_EVAL_227;
  assign _EVAL_265 = _EVAL_307 & _EVAL_71;
  assign _EVAL_50 = _EVAL_162 | _EVAL_3;
  assign _EVAL_276 = ~_EVAL_287;
  assign _EVAL_192 = _EVAL_5 & _EVAL_31;
  assign _EVAL_271 = 2'h1 << _EVAL_14;
  assign _EVAL_154 = ~_EVAL_308;
  assign _EVAL_174 = ~_EVAL_251;
  assign _EVAL_187 = _EVAL_273 == 32'h0;
  assign _EVAL_106 = ~_EVAL_83;
  assign _EVAL_309 = {_EVAL_200,_EVAL_58,_EVAL_122,_EVAL_278};
  assign _EVAL_207 = _EVAL_250[5:0];
  assign _EVAL_136 = ~_EVAL_267;
  assign _EVAL_172 = {{24'd0}, _EVAL_81};
  assign _EVAL_273 = _EVAL_13 & _EVAL_172;
  assign _EVAL_146 = _EVAL_129 & _EVAL_246;
  assign _EVAL_224 = _EVAL_161;
  assign _EVAL_63 = {1'b0,$signed(_EVAL_151)};
  assign _EVAL_204 = 2'h1 << _EVAL_61;
  assign _EVAL_252 = ~_EVAL_91;
  assign _EVAL_62 = ~_EVAL_15;
  assign _EVAL_272 = _EVAL_134 ? 2'h1 : 2'h0;
  assign _EVAL_155 = ~_EVAL_309;
  assign _EVAL_289 = _EVAL_111 | _EVAL_3;
  assign _EVAL_214 = ~_EVAL_109;
  assign _EVAL_101 = _EVAL_222 | _EVAL_90;
  assign _EVAL_151 = _EVAL_13 ^ 32'h3000;
  assign _EVAL_231 = ~_EVAL_185;
  assign _EVAL_213 = _EVAL_144 | _EVAL_90;
  assign _EVAL_229 = ~_EVAL_176;
  assign _EVAL_54 = _EVAL_260 | _EVAL_3;
  assign _EVAL_53 = ~_EVAL_193;
  assign _EVAL_188 = _EVAL_9 <= 3'h3;
  assign _EVAL_301 = _EVAL_4 == 3'h5;
  assign _EVAL_244 = _EVAL_171 | _EVAL_3;
  assign _EVAL_170 = _EVAL_2 == 3'h0;
  assign _EVAL_108 = _EVAL_11 & _EVAL_40;
  assign _EVAL_236 = ~_EVAL_54;
  assign _EVAL_117 = _EVAL_13 == _EVAL_141;
  assign _EVAL_316 = _EVAL_211[7:0];
  assign _EVAL_303 = _EVAL_9 != 3'h0;
  assign _EVAL_197 = $signed(_EVAL_237) == 33'sh0;
  assign _EVAL_111 = _EVAL_14 == _EVAL_86;
  assign _EVAL_129 = _EVAL_7 & _EVAL_11;
  assign _EVAL_22 = ~_EVAL_244;
  assign _EVAL_19 = _EVAL_5 & _EVAL_132;
  assign _EVAL_313 = _EVAL_0 <= 4'h8;
  assign _EVAL_171 = _EVAL_307 & _EVAL_164;
  assign _EVAL_48 = ~_EVAL_143;
  assign _EVAL_247 = ~_EVAL_33;
  assign _EVAL_58 = _EVAL_315 | _EVAL_297;
  assign _EVAL_78 = _EVAL_5 & _EVAL_72;
  assign _EVAL_134 = _EVAL_146 & _EVAL_145;
  assign _EVAL_248 = ~_EVAL_153;
  assign _EVAL_232 = _EVAL_251 != _EVAL_152;
  assign _EVAL_269 = _EVAL_13 ^ 32'h20000000;
  assign _EVAL_104 = _EVAL_95 | _EVAL_71;
  assign _EVAL_267 = _EVAL_219 == 6'h0;
  assign _EVAL_21 = _EVAL_216;
  assign _EVAL_51 = _EVAL_11 & _EVAL_229;
  assign _EVAL_137 = _EVAL_101 | _EVAL_3;
  assign _EVAL_80 = _EVAL_11 & _EVAL_314;
  assign _EVAL_120 = _EVAL_133 & _EVAL_240;
  assign _EVAL_91 = _EVAL_62 | _EVAL_3;
  assign _EVAL_18 = _EVAL_1 == _EVAL_309;
  assign _EVAL_268 = _EVAL_240 & _EVAL_239;
  assign _EVAL_317 = _EVAL_288 | _EVAL_3;
  assign _EVAL_261 = _EVAL_163 | _EVAL_3;
  assign _EVAL_227 = _EVAL_167 | _EVAL_3;
  assign _EVAL_226 = _EVAL_11 & _EVAL_170;
  assign _EVAL_132 = _EVAL_4 == 3'h2;
  assign _EVAL_57 = ~_EVAL;
  assign _EVAL_49 = _EVAL_251 | _EVAL_42;
  assign _EVAL_216 = $signed(_EVAL_68) & -33'shc000;
  assign _EVAL_253 = _EVAL_295 | _EVAL_3;
  assign _EVAL_99 = ~_EVAL_152;
  assign _EVAL_102 = _EVAL_9 <= 3'h4;
  assign _EVAL_38 = ~_EVAL_6;
  assign _EVAL_298 = _EVAL_0 == _EVAL_177;
  assign _EVAL_79 = _EVAL_206 | _EVAL_3;
  assign _EVAL_81 = ~_EVAL_316;
  assign _EVAL_35 = ~_EVAL_1;
  assign _EVAL_178 = ~_EVAL_253;
  assign _EVAL_89 = _EVAL_4 == 3'h4;
  assign _EVAL_237 = _EVAL_202;
  assign _EVAL_164 = _EVAL_148 | _EVAL_71;
  assign _EVAL_259 = _EVAL_307 & _EVAL_104;
  assign _EVAL_221 = _EVAL_8 & _EVAL_5;
  assign _EVAL_198 = _EVAL_96 | _EVAL_3;
  assign _EVAL_121 = _EVAL_248 | _EVAL_3;
  assign _EVAL_199 = _EVAL_5 & _EVAL_77;
  assign _EVAL_263 = _EVAL_187 | _EVAL_3;
  assign _EVAL_24 = _EVAL_2 == 3'h4;
  assign _EVAL_124 = _EVAL_35 == 4'h0;
  assign _EVAL_66 = $signed(_EVAL_157) & -33'sh2000;
  assign _EVAL_71 = $signed(_EVAL_220) == 33'sh0;
  assign _EVAL_43 = ~_EVAL_263;
  assign _EVAL_162 = _EVAL_10 == _EVAL_286;
  assign _EVAL_107 = plusarg_reader_out == 32'h0;
  assign _EVAL_70 = _EVAL_277 | _EVAL_3;
  assign _EVAL_297 = _EVAL_179 & _EVAL_311;
  assign _EVAL_110 = ~_EVAL_50;
  assign _EVAL_319 = _EVAL_28 | _EVAL_3;
  assign _EVAL_210 = _EVAL_280 + 32'h1;
  assign _EVAL_60 = _EVAL_221 | _EVAL_129;
  assign _EVAL_113 = _EVAL_103 | _EVAL_3;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_42 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_59 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_64 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_65 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_86 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_141 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_177 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_182 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_215 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_219 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_234 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_256 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_280 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_284 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_286 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_293 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_16) begin
    if (_EVAL_3) begin
      _EVAL_42 <= 1'h0;
    end else begin
      _EVAL_42 <= _EVAL_55;
    end
    if (_EVAL_3) begin
      _EVAL_59 <= 6'h0;
    end else if (_EVAL_129) begin
      if (_EVAL_176) begin
        if (_EVAL_264) begin
          _EVAL_59 <= _EVAL_127;
        end else begin
          _EVAL_59 <= 6'h0;
        end
      end else begin
        _EVAL_59 <= _EVAL_180;
      end
    end
    if (_EVAL_47) begin
      _EVAL_64 <= _EVAL_17;
    end
    if (_EVAL_47) begin
      _EVAL_65 <= _EVAL_12;
    end
    if (_EVAL_275) begin
      _EVAL_86 <= _EVAL_14;
    end
    if (_EVAL_275) begin
      _EVAL_141 <= _EVAL_13;
    end
    if (_EVAL_275) begin
      _EVAL_177 <= _EVAL_0;
    end
    if (_EVAL_275) begin
      _EVAL_182 <= _EVAL_4;
    end
    if (_EVAL_47) begin
      _EVAL_215 <= _EVAL_2;
    end
    if (_EVAL_3) begin
      _EVAL_219 <= 6'h0;
    end else if (_EVAL_221) begin
      if (_EVAL_267) begin
        if (_EVAL_230) begin
          _EVAL_219 <= _EVAL_160;
        end else begin
          _EVAL_219 <= 6'h0;
        end
      end else begin
        _EVAL_219 <= _EVAL_181;
      end
    end
    if (_EVAL_3) begin
      _EVAL_234 <= 6'h0;
    end else if (_EVAL_221) begin
      if (_EVAL_139) begin
        if (_EVAL_230) begin
          _EVAL_234 <= _EVAL_160;
        end else begin
          _EVAL_234 <= 6'h0;
        end
      end else begin
        _EVAL_234 <= _EVAL_207;
      end
    end
    if (_EVAL_3) begin
      _EVAL_256 <= 6'h0;
    end else if (_EVAL_129) begin
      if (_EVAL_246) begin
        if (_EVAL_264) begin
          _EVAL_256 <= _EVAL_127;
        end else begin
          _EVAL_256 <= 6'h0;
        end
      end else begin
        _EVAL_256 <= _EVAL_306;
      end
    end
    if (_EVAL_3) begin
      _EVAL_280 <= 32'h0;
    end else if (_EVAL_60) begin
      _EVAL_280 <= 32'h0;
    end else begin
      _EVAL_280 <= _EVAL_209;
    end
    if (_EVAL_47) begin
      _EVAL_284 <= _EVAL;
    end
    if (_EVAL_47) begin
      _EVAL_286 <= _EVAL_10;
    end
    if (_EVAL_275) begin
      _EVAL_293 <= _EVAL_9;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34632ca1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90e22a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c177d18d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc314e50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(369077f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(465fce12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7adf06e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4bae639)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_299) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca30466)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d8848d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bba0c2e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8be912f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa0abf92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57d2fec9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_134 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28a9879d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ce7531c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d89b8453)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1daf685a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(208dcbf8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3912be28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7f102fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d937c08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cf0dc75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e790f01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f3525b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6cbba41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9240abbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab5e459e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fe4c81a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26fecdf8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba2e4f70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23feba50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44d3f7da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7421a34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(175dafbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79d18ce6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40871b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddcb5f7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_73) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(741e66e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0f289ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59a1dfe4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2092f6b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae1ad682)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b06895e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(313d003e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b964e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c319d632)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c74db1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44754457)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fa6121d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48fa28e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ebdeb10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(978ab502)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a0c5e36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d893cab3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86ce4d2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46af7571)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b467402)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6861f0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf36ec7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14a18051)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(574c5cf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f652f07f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db772d11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2286dbcc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efe40a73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58cfa186)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb4e2c12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc2ac95a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ee80d56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df56b9a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60dac0f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37948ada)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ff33e01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(383e8c8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_115 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ba8c988)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3475bd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(440b477f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bd9318a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4cc4c9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_73) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1557a2c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47acfcf1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_299) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91869bd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7b8d717)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
