//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_73_assert(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [13:0] _EVAL_2,
  input         _EVAL_3,
  input  [1:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [3:0]  _EVAL_13,
  input  [3:0]  _EVAL_14,
  input  [2:0]  _EVAL_15,
  input  [3:0]  _EVAL_16,
  input  [2:0]  _EVAL_17,
  input         _EVAL_18
);
  wire  _EVAL_19;
  wire  _EVAL_20;
  reg [2:0] _EVAL_21;
  reg [31:0] _RAND_0;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire [5:0] _EVAL_24;
  wire  _EVAL_25;
  wire [6:0] _EVAL_26;
  wire  _EVAL_27;
  reg [5:0] _EVAL_28;
  reg [31:0] _RAND_1;
  wire  _EVAL_29;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire [7:0] _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire [4:0] _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire [4:0] _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire [4:0] _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  reg [5:0] _EVAL_54;
  reg [31:0] _RAND_2;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire [1:0] _EVAL_58;
  reg [1:0] _EVAL_59;
  reg [31:0] _RAND_3;
  wire  _EVAL_60;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire [32:0] _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire [14:0] _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire [4:0] _EVAL_87;
  wire  _EVAL_88;
  wire [3:0] _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  reg [5:0] _EVAL_94;
  reg [31:0] _RAND_4;
  wire  _EVAL_95;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire [6:0] _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  reg  _EVAL_116;
  reg [31:0] _RAND_5;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire [7:0] _EVAL_123;
  wire  _EVAL_124;
  wire [5:0] _EVAL_125;
  reg [13:0] _EVAL_126;
  reg [31:0] _RAND_6;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire [7:0] _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire [5:0] _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire [7:0] _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire [5:0] _EVAL_153;
  wire  _EVAL_154;
  wire [4:0] _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  reg  _EVAL_163;
  reg [31:0] _RAND_7;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire [5:0] _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [3:0] _EVAL_174;
  wire  _EVAL_175;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  reg [31:0] _EVAL_182;
  reg [31:0] _RAND_8;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire [3:0] _EVAL_189;
  reg [2:0] _EVAL_190;
  reg [31:0] _RAND_9;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire [14:0] _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire [7:0] _EVAL_205;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire [22:0] _EVAL_212;
  wire  _EVAL_213;
  reg [5:0] _EVAL_214;
  reg [31:0] _RAND_10;
  wire [7:0] _EVAL_215;
  reg [3:0] _EVAL_216;
  reg [31:0] _RAND_11;
  wire  _EVAL_217;
  wire [7:0] _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  reg [2:0] _EVAL_223;
  reg [31:0] _RAND_12;
  wire  _EVAL_224;
  wire [3:0] _EVAL_225;
  wire [13:0] _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  reg [2:0] _EVAL_233;
  reg [31:0] _RAND_13;
  wire [4:0] _EVAL_234;
  wire [31:0] _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire [5:0] _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire [6:0] _EVAL_244;
  wire [1:0] _EVAL_245;
  wire [7:0] _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire [1:0] _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  reg [2:0] _EVAL_258;
  reg [31:0] _RAND_14;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire [14:0] _EVAL_267;
  wire [13:0] _EVAL_268;
  wire [4:0] _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire [13:0] _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire [6:0] _EVAL_279;
  reg [3:0] _EVAL_280;
  reg [31:0] _RAND_15;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire [1:0] _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire [4:0] _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire [22:0] _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  reg [4:0] _EVAL_299;
  reg [31:0] _RAND_16;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_132 = _EVAL_176 | _EVAL_6;
  assign _EVAL_101 = _EVAL_4 == 2'h0;
  assign _EVAL_285 = _EVAL_245 | 2'h1;
  assign _EVAL_215 = _EVAL_212[7:0];
  assign _EVAL_179 = _EVAL_8 & _EVAL_20;
  assign _EVAL_43 = _EVAL_265 | _EVAL_6;
  assign _EVAL_102 = _EVAL_2 == _EVAL_126;
  assign _EVAL_164 = _EVAL_52 | _EVAL_6;
  assign _EVAL_270 = _EVAL_41 != _EVAL_47;
  assign _EVAL_91 = ~_EVAL_84;
  assign _EVAL_181 = _EVAL_238 & _EVAL_68;
  assign _EVAL_31 = _EVAL_5 <= 3'h3;
  assign _EVAL_36 = _EVAL_8 & _EVAL_75;
  assign _EVAL_154 = _EVAL_285[1];
  assign _EVAL_247 = ~_EVAL_172;
  assign _EVAL_240 = ~_EVAL_56;
  assign _EVAL_98 = ~_EVAL_185;
  assign _EVAL_275 = ~_EVAL_108;
  assign _EVAL_145 = _EVAL_16 <= 4'h2;
  assign _EVAL_142 = _EVAL_7 == 3'h1;
  assign _EVAL_77 = ~_EVAL_184;
  assign _EVAL_24 = _EVAL_148[7:2];
  assign _EVAL_235 = _EVAL_64[31:0];
  assign _EVAL_128 = ~_EVAL_19;
  assign _EVAL_241 = _EVAL_109[5:0];
  assign _EVAL_55 = _EVAL_15 == 3'h5;
  assign _EVAL_39 = ~_EVAL_147;
  assign _EVAL_184 = _EVAL_166 | _EVAL_6;
  assign _EVAL_290 = _EVAL_195 | _EVAL_6;
  assign _EVAL_23 = _EVAL_44 | _EVAL_162;
  assign _EVAL_114 = _EVAL_250 == 2'h1;
  assign _EVAL_34 = _EVAL_101 | _EVAL_6;
  assign _EVAL_67 = ~_EVAL_164;
  assign _EVAL_62 = _EVAL_45 | _EVAL_6;
  assign _EVAL_125 = _EVAL_279[5:0];
  assign _EVAL_213 = _EVAL_255 | _EVAL_65;
  assign _EVAL_151 = _EVAL_150 | _EVAL_137;
  assign _EVAL_47 = _EVAL_33[4:0];
  assign _EVAL_177 = _EVAL_7 == 3'h5;
  assign _EVAL_266 = ~_EVAL_88;
  assign _EVAL_191 = _EVAL_8 & _EVAL_98;
  assign _EVAL_20 = _EVAL_15 == 3'h1;
  assign _EVAL_272 = _EVAL_2 & _EVAL_226;
  assign _EVAL_111 = _EVAL_286 & _EVAL_232;
  assign _EVAL_74 = _EVAL_8 & _EVAL_55;
  assign _EVAL_66 = _EVAL_159 | _EVAL_6;
  assign _EVAL_107 = _EVAL_5 <= 3'h1;
  assign _EVAL_58 = _EVAL_17[2:1];
  assign _EVAL_232 = _EVAL_247 & _EVAL_69;
  assign _EVAL_65 = _EVAL_286 & _EVAL_161;
  assign _EVAL_93 = _EVAL_178 | _EVAL_238;
  assign _EVAL_110 = _EVAL_16 >= 4'h2;
  assign _EVAL_149 = _EVAL_155[0];
  assign _EVAL_231 = _EVAL_12 & _EVAL_177;
  assign _EVAL_198 = _EVAL_4 != 2'h2;
  assign _EVAL_273 = _EVAL_15 == 3'h7;
  assign _EVAL_242 = ~_EVAL_83;
  assign _EVAL_197 = _EVAL_138 & _EVAL_275;
  assign _EVAL_217 = _EVAL_15 == 3'h0;
  assign _EVAL_99 = _EVAL_58 == 2'h1;
  assign _EVAL_48 = ~_EVAL_170;
  assign _EVAL_264 = _EVAL_7 <= 3'h6;
  assign _EVAL_113 = _EVAL_5 == 3'h0;
  assign _EVAL_238 = _EVAL_1 & _EVAL_12;
  assign _EVAL_57 = _EVAL_102 | _EVAL_6;
  assign _EVAL_56 = _EVAL_107 | _EVAL_6;
  assign _EVAL_69 = ~_EVAL_112;
  assign _EVAL_161 = _EVAL_247 & _EVAL_112;
  assign _EVAL_83 = _EVAL_87[0];
  assign _EVAL_106 = ~_EVAL_144;
  assign _EVAL_73 = {1'b0,$signed(_EVAL_268)};
  assign _EVAL_276 = _EVAL_287 | _EVAL_6;
  assign _EVAL_262 = _EVAL_105 | _EVAL_6;
  assign _EVAL_159 = _EVAL_271 | _EVAL_3;
  assign _EVAL_277 = $signed(_EVAL_199) == 15'sh0;
  assign _EVAL_169 = _EVAL_26[5:0];
  assign _EVAL_260 = ~_EVAL_219;
  assign _EVAL_259 = _EVAL_4 == _EVAL_59;
  assign _EVAL_173 = _EVAL_15 == 3'h2;
  assign _EVAL_220 = _EVAL_7 == 3'h0;
  assign _EVAL_180 = _EVAL_293 | _EVAL_6;
  assign _EVAL_225 = ~_EVAL_14;
  assign _EVAL_158 = ~_EVAL_85;
  assign _EVAL_269 = _EVAL_234 & _EVAL_288;
  assign _EVAL_183 = ~_EVAL_43;
  assign _EVAL_204 = ~_EVAL_221;
  assign _EVAL_75 = _EVAL_15 == 3'h6;
  assign _EVAL_118 = ~_EVAL_86;
  assign _EVAL_80 = _EVAL_8 & _EVAL_217;
  assign _EVAL_178 = _EVAL_18 & _EVAL_8;
  assign _EVAL_51 = _EVAL_150 | _EVAL_103;
  assign _EVAL_265 = _EVAL_17 == _EVAL_233;
  assign _EVAL_26 = _EVAL_214 - 6'h1;
  assign _EVAL_144 = _EVAL_299 != 5'h0;
  assign _EVAL_268 = _EVAL_2 ^ 14'h3000;
  assign _EVAL_119 = ~_EVAL_34;
  assign _EVAL_42 = _EVAL_242 | _EVAL_6;
  assign _EVAL_70 = _EVAL_133 | _EVAL_6;
  assign _EVAL_246 = 8'h1 << _EVAL;
  assign _EVAL_38 = _EVAL_5 <= 3'h4;
  assign _EVAL_187 = _EVAL_31 | _EVAL_6;
  assign _EVAL_92 = _EVAL_90 == 4'h0;
  assign _EVAL_288 = ~_EVAL_47;
  assign _EVAL_25 = _EVAL_250 == 2'h0;
  assign _EVAL_227 = _EVAL_71 | _EVAL_22;
  assign _EVAL_278 = ~_EVAL_78;
  assign _EVAL_41 = _EVAL_205[4:0];
  assign _EVAL_257 = ~_EVAL_122;
  assign _EVAL_196 = _EVAL_214 == 6'h0;
  assign _EVAL_193 = _EVAL_172 & _EVAL_69;
  assign _EVAL_103 = _EVAL_286 & _EVAL_193;
  assign _EVAL_19 = _EVAL_237 | _EVAL_6;
  assign _EVAL_76 = _EVAL_12 & _EVAL_142;
  assign _EVAL_104 = _EVAL_154 & _EVAL_172;
  assign _EVAL_292 = _EVAL_54 == 6'h0;
  assign _EVAL_136 = _EVAL_7 == 3'h2;
  assign _EVAL_109 = _EVAL_94 - 6'h1;
  assign _EVAL_281 = ~_EVAL_207;
  assign _EVAL_207 = _EVAL_264 | _EVAL_6;
  assign _EVAL_200 = _EVAL_225 == 4'h0;
  assign _EVAL_279 = _EVAL_28 - 6'h1;
  assign _EVAL_293 = _EVAL_14 == _EVAL_174;
  assign _EVAL_255 = _EVAL_110 | _EVAL_188;
  assign _EVAL_239 = ~_EVAL_6;
  assign _EVAL_298 = _EVAL_23 | _EVAL_6;
  assign _EVAL_84 = _EVAL_38 | _EVAL_6;
  assign _EVAL_88 = _EVAL_198 | _EVAL_6;
  assign _EVAL_123 = ~_EVAL_215;
  assign _EVAL_172 = _EVAL_2[1];
  assign _EVAL_205 = _EVAL_130 ? _EVAL_135 : 8'h0;
  assign _EVAL_146 = _EVAL_228 & _EVAL_277;
  assign _EVAL_252 = ~_EVAL_63;
  assign _EVAL_244 = _EVAL_54 - 6'h1;
  assign _EVAL_138 = _EVAL_238 & _EVAL_292;
  assign _EVAL_33 = _EVAL_197 ? _EVAL_246 : 8'h0;
  assign _EVAL_243 = ~_EVAL_68;
  assign _EVAL_165 = _EVAL_41 != 5'h0;
  assign _EVAL_221 = _EVAL_32 | _EVAL_6;
  assign _EVAL_295 = 23'hff << _EVAL_16;
  assign _EVAL_245 = 2'h1 << _EVAL_251;
  assign _EVAL_237 = _EVAL == _EVAL_21;
  assign _EVAL_105 = _EVAL_272 == 14'h0;
  assign _EVAL_143 = _EVAL_178 & _EVAL_185;
  assign _EVAL_22 = _EVAL_182 < plusarg_reader_out;
  assign _EVAL_32 = _EVAL_5 <= 3'h2;
  assign _EVAL_192 = _EVAL_15 == 3'h3;
  assign _EVAL_194 = ~_EVAL_298;
  assign _EVAL_254 = ~_EVAL_187;
  assign _EVAL_171 = _EVAL_201 | _EVAL_6;
  assign _EVAL_256 = ~_EVAL_261;
  assign _EVAL_287 = _EVAL_145 & _EVAL_277;
  assign _EVAL_188 = _EVAL_154 & _EVAL_247;
  assign _EVAL_224 = ~_EVAL_66;
  assign _EVAL_35 = ~_EVAL_296;
  assign _EVAL_291 = _EVAL_117 | _EVAL_6;
  assign _EVAL_139 = ~_EVAL_180;
  assign _EVAL_166 = ~_EVAL_10;
  assign _EVAL_261 = _EVAL_15[2];
  assign _EVAL_230 = _EVAL_4 <= 2'h2;
  assign _EVAL_286 = _EVAL_285[0];
  assign _EVAL_294 = _EVAL_8 & _EVAL_273;
  assign _EVAL_219 = _EVAL_146 | _EVAL_6;
  assign _EVAL_250 = _EVAL[2:1];
  assign _EVAL_121 = ~_EVAL_291;
  assign _EVAL_162 = _EVAL_17 == 3'h4;
  assign _EVAL_79 = _EVAL_12 & _EVAL_108;
  assign _EVAL_87 = _EVAL_299 >> _EVAL_17;
  assign _EVAL_202 = _EVAL_8 & _EVAL_173;
  assign _EVAL_236 = ~_EVAL_132;
  assign _EVAL_168 = _EVAL_230 | _EVAL_6;
  assign _EVAL_152 = ~_EVAL_276;
  assign _EVAL_108 = _EVAL_7 == 3'h6;
  assign _EVAL_249 = _EVAL_172 & _EVAL_112;
  assign _EVAL_153 = _EVAL_123[7:2];
  assign _EVAL_148 = ~_EVAL_218;
  assign _EVAL_209 = ~_EVAL_127;
  assign _EVAL_85 = _EVAL_92 | _EVAL_6;
  assign _EVAL_141 = _EVAL_244[5:0];
  assign _EVAL_289 = _EVAL_200 | _EVAL_6;
  assign _EVAL_46 = _EVAL_12 & _EVAL_243;
  assign _EVAL_53 = _EVAL_8 & _EVAL_274;
  assign _EVAL_49 = _EVAL_8 & _EVAL_192;
  assign _EVAL_160 = ~_EVAL_81;
  assign _EVAL_130 = _EVAL_178 & _EVAL_196;
  assign _EVAL_124 = ~_EVAL_165;
  assign _EVAL_72 = ~_EVAL_289;
  assign _EVAL_45 = _EVAL_13 == _EVAL_280;
  assign _EVAL_44 = _EVAL_99 | _EVAL_140;
  assign _EVAL_81 = _EVAL_271 | _EVAL_6;
  assign _EVAL_271 = ~_EVAL_9;
  assign _EVAL_50 = _EVAL_0 == _EVAL_116;
  assign _EVAL_228 = _EVAL_16 <= 4'h8;
  assign _EVAL_185 = _EVAL_94 == 6'h0;
  assign _EVAL_157 = ~_EVAL_62;
  assign _EVAL_251 = _EVAL_16[0];
  assign _EVAL_199 = _EVAL_267;
  assign _EVAL_150 = _EVAL_110 | _EVAL_104;
  assign _EVAL_40 = _EVAL_9 == _EVAL_163;
  assign _EVAL_170 = _EVAL_115 | _EVAL_6;
  assign _EVAL_135 = 8'h1 << _EVAL_17;
  assign _EVAL_29 = ~_EVAL_168;
  assign _EVAL_156 = _EVAL_210 | _EVAL_6;
  assign _EVAL_212 = 23'hff << _EVAL_13;
  assign _EVAL_274 = _EVAL_15 == 3'h4;
  assign _EVAL_248 = _EVAL_7 == 3'h4;
  assign _EVAL_120 = _EVAL == 3'h4;
  assign _EVAL_122 = _EVAL_113 | _EVAL_6;
  assign _EVAL_147 = _EVAL_40 | _EVAL_6;
  assign _EVAL_71 = _EVAL_106 | _EVAL_208;
  assign _EVAL_211 = ~_EVAL_70;
  assign _EVAL_210 = _EVAL_253 | _EVAL_120;
  assign _EVAL_86 = _EVAL_50 | _EVAL_6;
  assign _EVAL_68 = _EVAL_28 == 6'h0;
  assign _EVAL_296 = _EVAL_27 | _EVAL_6;
  assign _EVAL_253 = _EVAL_114 | _EVAL_25;
  assign _EVAL_95 = _EVAL_7[0];
  assign _EVAL_60 = ~_EVAL_203;
  assign _EVAL_208 = plusarg_reader_out == 32'h0;
  assign _EVAL_82 = ~_EVAL_290;
  assign _EVAL_203 = _EVAL_110 | _EVAL_6;
  assign _EVAL_112 = _EVAL_2[0];
  assign _EVAL_27 = _EVAL_5 == _EVAL_190;
  assign _EVAL_263 = ~_EVAL_42;
  assign _EVAL_100 = ~_EVAL_171;
  assign _EVAL_117 = ~_EVAL_3;
  assign _EVAL_284 = _EVAL_12 & _EVAL_220;
  assign _EVAL_133 = _EVAL_16 == _EVAL_216;
  assign _EVAL_63 = _EVAL_149 | _EVAL_6;
  assign _EVAL_174 = {_EVAL_151,_EVAL_51,_EVAL_213,_EVAL_283};
  assign _EVAL_226 = {{6'd0}, _EVAL_148};
  assign _EVAL_201 = _EVAL_15 == _EVAL_258;
  assign _EVAL_78 = _EVAL_259 | _EVAL_6;
  assign _EVAL_282 = _EVAL_12 & _EVAL_248;
  assign _EVAL_140 = _EVAL_58 == 2'h0;
  assign _EVAL_131 = ~_EVAL_57;
  assign _EVAL_218 = _EVAL_295[7:0];
  assign _EVAL_90 = _EVAL_14 & _EVAL_189;
  assign _EVAL_115 = _EVAL_270 | _EVAL_124;
  assign _EVAL_137 = _EVAL_286 & _EVAL_249;
  assign _EVAL_234 = _EVAL_299 | _EVAL_41;
  assign _EVAL_52 = _EVAL_5 != 3'h0;
  assign _EVAL_155 = _EVAL_37 >> _EVAL;
  assign _EVAL_267 = $signed(_EVAL_73) & -15'sh1000;
  assign _EVAL_175 = ~_EVAL_262;
  assign _EVAL_37 = _EVAL_41 | _EVAL_299;
  assign _EVAL_176 = _EVAL_13 >= 4'h2;
  assign _EVAL_189 = ~_EVAL_174;
  assign _EVAL_64 = _EVAL_182 + 32'h1;
  assign _EVAL_167 = ~_EVAL_156;
  assign _EVAL_283 = _EVAL_255 | _EVAL_111;
  assign _EVAL_195 = _EVAL_7 == _EVAL_223;
  assign _EVAL_297 = _EVAL_12 & _EVAL_136;
  assign _EVAL_127 = _EVAL_227 | _EVAL_6;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_21 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_28 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_54 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_59 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_94 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_116 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_126 = _RAND_6[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_163 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_182 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_190 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_214 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_216 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_223 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_233 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_258 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_280 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_299 = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_11) begin
    if (_EVAL_181) begin
      _EVAL_21 <= _EVAL;
    end
    if (_EVAL_6) begin
      _EVAL_28 <= 6'h0;
    end else if (_EVAL_238) begin
      if (_EVAL_68) begin
        if (_EVAL_95) begin
          _EVAL_28 <= _EVAL_153;
        end else begin
          _EVAL_28 <= 6'h0;
        end
      end else begin
        _EVAL_28 <= _EVAL_125;
      end
    end
    if (_EVAL_6) begin
      _EVAL_54 <= 6'h0;
    end else if (_EVAL_238) begin
      if (_EVAL_292) begin
        if (_EVAL_95) begin
          _EVAL_54 <= _EVAL_153;
        end else begin
          _EVAL_54 <= 6'h0;
        end
      end else begin
        _EVAL_54 <= _EVAL_141;
      end
    end
    if (_EVAL_181) begin
      _EVAL_59 <= _EVAL_4;
    end
    if (_EVAL_6) begin
      _EVAL_94 <= 6'h0;
    end else if (_EVAL_178) begin
      if (_EVAL_185) begin
        if (_EVAL_256) begin
          _EVAL_94 <= _EVAL_24;
        end else begin
          _EVAL_94 <= 6'h0;
        end
      end else begin
        _EVAL_94 <= _EVAL_241;
      end
    end
    if (_EVAL_181) begin
      _EVAL_116 <= _EVAL_0;
    end
    if (_EVAL_143) begin
      _EVAL_126 <= _EVAL_2;
    end
    if (_EVAL_181) begin
      _EVAL_163 <= _EVAL_9;
    end
    if (_EVAL_6) begin
      _EVAL_182 <= 32'h0;
    end else if (_EVAL_93) begin
      _EVAL_182 <= 32'h0;
    end else begin
      _EVAL_182 <= _EVAL_235;
    end
    if (_EVAL_143) begin
      _EVAL_190 <= _EVAL_5;
    end
    if (_EVAL_6) begin
      _EVAL_214 <= 6'h0;
    end else if (_EVAL_178) begin
      if (_EVAL_196) begin
        if (_EVAL_256) begin
          _EVAL_214 <= _EVAL_24;
        end else begin
          _EVAL_214 <= 6'h0;
        end
      end else begin
        _EVAL_214 <= _EVAL_169;
      end
    end
    if (_EVAL_143) begin
      _EVAL_216 <= _EVAL_16;
    end
    if (_EVAL_181) begin
      _EVAL_223 <= _EVAL_7;
    end
    if (_EVAL_143) begin
      _EVAL_233 <= _EVAL_17;
    end
    if (_EVAL_143) begin
      _EVAL_258 <= _EVAL_15;
    end
    if (_EVAL_181) begin
      _EVAL_280 <= _EVAL_13;
    end
    if (_EVAL_6) begin
      _EVAL_299 <= 5'h0;
    end else begin
      _EVAL_299 <= _EVAL_269;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16035bba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1d4d4de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3cd76ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6600093)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b483d81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44065d6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c8b4e35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_211) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b109093e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7641805b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33f2bb39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(754d77ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ebdd70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cedcd6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c009526)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e008bad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73b86229)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8db2b9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7307629)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cc1288a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7de07ba9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7747464)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83c7a0ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59fbd93c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48438429)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c633b442)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83ee08f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_240) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51c517e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0438ece)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(705b9f2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b196ad8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bcf011f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1801ab97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bfb9c99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33a02578)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf471f81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5b8d5c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61f15133)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fea3ffc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69316254)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e06df185)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18101297)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(242bad5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e69b2676)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfbc6cac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6609087)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5814e3c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(523dedc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d474fa9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e478dbe4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fea0a420)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b96d5a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ae235de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e91a13b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_211) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7034c5a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15278994)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a80aedb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97501406)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a61c207)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87d20865)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48d5f826)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa207680)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a32bd95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(505218d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13ebe3df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bde3e9d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52d3a646)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4befdaf3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54115758)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_240) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(723bef08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ac78b63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(108c62c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a745e020)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ee057e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5719096b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(805261d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7b0912b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc2a51df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4078c87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(851a4fc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d16ef88b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f326f456)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8893c3fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4fafe02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(713346e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1970ecae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84f0f370)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a770bdc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9e24d41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85ba1920)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_297 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(473195d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0dc638a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
