//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_134(
  output [2:0]  _EVAL,
  input  [8:0]  _EVAL_0,
  input  [31:0] _EVAL_1,
  output        _EVAL_2,
  output        _EVAL_3,
  output [8:0]  _EVAL_4,
  output [31:0] _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  output        _EVAL_8,
  input         _EVAL_9,
  output [1:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  input         _EVAL_12,
  output        _EVAL_13,
  input         _EVAL_14,
  input  [3:0]  _EVAL_15,
  input         _EVAL_16,
  input  [31:0] _EVAL_17,
  output        _EVAL_18,
  output [31:0] _EVAL_19,
  input  [1:0]  _EVAL_20,
  output [3:0]  _EVAL_21,
  output [2:0]  _EVAL_22,
  output [1:0]  _EVAL_23,
  output        _EVAL_24,
  input  [2:0]  _EVAL_25,
  output        _EVAL_26,
  output        _EVAL_27,
  input         _EVAL_28
);
  wire  AsyncQueueSource__EVAL;
  wire [31:0] AsyncQueueSource__EVAL_0;
  wire  AsyncQueueSource__EVAL_1;
  wire  AsyncQueueSource__EVAL_2;
  wire [8:0] AsyncQueueSource__EVAL_3;
  wire [8:0] AsyncQueueSource__EVAL_4;
  wire  AsyncQueueSource__EVAL_5;
  wire  AsyncQueueSource__EVAL_6;
  wire [2:0] AsyncQueueSource__EVAL_7;
  wire [3:0] AsyncQueueSource__EVAL_8;
  wire [3:0] AsyncQueueSource__EVAL_9;
  wire [31:0] AsyncQueueSource__EVAL_10;
  wire  AsyncQueueSource__EVAL_11;
  wire [2:0] AsyncQueueSource__EVAL_12;
  wire  AsyncQueueSink__EVAL;
  wire [1:0] AsyncQueueSink__EVAL_0;
  wire  AsyncQueueSink__EVAL_1;
  wire  AsyncQueueSink__EVAL_2;
  wire  AsyncQueueSink__EVAL_3;
  wire [2:0] AsyncQueueSink__EVAL_4;
  wire [31:0] AsyncQueueSink__EVAL_5;
  wire [1:0] AsyncQueueSink__EVAL_6;
  wire  AsyncQueueSink__EVAL_7;
  wire  AsyncQueueSink__EVAL_8;
  wire [1:0] AsyncQueueSink__EVAL_9;
  wire  AsyncQueueSink__EVAL_10;
  wire [2:0] AsyncQueueSink__EVAL_11;
  wire [31:0] AsyncQueueSink__EVAL_12;
  wire  AsyncQueueSink__EVAL_13;
  wire  AsyncQueueSink__EVAL_14;
  wire  AsyncQueueSink__EVAL_15;
  wire  AsyncQueueSink__EVAL_16;
  _EVAL_131 AsyncQueueSource (
    ._EVAL(AsyncQueueSource__EVAL),
    ._EVAL_0(AsyncQueueSource__EVAL_0),
    ._EVAL_1(AsyncQueueSource__EVAL_1),
    ._EVAL_2(AsyncQueueSource__EVAL_2),
    ._EVAL_3(AsyncQueueSource__EVAL_3),
    ._EVAL_4(AsyncQueueSource__EVAL_4),
    ._EVAL_5(AsyncQueueSource__EVAL_5),
    ._EVAL_6(AsyncQueueSource__EVAL_6),
    ._EVAL_7(AsyncQueueSource__EVAL_7),
    ._EVAL_8(AsyncQueueSource__EVAL_8),
    ._EVAL_9(AsyncQueueSource__EVAL_9),
    ._EVAL_10(AsyncQueueSource__EVAL_10),
    ._EVAL_11(AsyncQueueSource__EVAL_11),
    ._EVAL_12(AsyncQueueSource__EVAL_12)
  );
  _EVAL_133 AsyncQueueSink (
    ._EVAL(AsyncQueueSink__EVAL),
    ._EVAL_0(AsyncQueueSink__EVAL_0),
    ._EVAL_1(AsyncQueueSink__EVAL_1),
    ._EVAL_2(AsyncQueueSink__EVAL_2),
    ._EVAL_3(AsyncQueueSink__EVAL_3),
    ._EVAL_4(AsyncQueueSink__EVAL_4),
    ._EVAL_5(AsyncQueueSink__EVAL_5),
    ._EVAL_6(AsyncQueueSink__EVAL_6),
    ._EVAL_7(AsyncQueueSink__EVAL_7),
    ._EVAL_8(AsyncQueueSink__EVAL_8),
    ._EVAL_9(AsyncQueueSink__EVAL_9),
    ._EVAL_10(AsyncQueueSink__EVAL_10),
    ._EVAL_11(AsyncQueueSink__EVAL_11),
    ._EVAL_12(AsyncQueueSink__EVAL_12),
    ._EVAL_13(AsyncQueueSink__EVAL_13),
    ._EVAL_14(AsyncQueueSink__EVAL_14),
    ._EVAL_15(AsyncQueueSink__EVAL_15),
    ._EVAL_16(AsyncQueueSink__EVAL_16)
  );
  assign AsyncQueueSink__EVAL_6 = _EVAL_20;
  assign _EVAL_10 = AsyncQueueSink__EVAL_9;
  assign _EVAL_27 = AsyncQueueSink__EVAL_15;
  assign _EVAL_4 = AsyncQueueSource__EVAL_3;
  assign AsyncQueueSource__EVAL_11 = _EVAL_6;
  assign _EVAL_24 = AsyncQueueSink__EVAL_10;
  assign _EVAL = AsyncQueueSink__EVAL_11;
  assign AsyncQueueSource__EVAL = _EVAL_28;
  assign _EVAL_23 = AsyncQueueSink__EVAL_0;
  assign AsyncQueueSink__EVAL_1 = _EVAL_7;
  assign _EVAL_13 = AsyncQueueSink__EVAL_3;
  assign AsyncQueueSink__EVAL_8 = _EVAL_14;
  assign AsyncQueueSink__EVAL_16 = _EVAL_12;
  assign AsyncQueueSource__EVAL_9 = _EVAL_15;
  assign _EVAL_8 = AsyncQueueSource__EVAL_2;
  assign AsyncQueueSource__EVAL_6 = _EVAL_16;
  assign AsyncQueueSource__EVAL_10 = _EVAL_17;
  assign _EVAL_22 = AsyncQueueSource__EVAL_7;
  assign AsyncQueueSink__EVAL_5 = _EVAL_1;
  assign _EVAL_26 = AsyncQueueSink__EVAL_14;
  assign AsyncQueueSource__EVAL_12 = _EVAL_11;
  assign _EVAL_3 = AsyncQueueSource__EVAL_5;
  assign _EVAL_2 = AsyncQueueSink__EVAL_7;
  assign _EVAL_18 = AsyncQueueSink__EVAL_13;
  assign _EVAL_21 = AsyncQueueSource__EVAL_8;
  assign AsyncQueueSink__EVAL = _EVAL_9;
  assign AsyncQueueSource__EVAL_1 = _EVAL_7;
  assign AsyncQueueSink__EVAL_2 = _EVAL_16;
  assign AsyncQueueSink__EVAL_4 = _EVAL_25;
  assign _EVAL_19 = AsyncQueueSink__EVAL_12;
  assign _EVAL_5 = AsyncQueueSource__EVAL_0;
  assign AsyncQueueSource__EVAL_4 = _EVAL_0;
endmodule
