//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_31_assert(
  input  [2:0]  _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [3:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [1:0]  _EVAL_12,
  input  [3:0]  _EVAL_13,
  input         _EVAL_14,
  input  [2:0]  _EVAL_15,
  input  [29:0] _EVAL_16,
  input         _EVAL_17,
  input  [3:0]  _EVAL_18
);
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  reg [31:0] _EVAL_22;
  reg [31:0] _RAND_0;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire [29:0] _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire [3:0] _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire [1:0] _EVAL_35;
  wire [1:0] _EVAL_36;
  wire  _EVAL_37;
  wire [30:0] _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire [4:0] _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire [7:0] _EVAL_56;
  wire  _EVAL_57;
  wire [4:0] _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire [5:0] _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  reg [5:0] _EVAL_72;
  reg [31:0] _RAND_1;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire [29:0] _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  reg [1:0] _EVAL_90;
  reg [31:0] _RAND_2;
  wire  _EVAL_91;
  wire [29:0] _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire [30:0] _EVAL_101;
  wire  _EVAL_102;
  wire [6:0] _EVAL_103;
  wire [30:0] _EVAL_104;
  wire  _EVAL_105;
  wire [7:0] _EVAL_106;
  wire  _EVAL_107;
  wire [7:0] _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire [5:0] _EVAL_112;
  wire [3:0] _EVAL_113;
  wire [4:0] _EVAL_114;
  reg [29:0] _EVAL_115;
  reg [31:0] _RAND_3;
  wire  _EVAL_116;
  wire [29:0] _EVAL_117;
  wire  _EVAL_118;
  wire [30:0] _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire [4:0] _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  reg [2:0] _EVAL_153;
  reg [31:0] _RAND_4;
  wire  _EVAL_154;
  wire [3:0] _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire [29:0] _EVAL_159;
  reg [2:0] _EVAL_160;
  reg [31:0] _RAND_5;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire [30:0] _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire [22:0] _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  reg [5:0] _EVAL_175;
  reg [31:0] _RAND_6;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire [30:0] _EVAL_178;
  wire [7:0] _EVAL_179;
  wire [6:0] _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  reg [2:0] _EVAL_185;
  reg [31:0] _RAND_7;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  reg  _EVAL_197;
  reg [31:0] _RAND_8;
  wire  _EVAL_198;
  wire [32:0] _EVAL_199;
  wire [30:0] _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire [5:0] _EVAL_216;
  reg [4:0] _EVAL_217;
  reg [31:0] _RAND_9;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire [4:0] _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire [30:0] _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire [7:0] _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire [31:0] plusarg_reader_out;
  reg [3:0] _EVAL_234;
  reg [31:0] _RAND_10;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  reg [5:0] _EVAL_245;
  reg [31:0] _RAND_11;
  wire  _EVAL_246;
  wire [31:0] _EVAL_248;
  reg  _EVAL_249;
  reg [31:0] _RAND_12;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_253;
  wire [6:0] _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire [4:0] _EVAL_258;
  wire  _EVAL_259;
  wire [7:0] _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  reg [3:0] _EVAL_263;
  reg [31:0] _RAND_13;
  wire  _EVAL_264;
  wire  _EVAL_265;
  reg [2:0] _EVAL_266;
  reg [31:0] _RAND_14;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  reg [5:0] _EVAL_270;
  reg [31:0] _RAND_15;
  wire [7:0] _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire [5:0] _EVAL_275;
  wire [30:0] _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire [22:0] _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire [4:0] _EVAL_283;
  wire [4:0] _EVAL_284;
  reg [2:0] _EVAL_285;
  reg [31:0] _RAND_16;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire [5:0] _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire [3:0] _EVAL_299;
  wire [30:0] _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire [30:0] _EVAL_311;
  wire [7:0] _EVAL_312;
  wire [30:0] _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire [1:0] _EVAL_316;
  wire [5:0] _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire  _EVAL_321;
  wire  _EVAL_322;
  wire [1:0] _EVAL_323;
  wire  _EVAL_324;
  wire  _EVAL_325;
  wire [6:0] _EVAL_326;
  wire  _EVAL_327;
  wire  _EVAL_328;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_161 = _EVAL_127[0];
  assign _EVAL_87 = _EVAL_5 >= 4'h2;
  assign _EVAL_246 = plusarg_reader_out == 32'h0;
  assign _EVAL_193 = ~_EVAL_10;
  assign _EVAL_159 = _EVAL_16 ^ 30'h20000000;
  assign _EVAL_224 = _EVAL_68 | _EVAL_9;
  assign _EVAL_35 = _EVAL_15[2:1];
  assign _EVAL_117 = _EVAL_16 ^ 30'h2000000;
  assign _EVAL_322 = _EVAL_6[2];
  assign _EVAL_147 = _EVAL_148 | _EVAL_9;
  assign _EVAL_239 = _EVAL_264 | _EVAL_172;
  assign _EVAL_293 = ~_EVAL_83;
  assign _EVAL_21 = _EVAL_51 != 5'h0;
  assign _EVAL_210 = ~_EVAL_19;
  assign _EVAL_273 = _EVAL_0 == 3'h2;
  assign _EVAL_83 = _EVAL_63 | _EVAL_9;
  assign _EVAL_158 = _EVAL_302 | _EVAL_107;
  assign _EVAL_106 = 8'h1 << _EVAL;
  assign _EVAL_201 = ~_EVAL_309;
  assign _EVAL_142 = _EVAL_14 & _EVAL_286;
  assign _EVAL_171 = 23'hff << _EVAL_5;
  assign _EVAL_74 = _EVAL_149 & _EVAL_32;
  assign _EVAL_116 = _EVAL_109 | _EVAL_9;
  assign _EVAL_44 = _EVAL_6 == 3'h5;
  assign _EVAL_25 = _EVAL_16 & _EVAL_92;
  assign _EVAL_99 = ~_EVAL_181;
  assign _EVAL_139 = _EVAL_16[0];
  assign _EVAL_323 = 2'h1 << _EVAL_218;
  assign _EVAL_324 = _EVAL_43 | _EVAL_320;
  assign _EVAL_89 = _EVAL_42 | _EVAL_9;
  assign _EVAL_103 = _EVAL_270 - 6'h1;
  assign _EVAL_237 = _EVAL_205 | _EVAL_321;
  assign _EVAL_306 = _EVAL_14 & _EVAL_213;
  assign _EVAL_181 = _EVAL_245 == 6'h0;
  assign _EVAL_123 = ~_EVAL_189;
  assign _EVAL_230 = _EVAL_187 ? _EVAL_260 : 8'h0;
  assign _EVAL_219 = _EVAL_195 & _EVAL_139;
  assign _EVAL_95 = $signed(_EVAL_104) == 31'sh0;
  assign _EVAL_108 = ~_EVAL_312;
  assign _EVAL_88 = _EVAL_164 | _EVAL_9;
  assign _EVAL_218 = _EVAL_5[0];
  assign _EVAL_110 = ~_EVAL_303;
  assign _EVAL_101 = $signed(_EVAL_226) & -31'sh1000;
  assign _EVAL_145 = _EVAL_66 | _EVAL_9;
  assign _EVAL_144 = _EVAL_41 | _EVAL_9;
  assign _EVAL_192 = _EVAL_8 & _EVAL_273;
  assign _EVAL_275 = _EVAL_254[5:0];
  assign _EVAL_178 = {1'b0,$signed(_EVAL_159)};
  assign _EVAL_292 = _EVAL_75 | _EVAL_10;
  assign _EVAL_315 = _EVAL_149 & _EVAL_219;
  assign _EVAL_62 = _EVAL_113 == 4'h0;
  assign _EVAL_213 = _EVAL_6 == 3'h6;
  assign _EVAL_327 = ~_EVAL_168;
  assign _EVAL_81 = _EVAL_203 | _EVAL_9;
  assign _EVAL_29 = ~_EVAL_54;
  assign _EVAL_124 = ~_EVAL_166;
  assign _EVAL_291 = _EVAL_108[7:2];
  assign _EVAL_135 = _EVAL_149 & _EVAL_294;
  assign _EVAL_229 = _EVAL_0 <= 3'h6;
  assign _EVAL_325 = ~_EVAL_88;
  assign _EVAL_251 = _EVAL_320 & _EVAL_181;
  assign _EVAL_163 = ~_EVAL_314;
  assign _EVAL_200 = {1'b0,$signed(_EVAL_16)};
  assign _EVAL_111 = _EVAL_36[1];
  assign _EVAL_42 = _EVAL_28 == 4'h0;
  assign _EVAL_269 = _EVAL_43 & _EVAL_169;
  assign _EVAL_126 = _EVAL_111 & _EVAL_319;
  assign _EVAL_208 = _EVAL_231 | _EVAL_136;
  assign _EVAL_262 = _EVAL_137 | _EVAL_9;
  assign _EVAL_286 = ~_EVAL_152;
  assign _EVAL_281 = _EVAL_71 | _EVAL_9;
  assign _EVAL_130 = _EVAL_8 & _EVAL_257;
  assign _EVAL_146 = $signed(_EVAL_119) == 31'sh0;
  assign _EVAL_206 = ~_EVAL_64;
  assign _EVAL_290 = _EVAL_7 == _EVAL_249;
  assign _EVAL_272 = _EVAL_39 | _EVAL_246;
  assign _EVAL_250 = _EVAL_217 != 5'h0;
  assign _EVAL_70 = ~_EVAL_223;
  assign _EVAL_143 = _EVAL_0 == 3'h4;
  assign _EVAL_156 = {_EVAL_204,_EVAL_207,_EVAL_242,_EVAL_328};
  assign _EVAL_125 = _EVAL_18 == _EVAL_156;
  assign _EVAL_67 = _EVAL_4 == _EVAL_285;
  assign _EVAL_274 = ~_EVAL_211;
  assign _EVAL_127 = _EVAL_284 >> _EVAL_15;
  assign _EVAL_24 = ~_EVAL_3;
  assign _EVAL_19 = _EVAL_277 | _EVAL_9;
  assign _EVAL_204 = _EVAL_308 | _EVAL_135;
  assign _EVAL_66 = _EVAL_4 <= 3'h3;
  assign _EVAL_112 = _EVAL_180[5:0];
  assign _EVAL_300 = _EVAL_276;
  assign _EVAL_47 = _EVAL_55 | _EVAL_146;
  assign _EVAL_45 = ~_EVAL_261;
  assign _EVAL_326 = _EVAL_175 - 6'h1;
  assign _EVAL_34 = _EVAL_6 == 3'h3;
  assign _EVAL_312 = _EVAL_279[7:0];
  assign _EVAL_57 = ~_EVAL_183;
  assign _EVAL_148 = _EVAL_4 <= 3'h1;
  assign _EVAL_174 = _EVAL_73 | _EVAL_9;
  assign _EVAL_32 = _EVAL_319 & _EVAL_84;
  assign _EVAL_65 = _EVAL_13 >= 4'h2;
  assign _EVAL_259 = ~_EVAL_102;
  assign _EVAL_241 = _EVAL_6 == _EVAL_266;
  assign _EVAL_30 = _EVAL_190 & _EVAL_47;
  assign _EVAL_278 = _EVAL_8 & _EVAL_99;
  assign _EVAL_187 = _EVAL_280 & _EVAL_327;
  assign _EVAL_170 = _EVAL_0 == 3'h1;
  assign _EVAL_209 = _EVAL_48 | _EVAL_9;
  assign _EVAL_94 = _EVAL_0 == 3'h0;
  assign _EVAL_260 = 8'h1 << _EVAL_15;
  assign _EVAL_162 = _EVAL_158 | _EVAL_9;
  assign _EVAL_316 = _EVAL[2:1];
  assign _EVAL_309 = _EVAL_290 | _EVAL_9;
  assign _EVAL_191 = _EVAL_173 | _EVAL_9;
  assign _EVAL_307 = _EVAL_0[0];
  assign _EVAL_228 = _EVAL_22 < plusarg_reader_out;
  assign _EVAL_182 = ~_EVAL_9;
  assign _EVAL_68 = _EVAL_25 == 30'h0;
  assign _EVAL_248 = _EVAL_199[31:0];
  assign _EVAL_52 = $signed(_EVAL_311) == 31'sh0;
  assign _EVAL_152 = _EVAL_270 == 6'h0;
  assign _EVAL_71 = _EVAL_4 <= 3'h4;
  assign _EVAL_253 = _EVAL_30 | _EVAL_9;
  assign _EVAL_226 = {1'b0,$signed(_EVAL_78)};
  assign _EVAL_169 = _EVAL_72 == 6'h0;
  assign _EVAL_102 = _EVAL_208 | _EVAL_9;
  assign _EVAL_294 = _EVAL_319 & _EVAL_139;
  assign _EVAL_222 = _EVAL_8 & _EVAL_94;
  assign _EVAL_186 = ~_EVAL_157;
  assign _EVAL_119 = _EVAL_38;
  assign _EVAL_282 = _EVAL_62 | _EVAL_9;
  assign _EVAL_256 = ~_EVAL_282;
  assign _EVAL_46 = _EVAL_12 != 2'h2;
  assign _EVAL_231 = _EVAL_265 & _EVAL_52;
  assign _EVAL_128 = _EVAL_4 == 3'h0;
  assign _EVAL_36 = _EVAL_323 | 2'h1;
  assign _EVAL_176 = ~_EVAL_162;
  assign _EVAL_73 = _EVAL_272 | _EVAL_228;
  assign _EVAL_132 = ~_EVAL_227;
  assign _EVAL_180 = _EVAL_245 - 6'h1;
  assign _EVAL_98 = ~_EVAL_224;
  assign _EVAL_79 = _EVAL_85 | _EVAL_95;
  assign _EVAL_58 = _EVAL_217 >> _EVAL;
  assign _EVAL_308 = _EVAL_87 | _EVAL_126;
  assign _EVAL_299 = ~_EVAL_156;
  assign _EVAL_212 = _EVAL_149 & _EVAL_298;
  assign _EVAL_223 = _EVAL_241 | _EVAL_9;
  assign _EVAL_164 = _EVAL_237 | _EVAL_198;
  assign _EVAL_319 = _EVAL_16[1];
  assign _EVAL_267 = ~_EVAL_89;
  assign _EVAL_55 = _EVAL_297 | _EVAL_95;
  assign _EVAL_33 = _EVAL_215 | _EVAL_9;
  assign _EVAL_214 = _EVAL_14 & _EVAL_105;
  assign _EVAL_91 = _EVAL_8 & _EVAL_170;
  assign _EVAL_172 = _EVAL_35 == 2'h0;
  assign _EVAL_216 = _EVAL_271[7:2];
  assign _EVAL_305 = ~_EVAL_253;
  assign _EVAL_167 = _EVAL_79 | _EVAL_146;
  assign _EVAL_321 = _EVAL_316 == 2'h0;
  assign _EVAL_221 = ~_EVAL_81;
  assign _EVAL_189 = _EVAL_65 | _EVAL_9;
  assign _EVAL_75 = ~_EVAL_11;
  assign _EVAL_137 = _EVAL_0 == _EVAL_153;
  assign _EVAL_328 = _EVAL_141 | _EVAL_212;
  assign _EVAL_165 = $signed(_EVAL_200) & -31'sh5000;
  assign _EVAL_43 = _EVAL_1 & _EVAL_14;
  assign _EVAL_283 = _EVAL_230[4:0];
  assign _EVAL_28 = ~_EVAL_18;
  assign _EVAL_76 = ~_EVAL_184;
  assign _EVAL_120 = ~_EVAL_177;
  assign _EVAL_311 = _EVAL_101;
  assign _EVAL_296 = ~_EVAL_20;
  assign _EVAL_92 = {{22'd0}, _EVAL_271};
  assign _EVAL_177 = _EVAL_292 | _EVAL_9;
  assign _EVAL_255 = ~_EVAL_154;
  assign _EVAL_151 = ~_EVAL_262;
  assign _EVAL_276 = $signed(_EVAL_313) & -31'sh1000000;
  assign _EVAL_105 = _EVAL_6 == 3'h0;
  assign _EVAL_233 = ~_EVAL_304;
  assign _EVAL_168 = _EVAL_0 == 3'h6;
  assign _EVAL_264 = _EVAL_35 == 2'h1;
  assign _EVAL_39 = ~_EVAL_250;
  assign _EVAL_84 = ~_EVAL_139;
  assign _EVAL_38 = $signed(_EVAL_178) & -31'sh2000;
  assign _EVAL_64 = _EVAL_133 | _EVAL_9;
  assign _EVAL_49 = ~_EVAL_131;
  assign _EVAL_302 = _EVAL_51 != _EVAL_283;
  assign _EVAL_280 = _EVAL_320 & _EVAL_236;
  assign _EVAL_254 = _EVAL_72 - 6'h1;
  assign _EVAL_114 = ~_EVAL_283;
  assign _EVAL_133 = _EVAL_4 <= 3'h2;
  assign _EVAL_284 = _EVAL_51 | _EVAL_217;
  assign _EVAL_136 = _EVAL_190 & _EVAL_146;
  assign _EVAL_314 = _EVAL_24 | _EVAL_9;
  assign _EVAL_134 = _EVAL_6 == 3'h1;
  assign _EVAL_179 = _EVAL_269 ? _EVAL_106 : 8'h0;
  assign _EVAL_257 = _EVAL_0 == 3'h5;
  assign _EVAL_184 = _EVAL_128 | _EVAL_9;
  assign _EVAL_195 = ~_EVAL_319;
  assign _EVAL_227 = _EVAL_287 | _EVAL_9;
  assign _EVAL_205 = _EVAL_316 == 2'h1;
  assign _EVAL_295 = _EVAL_13 == _EVAL_263;
  assign _EVAL_258 = _EVAL_217 | _EVAL_51;
  assign _EVAL_243 = ~_EVAL_144;
  assign _EVAL_289 = ~_EVAL_33;
  assign _EVAL_297 = _EVAL_52 | _EVAL_85;
  assign _EVAL_54 = _EVAL_240 | _EVAL_9;
  assign _EVAL_27 = ~_EVAL_281;
  assign _EVAL_183 = _EVAL_125 | _EVAL_9;
  assign _EVAL_59 = _EVAL_14 & _EVAL_44;
  assign _EVAL_287 = _EVAL == _EVAL_160;
  assign _EVAL_140 = ~_EVAL_147;
  assign _EVAL_77 = _EVAL_58[0];
  assign _EVAL_261 = _EVAL_23 | _EVAL_9;
  assign _EVAL_242 = _EVAL_141 | _EVAL_315;
  assign _EVAL_150 = _EVAL_8 & _EVAL_143;
  assign _EVAL_26 = _EVAL_14 & _EVAL_34;
  assign _EVAL_298 = _EVAL_195 & _EVAL_84;
  assign _EVAL_190 = _EVAL_5 <= 4'h2;
  assign _EVAL_279 = 23'hff << _EVAL_13;
  assign _EVAL_121 = _EVAL_6 == 3'h2;
  assign _EVAL_109 = ~_EVAL_77;
  assign _EVAL_303 = _EVAL_235 | _EVAL_9;
  assign _EVAL_23 = _EVAL_12 <= 2'h2;
  assign _EVAL_51 = _EVAL_179[4:0];
  assign _EVAL_97 = ~_EVAL_145;
  assign _EVAL_194 = _EVAL_6 == 3'h7;
  assign _EVAL_225 = _EVAL_190 & _EVAL_167;
  assign _EVAL_53 = _EVAL_190 & _EVAL_79;
  assign _EVAL_60 = ~_EVAL_209;
  assign _EVAL_207 = _EVAL_308 | _EVAL_74;
  assign _EVAL_215 = _EVAL_11 == _EVAL_197;
  assign _EVAL_104 = _EVAL_165;
  assign _EVAL_173 = _EVAL_239 | _EVAL_40;
  assign _EVAL_238 = _EVAL_14 & _EVAL_134;
  assign _EVAL_48 = _EVAL_5 == _EVAL_234;
  assign _EVAL_196 = ~_EVAL_202;
  assign _EVAL_232 = ~_EVAL_322;
  assign _EVAL_141 = _EVAL_87 | _EVAL_93;
  assign _EVAL_41 = _EVAL_12 == 2'h0;
  assign _EVAL_198 = _EVAL == 3'h4;
  assign _EVAL_318 = ~_EVAL_310;
  assign _EVAL_301 = _EVAL_14 & _EVAL_194;
  assign _EVAL_202 = _EVAL_161 | _EVAL_9;
  assign _EVAL_93 = _EVAL_111 & _EVAL_195;
  assign _EVAL_149 = _EVAL_36[0];
  assign _EVAL_240 = _EVAL_15 == _EVAL_185;
  assign _EVAL_203 = _EVAL_4 != 3'h0;
  assign _EVAL_20 = _EVAL_46 | _EVAL_9;
  assign _EVAL_69 = _EVAL_6 == 3'h4;
  assign _EVAL_78 = _EVAL_16 ^ 30'h3000;
  assign _EVAL_61 = _EVAL_326[5:0];
  assign _EVAL_277 = _EVAL_231 | _EVAL_53;
  assign _EVAL_265 = _EVAL_5 <= 4'h8;
  assign _EVAL_56 = _EVAL_171[7:0];
  assign _EVAL_82 = _EVAL_231 | _EVAL_225;
  assign _EVAL_268 = _EVAL_43 & _EVAL_152;
  assign _EVAL_40 = _EVAL_15 == 3'h4;
  assign _EVAL_199 = _EVAL_22 + 32'h1;
  assign _EVAL_113 = _EVAL_18 & _EVAL_299;
  assign _EVAL_320 = _EVAL_17 & _EVAL_8;
  assign _EVAL_310 = _EVAL_295 | _EVAL_9;
  assign _EVAL_244 = _EVAL_8 & _EVAL_168;
  assign _EVAL_271 = ~_EVAL_56;
  assign _EVAL_63 = _EVAL_12 == _EVAL_90;
  assign _EVAL_138 = ~_EVAL_116;
  assign _EVAL_317 = _EVAL_103[5:0];
  assign _EVAL_157 = _EVAL_75 | _EVAL_9;
  assign _EVAL_96 = _EVAL_14 & _EVAL_121;
  assign _EVAL_131 = _EVAL_82 | _EVAL_9;
  assign _EVAL_211 = _EVAL_229 | _EVAL_9;
  assign _EVAL_166 = _EVAL_67 | _EVAL_9;
  assign _EVAL_220 = _EVAL_258 & _EVAL_114;
  assign _EVAL_37 = _EVAL_14 & _EVAL_69;
  assign _EVAL_313 = {1'b0,$signed(_EVAL_117)};
  assign _EVAL_85 = $signed(_EVAL_300) == 31'sh0;
  assign _EVAL_154 = _EVAL_87 | _EVAL_9;
  assign _EVAL_118 = ~_EVAL_174;
  assign _EVAL_107 = ~_EVAL_21;
  assign _EVAL_235 = _EVAL_16 == _EVAL_115;
  assign _EVAL_304 = _EVAL_193 | _EVAL_9;
  assign _EVAL_100 = ~_EVAL_191;
  assign _EVAL_236 = _EVAL_175 == 6'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_22 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_72 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_90 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_115 = _RAND_3[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_153 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_160 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_175 = _RAND_6[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_185 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_197 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_217 = _RAND_9[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_234 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_245 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_249 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_263 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_266 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_270 = _RAND_15[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_285 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_2) begin
    if (_EVAL_9) begin
      _EVAL_22 <= 32'h0;
    end else if (_EVAL_324) begin
      _EVAL_22 <= 32'h0;
    end else begin
      _EVAL_22 <= _EVAL_248;
    end
    if (_EVAL_9) begin
      _EVAL_72 <= 6'h0;
    end else if (_EVAL_43) begin
      if (_EVAL_169) begin
        if (_EVAL_232) begin
          _EVAL_72 <= _EVAL_216;
        end else begin
          _EVAL_72 <= 6'h0;
        end
      end else begin
        _EVAL_72 <= _EVAL_275;
      end
    end
    if (_EVAL_251) begin
      _EVAL_90 <= _EVAL_12;
    end
    if (_EVAL_268) begin
      _EVAL_115 <= _EVAL_16;
    end
    if (_EVAL_251) begin
      _EVAL_153 <= _EVAL_0;
    end
    if (_EVAL_268) begin
      _EVAL_160 <= _EVAL;
    end
    if (_EVAL_9) begin
      _EVAL_175 <= 6'h0;
    end else if (_EVAL_320) begin
      if (_EVAL_236) begin
        if (_EVAL_307) begin
          _EVAL_175 <= _EVAL_291;
        end else begin
          _EVAL_175 <= 6'h0;
        end
      end else begin
        _EVAL_175 <= _EVAL_61;
      end
    end
    if (_EVAL_251) begin
      _EVAL_185 <= _EVAL_15;
    end
    if (_EVAL_251) begin
      _EVAL_197 <= _EVAL_11;
    end
    if (_EVAL_9) begin
      _EVAL_217 <= 5'h0;
    end else begin
      _EVAL_217 <= _EVAL_220;
    end
    if (_EVAL_268) begin
      _EVAL_234 <= _EVAL_5;
    end
    if (_EVAL_9) begin
      _EVAL_245 <= 6'h0;
    end else if (_EVAL_320) begin
      if (_EVAL_181) begin
        if (_EVAL_307) begin
          _EVAL_245 <= _EVAL_291;
        end else begin
          _EVAL_245 <= 6'h0;
        end
      end else begin
        _EVAL_245 <= _EVAL_112;
      end
    end
    if (_EVAL_251) begin
      _EVAL_249 <= _EVAL_7;
    end
    if (_EVAL_251) begin
      _EVAL_263 <= _EVAL_13;
    end
    if (_EVAL_268) begin
      _EVAL_266 <= _EVAL_6;
    end
    if (_EVAL_9) begin
      _EVAL_270 <= 6'h0;
    end else if (_EVAL_43) begin
      if (_EVAL_152) begin
        if (_EVAL_232) begin
          _EVAL_270 <= _EVAL_216;
        end else begin
          _EVAL_270 <= 6'h0;
        end
      end else begin
        _EVAL_270 <= _EVAL_317;
      end
    end
    if (_EVAL_268) begin
      _EVAL_285 <= _EVAL_4;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(284cd84c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_255) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d570b077)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_318) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_325) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7590f0ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26a98f31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d537fe04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(525211a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e027cde5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67d0105b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f70a8e92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c42778d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_325) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e60784a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec2abebe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9df9454)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3aff28cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(623579c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c59b7b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c9e9ed0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f9ff6e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33827917)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_325) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba34b342)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_305) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(474ebf8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(924db437)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd93d3b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c431e0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7135f0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2951cbf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1983cc91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49d4003d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87a49b09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7287d107)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c6c2e17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f87ac590)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34e32532)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4ae42ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_325) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64047657)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35327474)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_325) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f86db1a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bce2981)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c40694d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba7a6a4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1b14d8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc384e38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bb168e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3089b1df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f8b8f21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_325) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5a26738)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27ebfe9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_305) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_305) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9381c7ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5c5086f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_255) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35f0258)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73bb6104)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e23bdf8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7d9ba3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f201133e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_325) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c850e35e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_255) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6703368)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33e12083)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_325) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7400dd52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9938923)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_318) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(592a0218)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f557b4e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b58c0742)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_325) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83a2025a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93aaa186)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4028b1d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_325) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0c644af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(466786df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24063f72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_325) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_325) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32d88cc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(febdf8e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8970a1a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3325e1d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_8 & _EVAL_274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_325) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd46516c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_325) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d2a0754)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cc9c12f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec4f0de1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a6fccbf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16d5b89a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a63fd1ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_255) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adb618e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67d81002)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52b2d283)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_325) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91e284db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63f31ebf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ba6358)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_26 & _EVAL_305) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_8 & _EVAL_274) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f848b459)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(effb58ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b20b1fe4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1577048)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_325) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51fe5092)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_130 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8575024b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
