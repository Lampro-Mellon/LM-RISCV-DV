//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_141_assert(
  input          _EVAL,
  input  [2:0]   _EVAL_0,
  input          _EVAL_2,
  input  [2:0]   _EVAL_5,
  input  [2:0]   _EVAL_13,
  input  [1:0]   _EVAL_14,
  input  [2:0]   _EVAL_15,
  input          _EVAL_20,
  input  [8:0]   _EVAL_21,
  input  [31:0]  _EVAL_26,
  input  [3:0]   _EVAL_28,
  input  [3:0]   _EVAL_29,
  input          _EVAL_30,
  input          _EVAL_32,
  input          _EVAL_33,
  input          _EVAL_34,
  input  [11:0]  _EVAL_36,
  input          _EVAL_38,
  input  [2:0]   _EVAL_39,
  input  [1:0]   _EVAL_40,
  input          _EVAL_41,
  input  [31:0]  _EVAL_83,
  input          _EVAL_200,
  input          _EVAL_209,
  input          _EVAL_360,
  input          _EVAL_421,
  input          _EVAL_468,
  input          _EVAL_470,
  input          _EVAL_474,
  input  [31:0]  _EVAL_575,
  input  [1:0]   _EVAL_612,
  input          _EVAL_624,
  input          _EVAL_724,
  input          _EVAL_829,
  input          _EVAL_926,
  input          _EVAL_952,
  input          _EVAL_1049,
  input          _EVAL_1183,
  input          _EVAL_1184,
  input          _EVAL_1191,
  input          _EVAL_1335,
  input          _EVAL_1337,
  input          _EVAL_1376,
  input          _EVAL_1400,
  input          _EVAL_1523,
  input          _EVAL_1575,
  input          _EVAL_1589,
  input          _EVAL_1681,
  input          _EVAL_1752,
  input          _EVAL_1761,
  input          _EVAL_1830,
  input          _EVAL_1834,
  input          _EVAL_1841,
  input          _EVAL_1856,
  input          _EVAL_1871,
  input          _EVAL_1888,
  input          _EVAL_1897,
  input          _EVAL_1945,
  input  [1:0]   _EVAL_1987,
  input          _EVAL_2004,
  input          _EVAL_2018,
  input          _EVAL_2029,
  input          _EVAL_2061,
  input          _EVAL_2188,
  input          _EVAL_2262,
  input  [31:0]  _EVAL_2363,
  input          _EVAL_2400,
  input          _EVAL_2488,
  input          _EVAL_2499,
  input          _EVAL_2571,
  input          _EVAL_2583,
  input          _EVAL_2594,
  input  [2:0]   _EVAL_2628,
  input          _EVAL_2643,
  input          _EVAL_2651,
  input          _EVAL_2655,
  input  [7:0]   _EVAL_2662,
  input          _EVAL_2714,
  input  [511:0] _EVAL_2743,
  input          _EVAL_2828,
  input          _EVAL_2845,
  input  [7:0]   _EVAL_2864,
  input          _EVAL_2988,
  input          _EVAL_3155,
  input          _EVAL_3264,
  input          _EVAL_3268,
  input          _EVAL_3425,
  input  [7:0]   _EVAL_3474,
  input          _EVAL_3485,
  input          _EVAL_3507,
  input          _EVAL_3519,
  input          _EVAL_3588,
  input          _EVAL_3670,
  input          _EVAL_3701,
  input  [7:0]   _EVAL_3750,
  input          _EVAL_3836
);
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_50;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_57;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_62;
  wire  _EVAL_64;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_77;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_89;
  wire  _EVAL_91;
  wire  _EVAL_96;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_112;
  wire  _EVAL_114;
  wire  _EVAL_116;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_122;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_140;
  wire  _EVAL_142;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_155;
  wire  _EVAL_157;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_168;
  wire  _EVAL_170;
  wire  _EVAL_173;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_183;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_199;
  wire  _EVAL_201;
  wire  _EVAL_203;
  wire  _EVAL_208;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_213;
  wire  _EVAL_216;
  wire  _EVAL_218;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_224;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_235;
  wire  _EVAL_240;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_250;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_267;
  wire  _EVAL_269;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_281;
  wire  _EVAL_283;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_305;
  wire [2:0] _EVAL_307;
  wire [3:0] _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_321;
  wire  _EVAL_322;
  wire  _EVAL_326;
  wire  _EVAL_328;
  wire  _EVAL_330;
  wire  _EVAL_335;
  wire  _EVAL_336;
  wire  _EVAL_337;
  wire  _EVAL_338;
  wire  _EVAL_340;
  wire  _EVAL_341;
  wire  _EVAL_342;
  wire  _EVAL_345;
  wire  _EVAL_346;
  wire  _EVAL_348;
  wire  _EVAL_349;
  wire  _EVAL_350;
  wire  _EVAL_352;
  wire  _EVAL_355;
  wire  _EVAL_356;
  wire  _EVAL_357;
  wire  _EVAL_358;
  wire  _EVAL_359;
  wire  _EVAL_361;
  wire  _EVAL_364;
  wire  _EVAL_367;
  wire  _EVAL_369;
  wire  _EVAL_371;
  wire  _EVAL_373;
  wire  _EVAL_376;
  wire  _EVAL_379;
  wire  _EVAL_380;
  wire  _EVAL_381;
  wire  _EVAL_383;
  wire  _EVAL_385;
  wire  _EVAL_387;
  wire  _EVAL_388;
  wire  _EVAL_390;
  wire  _EVAL_391;
  wire  _EVAL_394;
  wire  _EVAL_396;
  wire  _EVAL_398;
  wire  _EVAL_400;
  wire  _EVAL_404;
  wire  _EVAL_405;
  wire  _EVAL_408;
  wire  _EVAL_410;
  wire  _EVAL_411;
  wire  _EVAL_413;
  wire  _EVAL_414;
  wire  _EVAL_416;
  wire  _EVAL_418;
  wire  _EVAL_422;
  wire  _EVAL_423;
  wire  _EVAL_424;
  wire  _EVAL_425;
  wire  _EVAL_426;
  wire  _EVAL_427;
  wire  _EVAL_428;
  wire  _EVAL_429;
  wire  _EVAL_430;
  wire  _EVAL_433;
  wire  _EVAL_435;
  wire  _EVAL_437;
  wire  _EVAL_438;
  wire  _EVAL_440;
  wire  _EVAL_441;
  wire  _EVAL_443;
  wire  _EVAL_444;
  wire  _EVAL_445;
  wire  _EVAL_446;
  wire  _EVAL_447;
  wire  _EVAL_449;
  wire  _EVAL_452;
  wire  _EVAL_453;
  wire  _EVAL_454;
  wire  _EVAL_455;
  wire  _EVAL_456;
  wire  _EVAL_457;
  wire  _EVAL_460;
  wire  _EVAL_461;
  wire  _EVAL_462;
  wire  _EVAL_465;
  wire  _EVAL_466;
  wire  TLMonitor_1__EVAL;
  wire  TLMonitor_1__EVAL_0;
  wire  TLMonitor_1__EVAL_1;
  wire  TLMonitor_1__EVAL_2;
  wire [3:0] TLMonitor_1__EVAL_3;
  wire [2:0] TLMonitor_1__EVAL_4;
  wire [1:0] TLMonitor_1__EVAL_5;
  wire [2:0] TLMonitor_1__EVAL_6;
  wire  TLMonitor_1__EVAL_7;
  wire [11:0] TLMonitor_1__EVAL_8;
  wire [1:0] TLMonitor_1__EVAL_9;
  wire [2:0] TLMonitor_1__EVAL_10;
  wire [2:0] TLMonitor_1__EVAL_11;
  wire  TLMonitor_1__EVAL_12;
  wire  TLMonitor_1__EVAL_13;
  wire [2:0] TLMonitor_1__EVAL_14;
  wire  _EVAL_469;
  wire  _EVAL_472;
  wire  _EVAL_475;
  wire  _EVAL_476;
  wire  _EVAL_478;
  wire  _EVAL_482;
  wire  _EVAL_483;
  wire  _EVAL_489;
  wire  _EVAL_490;
  wire  _EVAL_491;
  wire  _EVAL_494;
  wire  _EVAL_495;
  wire  _EVAL_496;
  wire  _EVAL_500;
  wire  _EVAL_501;
  wire  _EVAL_503;
  wire  _EVAL_504;
  wire  _EVAL_507;
  wire  _EVAL_508;
  wire  _EVAL_511;
  wire  _EVAL_513;
  wire  _EVAL_515;
  wire  _EVAL_517;
  wire  _EVAL_518;
  wire  _EVAL_520;
  wire  _EVAL_521;
  wire  _EVAL_523;
  wire  _EVAL_524;
  wire  _EVAL_525;
  wire  _EVAL_528;
  wire  _EVAL_529;
  wire  _EVAL_531;
  wire  _EVAL_532;
  wire  _EVAL_534;
  wire  _EVAL_535;
  wire  _EVAL_536;
  wire  _EVAL_537;
  wire  _EVAL_539;
  wire  _EVAL_543;
  wire  _EVAL_544;
  wire  _EVAL_548;
  wire  _EVAL_550;
  wire  _EVAL_553;
  wire  _EVAL_556;
  wire  _EVAL_557;
  wire  _EVAL_560;
  wire  _EVAL_561;
  wire  _EVAL_562;
  wire  _EVAL_564;
  wire  _EVAL_568;
  wire  _EVAL_570;
  wire  _EVAL_573;
  wire  _EVAL_574;
  wire  _EVAL_576;
  wire  _EVAL_578;
  wire  _EVAL_579;
  wire  _EVAL_580;
  wire  _EVAL_581;
  wire  _EVAL_582;
  wire  _EVAL_584;
  wire  _EVAL_586;
  wire  _EVAL_587;
  wire  _EVAL_588;
  wire  _EVAL_589;
  wire  _EVAL_591;
  wire  _EVAL_593;
  wire  _EVAL_594;
  wire  _EVAL_595;
  wire  _EVAL_596;
  wire  _EVAL_597;
  wire  _EVAL_598;
  wire  _EVAL_600;
  wire  _EVAL_603;
  wire  _EVAL_604;
  wire  _EVAL_609;
  wire  _EVAL_610;
  wire  _EVAL_615;
  wire  _EVAL_618;
  wire  _EVAL_621;
  wire  _EVAL_623;
  wire  _EVAL_625;
  wire  _EVAL_626;
  wire  _EVAL_627;
  wire  _EVAL_629;
  wire  _EVAL_631;
  wire  _EVAL_632;
  wire  _EVAL_633;
  wire  _EVAL_635;
  wire  _EVAL_637;
  wire  _EVAL_639;
  wire  _EVAL_640;
  wire  _EVAL_641;
  wire  _EVAL_643;
  wire  _EVAL_644;
  wire  _EVAL_646;
  wire  _EVAL_647;
  wire  _EVAL_648;
  wire  _EVAL_652;
  wire  _EVAL_655;
  wire  _EVAL_656;
  wire  _EVAL_657;
  wire  _EVAL_658;
  wire  _EVAL_660;
  wire  _EVAL_661;
  wire  _EVAL_663;
  wire  _EVAL_664;
  wire  _EVAL_665;
  wire  _EVAL_666;
  wire  _EVAL_667;
  wire  _EVAL_668;
  wire  _EVAL_670;
  wire  _EVAL_671;
  wire  _EVAL_672;
  wire [3:0] _EVAL_673;
  wire  _EVAL_675;
  wire  _EVAL_676;
  wire  _EVAL_677;
  wire  _EVAL_678;
  wire  _EVAL_680;
  wire  _EVAL_681;
  wire  _EVAL_682;
  wire  _EVAL_684;
  wire  _EVAL_687;
  wire  _EVAL_688;
  wire  _EVAL_690;
  wire  _EVAL_691;
  wire  _EVAL_693;
  wire  _EVAL_694;
  wire  _EVAL_695;
  wire  _EVAL_698;
  wire  _EVAL_701;
  wire  _EVAL_703;
  wire  _EVAL_704;
  wire  _EVAL_706;
  wire  _EVAL_708;
  wire  _EVAL_709;
  wire  _EVAL_712;
  wire  _EVAL_714;
  wire  _EVAL_715;
  wire  _EVAL_716;
  wire  _EVAL_717;
  wire  _EVAL_718;
  wire  _EVAL_720;
  wire  _EVAL_726;
  wire  _EVAL_729;
  wire  _EVAL_731;
  wire  _EVAL_732;
  wire  _EVAL_733;
  wire  _EVAL_737;
  wire  _EVAL_738;
  wire  _EVAL_740;
  wire  _EVAL_741;
  wire  _EVAL_742;
  wire  _EVAL_743;
  wire  _EVAL_745;
  wire  _EVAL_746;
  wire  _EVAL_747;
  wire  _EVAL_749;
  wire  _EVAL_750;
  wire  _EVAL_755;
  wire  _EVAL_756;
  wire  _EVAL_758;
  wire  _EVAL_761;
  wire  _EVAL_764;
  wire  _EVAL_767;
  wire  _EVAL_770;
  wire  _EVAL_772;
  wire  _EVAL_773;
  wire  _EVAL_775;
  wire  _EVAL_776;
  wire  _EVAL_777;
  wire  _EVAL_778;
  wire  _EVAL_779;
  wire  _EVAL_780;
  wire  _EVAL_781;
  wire  _EVAL_782;
  wire  _EVAL_783;
  wire  _EVAL_786;
  wire  _EVAL_787;
  wire  _EVAL_791;
  wire  _EVAL_794;
  wire  _EVAL_796;
  wire  _EVAL_798;
  wire  _EVAL_800;
  wire  _EVAL_801;
  wire  _EVAL_803;
  wire  _EVAL_804;
  wire  _EVAL_805;
  wire  _EVAL_806;
  wire  _EVAL_807;
  wire  _EVAL_810;
  wire  _EVAL_811;
  wire  _EVAL_812;
  wire  _EVAL_813;
  wire  _EVAL_814;
  wire  _EVAL_816;
  wire  _EVAL_818;
  wire  _EVAL_821;
  wire  _EVAL_823;
  wire  _EVAL_824;
  wire  _EVAL_825;
  wire  _EVAL_826;
  wire  _EVAL_827;
  wire  _EVAL_828;
  wire  _EVAL_830;
  wire  _EVAL_831;
  wire  _EVAL_834;
  wire  _EVAL_838;
  wire  _EVAL_839;
  wire  _EVAL_840;
  wire  _EVAL_843;
  wire  _EVAL_844;
  wire  _EVAL_845;
  wire  _EVAL_848;
  wire  _EVAL_850;
  wire  _EVAL_852;
  wire  _EVAL_853;
  wire  _EVAL_854;
  wire  _EVAL_855;
  wire  _EVAL_856;
  wire  _EVAL_860;
  wire  _EVAL_862;
  wire  _EVAL_864;
  wire  _EVAL_865;
  wire  _EVAL_871;
  wire  _EVAL_872;
  wire  _EVAL_873;
  wire  _EVAL_874;
  wire  _EVAL_877;
  wire  _EVAL_878;
  wire  _EVAL_880;
  wire  _EVAL_883;
  wire  _EVAL_884;
  wire  _EVAL_885;
  wire  _EVAL_887;
  wire  _EVAL_888;
  wire  _EVAL_889;
  wire  _EVAL_892;
  wire  _EVAL_893;
  wire  _EVAL_894;
  wire  _EVAL_896;
  wire  _EVAL_897;
  wire  _EVAL_898;
  wire  _EVAL_899;
  wire  _EVAL_901;
  wire  _EVAL_902;
  wire  _EVAL_903;
  wire  _EVAL_904;
  wire  _EVAL_905;
  wire  _EVAL_907;
  wire  _EVAL_911;
  wire  _EVAL_913;
  wire  _EVAL_914;
  wire  _EVAL_917;
  wire  _EVAL_918;
  wire  _EVAL_919;
  wire  _EVAL_920;
  wire  _EVAL_923;
  wire  _EVAL_924;
  wire  _EVAL_925;
  wire  _EVAL_927;
  wire  _EVAL_928;
  wire  _EVAL_929;
  wire  _EVAL_932;
  wire  _EVAL_933;
  wire  _EVAL_935;
  wire  _EVAL_936;
  wire  _EVAL_937;
  wire  _EVAL_938;
  wire  _EVAL_939;
  wire  _EVAL_940;
  wire  _EVAL_944;
  wire  _EVAL_945;
  wire  _EVAL_947;
  wire  _EVAL_948;
  wire  _EVAL_950;
  wire  _EVAL_953;
  wire  _EVAL_954;
  wire  _EVAL_955;
  wire  _EVAL_961;
  wire  _EVAL_962;
  wire  _EVAL_966;
  wire  _EVAL_970;
  wire  _EVAL_971;
  wire  _EVAL_973;
  wire  _EVAL_974;
  wire  _EVAL_975;
  wire  _EVAL_976;
  wire  _EVAL_977;
  wire  _EVAL_978;
  wire  _EVAL_979;
  wire  _EVAL_980;
  wire  _EVAL_981;
  wire  _EVAL_983;
  wire  _EVAL_986;
  wire  _EVAL_988;
  wire  _EVAL_989;
  wire  _EVAL_992;
  wire  _EVAL_994;
  wire  _EVAL_998;
  wire  _EVAL_999;
  wire  _EVAL_1001;
  wire  _EVAL_1002;
  wire  _EVAL_1005;
  wire  _EVAL_1006;
  wire  _EVAL_1009;
  wire  _EVAL_1011;
  wire  _EVAL_1013;
  wire  _EVAL_1016;
  wire  _EVAL_1017;
  wire  _EVAL_1022;
  wire  _EVAL_1024;
  wire  _EVAL_1025;
  wire  _EVAL_1028;
  wire  _EVAL_1029;
  wire  _EVAL_1032;
  wire  _EVAL_1033;
  wire  _EVAL_1042;
  wire  _EVAL_1043;
  wire  _EVAL_1048;
  wire  _EVAL_1053;
  wire  _EVAL_1054;
  wire  _EVAL_1055;
  wire  _EVAL_1056;
  wire  _EVAL_1058;
  wire  _EVAL_1059;
  wire  _EVAL_1060;
  wire [14:0] _EVAL_1061;
  wire  _EVAL_1062;
  wire  _EVAL_1063;
  wire  _EVAL_1064;
  wire  _EVAL_1065;
  wire  _EVAL_1067;
  wire  _EVAL_1068;
  wire  _EVAL_1070;
  wire  _EVAL_1072;
  wire  _EVAL_1074;
  wire  _EVAL_1075;
  wire  _EVAL_1076;
  wire  _EVAL_1078;
  wire  _EVAL_1079;
  wire  _EVAL_1080;
  wire  _EVAL_1083;
  wire  _EVAL_1085;
  wire  _EVAL_1088;
  wire  _EVAL_1090;
  wire  _EVAL_1091;
  wire  _EVAL_1092;
  wire  _EVAL_1093;
  wire  _EVAL_1094;
  wire  _EVAL_1100;
  wire  _EVAL_1102;
  wire  _EVAL_1103;
  wire  _EVAL_1105;
  wire  _EVAL_1106;
  wire  _EVAL_1107;
  wire  _EVAL_1108;
  wire  _EVAL_1111;
  wire  _EVAL_1112;
  wire  _EVAL_1113;
  wire  _EVAL_1117;
  wire  _EVAL_1118;
  wire  _EVAL_1119;
  wire  _EVAL_1120;
  wire  _EVAL_1122;
  wire  _EVAL_1126;
  wire  _EVAL_1128;
  wire  _EVAL_1129;
  wire  _EVAL_1130;
  wire  _EVAL_1134;
  wire  _EVAL_1137;
  wire  _EVAL_1141;
  wire  _EVAL_1142;
  wire  _EVAL_1143;
  wire  _EVAL_1144;
  wire  _EVAL_1146;
  wire  _EVAL_1148;
  wire  _EVAL_1153;
  wire  _EVAL_1156;
  wire  _EVAL_1157;
  wire  _EVAL_1158;
  wire  _EVAL_1161;
  wire  _EVAL_1162;
  wire  _EVAL_1164;
  wire  _EVAL_1165;
  wire  _EVAL_1168;
  wire  _EVAL_1169;
  wire  _EVAL_1171;
  wire  _EVAL_1172;
  wire  _EVAL_1173;
  wire  _EVAL_1178;
  wire  _EVAL_1179;
  wire  _EVAL_1187;
  wire  _EVAL_1188;
  wire  _EVAL_1189;
  wire  _EVAL_1190;
  wire  _EVAL_1192;
  wire  _EVAL_1193;
  wire  _EVAL_1195;
  wire  _EVAL_1197;
  wire  _EVAL_1199;
  wire  _EVAL_1201;
  wire  _EVAL_1202;
  wire  _EVAL_1203;
  wire  _EVAL_1204;
  wire  _EVAL_1205;
  wire  _EVAL_1207;
  wire  _EVAL_1208;
  wire [1:0] _EVAL_1209;
  wire  _EVAL_1210;
  wire  _EVAL_1212;
  wire  _EVAL_1214;
  wire  _EVAL_1216;
  wire  _EVAL_1222;
  wire  _EVAL_1223;
  wire  _EVAL_1225;
  wire  _EVAL_1227;
  wire  _EVAL_1229;
  wire  _EVAL_1232;
  wire  _EVAL_1233;
  wire  _EVAL_1234;
  wire  _EVAL_1235;
  wire  _EVAL_1236;
  wire  _EVAL_1239;
  wire  _EVAL_1241;
  wire  _EVAL_1242;
  wire  _EVAL_1245;
  wire  _EVAL_1246;
  wire  _EVAL_1247;
  wire  _EVAL_1248;
  wire  _EVAL_1249;
  wire  _EVAL_1250;
  wire  _EVAL_1252;
  wire  _EVAL_1253;
  wire  _EVAL_1254;
  wire  _EVAL_1255;
  wire  _EVAL_1256;
  wire  _EVAL_1259;
  wire  _EVAL_1260;
  wire  _EVAL_1262;
  wire  _EVAL_1263;
  wire  _EVAL_1264;
  wire  _EVAL_1265;
  wire  _EVAL_1266;
  wire  _EVAL_1267;
  wire  _EVAL_1272;
  wire  _EVAL_1277;
  wire  _EVAL_1278;
  wire  _EVAL_1279;
  wire  _EVAL_1280;
  wire  _EVAL_1281;
  wire  _EVAL_1282;
  wire  _EVAL_1283;
  wire  _EVAL_1284;
  wire  _EVAL_1286;
  wire  _EVAL_1287;
  wire  _EVAL_1288;
  wire  _EVAL_1289;
  wire  _EVAL_1291;
  wire  _EVAL_1292;
  wire  _EVAL_1293;
  wire  _EVAL_1294;
  wire  _EVAL_1295;
  wire  _EVAL_1296;
  wire  _EVAL_1298;
  wire  _EVAL_1299;
  wire  _EVAL_1300;
  wire  _EVAL_1301;
  wire  _EVAL_1302;
  wire  _EVAL_1305;
  wire  _EVAL_1306;
  wire  _EVAL_1308;
  wire  _EVAL_1309;
  wire  _EVAL_1310;
  wire  _EVAL_1313;
  wire  _EVAL_1315;
  wire  _EVAL_1316;
  wire  _EVAL_1317;
  wire  _EVAL_1318;
  wire  _EVAL_1320;
  wire  _EVAL_1322;
  wire  _EVAL_1323;
  wire  _EVAL_1327;
  wire  _EVAL_1329;
  wire  _EVAL_1330;
  wire  _EVAL_1333;
  wire  _EVAL_1336;
  wire  _EVAL_1338;
  wire  _EVAL_1340;
  wire  _EVAL_1342;
  wire  _EVAL_1344;
  wire  _EVAL_1345;
  wire  _EVAL_1346;
  wire  _EVAL_1349;
  wire  _EVAL_1352;
  wire  _EVAL_1353;
  wire  _EVAL_1354;
  wire  _EVAL_1355;
  wire  _EVAL_1356;
  wire  _EVAL_1359;
  wire  _EVAL_1361;
  wire  _EVAL_1363;
  wire  _EVAL_1364;
  wire  _EVAL_1369;
  wire  _EVAL_1371;
  wire  _EVAL_1372;
  wire  _EVAL_1373;
  wire  _EVAL_1378;
  wire  _EVAL_1379;
  wire  _EVAL_1381;
  wire  _EVAL_1382;
  wire  _EVAL_1384;
  wire  _EVAL_1385;
  wire  _EVAL_1386;
  wire  _EVAL_1387;
  wire  _EVAL_1388;
  wire  _EVAL_1389;
  wire  _EVAL_1391;
  wire  _EVAL_1393;
  wire  _EVAL_1394;
  wire  _EVAL_1396;
  wire  _EVAL_1397;
  wire  _EVAL_1398;
  wire  _EVAL_1402;
  wire  _EVAL_1404;
  wire  _EVAL_1405;
  wire  _EVAL_1406;
  wire  _EVAL_1409;
  wire  _EVAL_1411;
  wire  _EVAL_1412;
  wire  _EVAL_1413;
  wire  _EVAL_1414;
  wire  _EVAL_1415;
  wire  _EVAL_1416;
  wire  _EVAL_1417;
  wire  _EVAL_1421;
  wire  _EVAL_1424;
  wire  _EVAL_1427;
  wire  _EVAL_1428;
  wire  _EVAL_1430;
  wire  _EVAL_1431;
  wire  _EVAL_1432;
  wire  _EVAL_1434;
  wire  _EVAL_1438;
  wire  _EVAL_1439;
  wire  _EVAL_1440;
  wire  _EVAL_1442;
  wire  _EVAL_1443;
  wire  _EVAL_1444;
  wire  _EVAL_1446;
  wire  _EVAL_1447;
  wire  _EVAL_1449;
  wire  _EVAL_1451;
  wire  _EVAL_1452;
  wire  _EVAL_1453;
  wire  _EVAL_1454;
  wire  _EVAL_1455;
  wire  _EVAL_1456;
  wire  _EVAL_1457;
  wire  _EVAL_1458;
  wire  _EVAL_1459;
  wire  _EVAL_1463;
  wire  _EVAL_1464;
  wire  _EVAL_1466;
  wire  _EVAL_1473;
  wire  _EVAL_1479;
  wire  _EVAL_1481;
  wire  _EVAL_1482;
  wire  _EVAL_1483;
  wire  _EVAL_1484;
  wire  _EVAL_1485;
  wire  _EVAL_1489;
  wire  _EVAL_1491;
  wire  _EVAL_1492;
  wire  _EVAL_1497;
  wire  _EVAL_1498;
  wire  _EVAL_1499;
  wire  _EVAL_1500;
  wire  _EVAL_1501;
  wire  _EVAL_1502;
  wire  _EVAL_1503;
  wire  _EVAL_1504;
  wire  _EVAL_1505;
  wire  _EVAL_1509;
  wire  _EVAL_1510;
  wire  _EVAL_1511;
  wire  _EVAL_1515;
  wire  _EVAL_1519;
  wire  _EVAL_1520;
  wire  _EVAL_1521;
  wire  _EVAL_1522;
  wire  _EVAL_1524;
  wire  _EVAL_1526;
  wire  _EVAL_1529;
  wire  _EVAL_1531;
  wire  _EVAL_1533;
  wire  _EVAL_1534;
  wire  _EVAL_1535;
  wire  _EVAL_1536;
  wire  _EVAL_1537;
  wire  _EVAL_1539;
  wire  _EVAL_1542;
  wire  _EVAL_1543;
  wire  _EVAL_1548;
  wire  _EVAL_1550;
  wire  _EVAL_1551;
  wire  _EVAL_1554;
  wire  _EVAL_1555;
  wire  _EVAL_1558;
  wire  _EVAL_1559;
  wire  _EVAL_1560;
  wire  _EVAL_1563;
  wire  _EVAL_1565;
  wire  _EVAL_1566;
  wire  _EVAL_1570;
  wire  _EVAL_1573;
  wire  _EVAL_1574;
  wire  _EVAL_1577;
  wire  _EVAL_1579;
  wire  _EVAL_1580;
  wire  _EVAL_1581;
  wire  _EVAL_1582;
  wire  _EVAL_1584;
  wire  _EVAL_1585;
  wire  _EVAL_1586;
  wire  _EVAL_1588;
  wire  _EVAL_1595;
  wire  _EVAL_1596;
  wire  _EVAL_1600;
  wire  _EVAL_1601;
  wire  _EVAL_1602;
  wire  _EVAL_1604;
  wire  _EVAL_1605;
  wire  _EVAL_1607;
  wire  _EVAL_1608;
  wire  _EVAL_1609;
  wire  _EVAL_1610;
  wire  _EVAL_1612;
  wire  _EVAL_1614;
  wire  _EVAL_1616;
  wire  _EVAL_1617;
  wire  _EVAL_1618;
  wire  _EVAL_1619;
  wire  _EVAL_1621;
  wire  _EVAL_1623;
  wire  _EVAL_1624;
  wire  _EVAL_1625;
  wire  _EVAL_1626;
  wire  _EVAL_1627;
  wire  _EVAL_1628;
  wire  _EVAL_1629;
  wire  _EVAL_1630;
  wire  _EVAL_1632;
  wire  _EVAL_1634;
  wire  _EVAL_1635;
  wire  _EVAL_1636;
  wire  _EVAL_1637;
  wire  _EVAL_1638;
  wire  _EVAL_1640;
  wire  _EVAL_1642;
  wire  _EVAL_1643;
  wire  _EVAL_1644;
  wire  _EVAL_1645;
  wire  _EVAL_1647;
  wire  _EVAL_1648;
  wire  _EVAL_1649;
  wire  _EVAL_1651;
  wire  _EVAL_1652;
  wire  _EVAL_1655;
  wire  _EVAL_1656;
  wire  _EVAL_1657;
  wire  _EVAL_1660;
  wire  _EVAL_1661;
  wire  _EVAL_1662;
  wire  _EVAL_1663;
  wire  _EVAL_1664;
  wire  _EVAL_1667;
  wire  _EVAL_1668;
  wire  _EVAL_1670;
  wire  _EVAL_1671;
  wire  _EVAL_1673;
  wire  _EVAL_1674;
  wire  _EVAL_1676;
  wire  _EVAL_1679;
  wire  _EVAL_1680;
  wire  _EVAL_1683;
  wire  _EVAL_1686;
  wire  _EVAL_1688;
  wire  _EVAL_1689;
  wire  _EVAL_1690;
  wire  _EVAL_1691;
  wire  _EVAL_1692;
  wire  _EVAL_1695;
  wire  _EVAL_1696;
  wire  _EVAL_1698;
  wire  _EVAL_1700;
  wire  _EVAL_1702;
  wire  _EVAL_1703;
  wire  _EVAL_1704;
  wire  _EVAL_1705;
  wire  _EVAL_1707;
  wire  _EVAL_1708;
  wire  _EVAL_1709;
  wire  _EVAL_1711;
  wire  _EVAL_1712;
  wire  _EVAL_1714;
  wire  _EVAL_1715;
  wire  _EVAL_1716;
  wire  _EVAL_1717;
  wire  _EVAL_1719;
  wire  _EVAL_1722;
  wire  _EVAL_1726;
  wire  _EVAL_1727;
  wire  _EVAL_1729;
  wire  _EVAL_1730;
  wire  _EVAL_1733;
  wire  _EVAL_1735;
  wire  _EVAL_1737;
  wire  _EVAL_1739;
  wire  _EVAL_1740;
  wire  _EVAL_1741;
  wire  _EVAL_1743;
  wire  _EVAL_1744;
  wire  _EVAL_1745;
  wire  _EVAL_1748;
  wire  _EVAL_1749;
  wire  _EVAL_1750;
  wire  _EVAL_1751;
  wire  _EVAL_1753;
  wire  _EVAL_1756;
  wire  _EVAL_1757;
  wire  _EVAL_1760;
  wire  _EVAL_1762;
  wire  _EVAL_1763;
  wire  _EVAL_1764;
  wire  _EVAL_1765;
  wire  _EVAL_1766;
  wire  _EVAL_1768;
  wire  _EVAL_1770;
  wire  _EVAL_1772;
  wire  _EVAL_1775;
  wire  _EVAL_1776;
  wire  _EVAL_1777;
  wire  _EVAL_1780;
  wire  _EVAL_1781;
  wire  _EVAL_1782;
  wire  _EVAL_1783;
  wire  _EVAL_1784;
  wire  _EVAL_1785;
  wire  _EVAL_1786;
  wire  _EVAL_1788;
  wire  _EVAL_1791;
  wire  _EVAL_1792;
  wire  _EVAL_1793;
  wire  _EVAL_1794;
  wire  _EVAL_1796;
  wire  _EVAL_1797;
  wire  _EVAL_1800;
  wire  _EVAL_1801;
  wire  _EVAL_1802;
  wire  _EVAL_1808;
  wire  _EVAL_1809;
  wire  _EVAL_1810;
  wire  _EVAL_1811;
  wire  _EVAL_1814;
  wire  _EVAL_1816;
  wire  _EVAL_1817;
  wire  _EVAL_1818;
  wire  _EVAL_1819;
  wire  _EVAL_1820;
  wire  _EVAL_1825;
  wire  _EVAL_1826;
  wire  _EVAL_1827;
  wire  _EVAL_1828;
  wire  _EVAL_1829;
  wire  _EVAL_1831;
  wire  _EVAL_1836;
  wire  _EVAL_1837;
  wire  _EVAL_1840;
  wire  _EVAL_1843;
  wire  _EVAL_1847;
  wire  _EVAL_1848;
  wire  _EVAL_1850;
  wire  _EVAL_1851;
  wire  _EVAL_1852;
  wire  _EVAL_1854;
  wire  _EVAL_1855;
  wire  _EVAL_1857;
  wire  _EVAL_1858;
  wire  _EVAL_1861;
  wire  _EVAL_1862;
  wire  _EVAL_1864;
  wire  _EVAL_1865;
  wire  _EVAL_1866;
  wire  _EVAL_1868;
  wire  _EVAL_1870;
  wire  _EVAL_1874;
  wire  _EVAL_1876;
  wire  _EVAL_1877;
  wire  _EVAL_1879;
  wire  _EVAL_1882;
  wire  _EVAL_1885;
  wire  _EVAL_1886;
  wire  _EVAL_1889;
  wire  _EVAL_1890;
  wire  _EVAL_1892;
  wire  _EVAL_1895;
  wire  _EVAL_1898;
  wire  _EVAL_1899;
  wire  _EVAL_1901;
  wire  _EVAL_1903;
  wire  _EVAL_1904;
  wire  _EVAL_1906;
  wire  _EVAL_1907;
  wire  _EVAL_1908;
  wire  _EVAL_1909;
  wire  _EVAL_1910;
  wire  _EVAL_1912;
  wire  _EVAL_1915;
  wire  _EVAL_1916;
  wire  _EVAL_1917;
  wire  _EVAL_1918;
  wire  _EVAL_1919;
  wire  _EVAL_1920;
  wire  _EVAL_1922;
  wire  _EVAL_1923;
  wire  _EVAL_1924;
  wire  _EVAL_1926;
  wire  _EVAL_1927;
  wire  _EVAL_1929;
  wire  _EVAL_1930;
  wire  _EVAL_1932;
  wire  _EVAL_1938;
  wire  _EVAL_1940;
  wire  _EVAL_1943;
  wire  _EVAL_1946;
  wire  _EVAL_1947;
  wire  _EVAL_1948;
  wire  _EVAL_1949;
  wire  _EVAL_1950;
  wire  _EVAL_1951;
  wire  _EVAL_1952;
  wire  _EVAL_1954;
  wire  _EVAL_1955;
  wire  _EVAL_1956;
  wire  _EVAL_1960;
  wire  _EVAL_1961;
  wire  _EVAL_1962;
  wire  _EVAL_1963;
  wire  _EVAL_1964;
  wire  _EVAL_1966;
  wire  _EVAL_1967;
  wire  _EVAL_1969;
  wire  _EVAL_1970;
  wire [3:0] _EVAL_1971;
  wire  _EVAL_1973;
  wire  _EVAL_1974;
  wire  _EVAL_1976;
  wire  _EVAL_1980;
  wire  _EVAL_1981;
  wire  _EVAL_1984;
  wire  _EVAL_1986;
  wire  _EVAL_1988;
  wire  _EVAL_1990;
  wire  _EVAL_1995;
  wire  _EVAL_1996;
  wire  _EVAL_1997;
  wire  _EVAL_1998;
  wire  _EVAL_1999;
  wire  _EVAL_2000;
  wire  _EVAL_2003;
  wire  _EVAL_2007;
  wire  _EVAL_2009;
  wire  _EVAL_2010;
  wire  _EVAL_2011;
  wire  _EVAL_2013;
  wire  _EVAL_2016;
  wire  _EVAL_2019;
  wire  _EVAL_2020;
  wire  _EVAL_2022;
  wire  _EVAL_2023;
  wire  _EVAL_2025;
  wire  _EVAL_2026;
  wire  _EVAL_2027;
  wire  _EVAL_2028;
  wire  _EVAL_2030;
  wire  _EVAL_2032;
  wire  _EVAL_2033;
  wire  _EVAL_2034;
  wire  _EVAL_2036;
  wire  _EVAL_2037;
  wire  _EVAL_2038;
  wire  _EVAL_2042;
  wire  _EVAL_2043;
  wire  _EVAL_2044;
  wire  _EVAL_2045;
  wire  _EVAL_2046;
  wire  _EVAL_2047;
  wire  _EVAL_2048;
  wire  _EVAL_2049;
  wire  _EVAL_2053;
  wire  _EVAL_2055;
  wire  _EVAL_2058;
  wire  _EVAL_2059;
  wire  _EVAL_2060;
  wire  _EVAL_2062;
  wire  _EVAL_2064;
  wire  _EVAL_2065;
  wire  _EVAL_2067;
  wire  _EVAL_2068;
  wire  _EVAL_2069;
  wire  _EVAL_2070;
  wire  _EVAL_2071;
  wire  _EVAL_2072;
  wire  _EVAL_2082;
  wire  _EVAL_2084;
  wire  _EVAL_2085;
  wire  _EVAL_2087;
  wire  _EVAL_2088;
  wire  _EVAL_2093;
  wire  _EVAL_2094;
  wire  _EVAL_2098;
  wire  _EVAL_2099;
  wire  _EVAL_2100;
  wire  _EVAL_2105;
  wire  _EVAL_2107;
  wire  _EVAL_2108;
  wire  _EVAL_2109;
  wire  _EVAL_2112;
  wire  _EVAL_2114;
  wire  _EVAL_2117;
  wire  _EVAL_2118;
  wire  _EVAL_2119;
  wire  _EVAL_2122;
  wire  _EVAL_2123;
  wire  _EVAL_2124;
  wire  _EVAL_2126;
  wire  _EVAL_2127;
  wire  _EVAL_2129;
  wire  _EVAL_2131;
  wire  _EVAL_2132;
  wire  _EVAL_2133;
  wire  _EVAL_2134;
  wire  _EVAL_2135;
  wire  _EVAL_2137;
  wire  _EVAL_2139;
  wire  _EVAL_2140;
  wire  _EVAL_2141;
  wire  _EVAL_2142;
  wire  _EVAL_2146;
  wire  _EVAL_2147;
  wire  _EVAL_2148;
  wire  _EVAL_2150;
  wire  _EVAL_2151;
  wire  _EVAL_2152;
  wire  _EVAL_2153;
  wire  _EVAL_2154;
  wire  _EVAL_2155;
  wire  _EVAL_2158;
  wire  _EVAL_2159;
  wire  _EVAL_2161;
  wire  _EVAL_2164;
  wire  _EVAL_2165;
  wire  _EVAL_2167;
  wire  _EVAL_2169;
  wire  _EVAL_2170;
  wire  _EVAL_2171;
  wire  _EVAL_2172;
  wire  _EVAL_2176;
  wire  _EVAL_2179;
  wire  _EVAL_2180;
  wire  _EVAL_2181;
  wire  _EVAL_2182;
  wire  _EVAL_2184;
  wire  _EVAL_2186;
  wire  _EVAL_2187;
  wire  _EVAL_2189;
  wire  _EVAL_2191;
  wire  _EVAL_2192;
  wire  _EVAL_2195;
  wire  _EVAL_2197;
  wire  _EVAL_2198;
  wire  _EVAL_2199;
  wire  _EVAL_2200;
  wire  _EVAL_2201;
  wire  _EVAL_2202;
  wire  _EVAL_2203;
  wire  _EVAL_2204;
  wire  _EVAL_2205;
  wire  _EVAL_2206;
  wire  _EVAL_2208;
  wire  _EVAL_2209;
  wire  _EVAL_2212;
  wire  _EVAL_2213;
  wire  _EVAL_2214;
  wire  _EVAL_2221;
  wire  _EVAL_2225;
  wire  _EVAL_2226;
  wire  _EVAL_2227;
  wire  _EVAL_2228;
  wire  _EVAL_2229;
  wire  _EVAL_2230;
  wire  _EVAL_2231;
  wire  _EVAL_2232;
  wire  _EVAL_2234;
  wire  _EVAL_2236;
  wire  _EVAL_2239;
  wire  _EVAL_2240;
  wire  _EVAL_2241;
  wire  _EVAL_2242;
  wire  _EVAL_2243;
  wire  _EVAL_2244;
  wire  _EVAL_2245;
  wire  _EVAL_2250;
  wire  _EVAL_2252;
  wire  _EVAL_2253;
  wire  _EVAL_2257;
  wire  _EVAL_2258;
  wire  _EVAL_2259;
  wire  _EVAL_2260;
  wire  _EVAL_2263;
  wire  _EVAL_2266;
  wire [4:0] _EVAL_2267;
  wire  _EVAL_2269;
  wire  _EVAL_2270;
  wire  _EVAL_2271;
  wire  _EVAL_2273;
  wire  _EVAL_2276;
  wire  _EVAL_2278;
  wire  _EVAL_2281;
  wire  _EVAL_2282;
  wire  _EVAL_2283;
  wire  _EVAL_2287;
  wire  _EVAL_2288;
  wire  _EVAL_2289;
  wire  _EVAL_2292;
  wire  _EVAL_2293;
  wire  _EVAL_2296;
  wire  _EVAL_2297;
  wire  _EVAL_2300;
  wire  _EVAL_2301;
  wire  _EVAL_2303;
  wire  _EVAL_2304;
  wire  _EVAL_2305;
  wire  _EVAL_2307;
  wire  _EVAL_2309;
  wire  _EVAL_2310;
  wire  _EVAL_2313;
  wire  _EVAL_2315;
  wire  _EVAL_2316;
  wire  _EVAL_2319;
  wire  _EVAL_2320;
  wire  _EVAL_2321;
  wire  _EVAL_2322;
  wire  _EVAL_2323;
  wire  _EVAL_2327;
  wire  _EVAL_2329;
  wire  _EVAL_2330;
  wire  _EVAL_2331;
  wire  _EVAL_2335;
  wire  _EVAL_2337;
  wire  _EVAL_2338;
  wire  _EVAL_2341;
  wire  _EVAL_2342;
  wire  _EVAL_2345;
  wire  _EVAL_2346;
  wire  _EVAL_2348;
  wire  _EVAL_2349;
  wire  _EVAL_2350;
  wire  _EVAL_2352;
  wire  _EVAL_2353;
  wire  _EVAL_2355;
  wire  _EVAL_2356;
  wire  _EVAL_2357;
  wire  _EVAL_2361;
  wire  _EVAL_2362;
  wire  _EVAL_2364;
  wire  _EVAL_2369;
  wire  _EVAL_2370;
  wire  _EVAL_2372;
  wire  _EVAL_2374;
  wire  _EVAL_2375;
  wire  _EVAL_2376;
  wire  _EVAL_2377;
  wire  _EVAL_2380;
  wire  _EVAL_2381;
  wire  _EVAL_2382;
  wire  _EVAL_2386;
  wire  _EVAL_2388;
  wire  _EVAL_2389;
  wire  _EVAL_2391;
  wire  _EVAL_2393;
  wire  _EVAL_2394;
  wire  _EVAL_2396;
  wire  _EVAL_2397;
  wire  _EVAL_2401;
  wire [11:0] _EVAL_2404;
  wire  _EVAL_2405;
  wire  _EVAL_2406;
  wire  _EVAL_2407;
  wire  _EVAL_2408;
  wire  _EVAL_2409;
  wire  _EVAL_2413;
  wire  _EVAL_2415;
  wire  _EVAL_2416;
  wire  _EVAL_2421;
  wire  _EVAL_2423;
  wire  _EVAL_2424;
  wire  _EVAL_2425;
  wire  _EVAL_2426;
  wire  _EVAL_2427;
  wire  _EVAL_2428;
  wire  _EVAL_2430;
  wire  _EVAL_2431;
  wire  _EVAL_2433;
  wire  _EVAL_2434;
  wire  _EVAL_2435;
  wire  _EVAL_2436;
  wire  _EVAL_2439;
  wire  _EVAL_2441;
  wire  _EVAL_2442;
  wire  _EVAL_2443;
  wire  _EVAL_2444;
  wire  _EVAL_2446;
  wire  _EVAL_2448;
  wire  _EVAL_2449;
  wire  _EVAL_2450;
  wire  _EVAL_2454;
  wire  _EVAL_2460;
  wire  _EVAL_2461;
  wire  _EVAL_2462;
  wire  _EVAL_2465;
  wire  _EVAL_2466;
  wire  _EVAL_2467;
  wire  _EVAL_2468;
  wire  _EVAL_2469;
  wire  _EVAL_2470;
  wire  _EVAL_2473;
  wire  _EVAL_2474;
  wire  _EVAL_2475;
  wire  _EVAL_2477;
  wire  _EVAL_2478;
  wire  _EVAL_2483;
  wire  _EVAL_2490;
  wire  _EVAL_2492;
  wire  _EVAL_2493;
  wire  _EVAL_2498;
  wire  _EVAL_2500;
  wire  _EVAL_2502;
  wire  _EVAL_2505;
  wire  _EVAL_2507;
  wire  _EVAL_2509;
  wire  _EVAL_2510;
  wire  _EVAL_2511;
  wire  _EVAL_2513;
  wire  _EVAL_2514;
  wire  _EVAL_2515;
  wire  _EVAL_2516;
  wire  _EVAL_2518;
  wire  _EVAL_2521;
  wire  _EVAL_2523;
  wire  _EVAL_2525;
  wire  _EVAL_2526;
  wire  _EVAL_2528;
  wire  _EVAL_2529;
  wire  _EVAL_2530;
  wire  _EVAL_2531;
  wire  _EVAL_2534;
  wire  _EVAL_2535;
  wire  _EVAL_2536;
  wire  _EVAL_2537;
  wire  _EVAL_2539;
  wire  _EVAL_2541;
  wire  _EVAL_2542;
  wire  _EVAL_2543;
  wire  _EVAL_2545;
  wire  _EVAL_2546;
  wire  _EVAL_2548;
  wire  _EVAL_2549;
  wire  _EVAL_2550;
  wire  _EVAL_2551;
  wire  _EVAL_2553;
  wire  _EVAL_2554;
  wire  _EVAL_2555;
  wire  _EVAL_2556;
  wire  _EVAL_2557;
  wire  _EVAL_2559;
  wire  _EVAL_2561;
  wire  _EVAL_2562;
  wire  _EVAL_2563;
  wire  _EVAL_2564;
  wire  _EVAL_2567;
  wire  _EVAL_2568;
  wire  _EVAL_2572;
  wire  _EVAL_2574;
  wire  _EVAL_2575;
  wire  _EVAL_2576;
  wire  _EVAL_2577;
  wire  _EVAL_2579;
  wire  _EVAL_2580;
  wire  _EVAL_2582;
  wire  _EVAL_2585;
  wire  _EVAL_2586;
  wire  _EVAL_2587;
  wire  _EVAL_2592;
  wire  _EVAL_2596;
  wire  _EVAL_2597;
  wire  _EVAL_2599;
  wire  _EVAL_2600;
  wire  _EVAL_2601;
  wire  _EVAL_2603;
  wire  _EVAL_2605;
  wire  _EVAL_2606;
  wire  _EVAL_2607;
  wire  _EVAL_2608;
  wire  _EVAL_2609;
  wire  _EVAL_2612;
  wire  _EVAL_2613;
  wire  _EVAL_2614;
  wire  _EVAL_2617;
  wire  _EVAL_2618;
  wire  _EVAL_2620;
  wire [1:0] TLMonitor__EVAL;
  wire  TLMonitor__EVAL_0;
  wire  TLMonitor__EVAL_1;
  wire  TLMonitor__EVAL_2;
  wire  TLMonitor__EVAL_3;
  wire  TLMonitor__EVAL_4;
  wire [1:0] TLMonitor__EVAL_5;
  wire [2:0] TLMonitor__EVAL_6;
  wire [3:0] TLMonitor__EVAL_7;
  wire  TLMonitor__EVAL_8;
  wire  TLMonitor__EVAL_9;
  wire  TLMonitor__EVAL_10;
  wire [2:0] TLMonitor__EVAL_11;
  wire [2:0] TLMonitor__EVAL_12;
  wire  TLMonitor__EVAL_13;
  wire [8:0] TLMonitor__EVAL_14;
  wire  _EVAL_2621;
  wire  _EVAL_2622;
  wire  _EVAL_2625;
  wire  _EVAL_2626;
  wire  _EVAL_2630;
  wire  _EVAL_2632;
  wire  _EVAL_2633;
  wire  _EVAL_2634;
  wire  _EVAL_2637;
  wire  _EVAL_2638;
  wire  _EVAL_2639;
  wire  _EVAL_2640;
  wire  _EVAL_2644;
  wire  _EVAL_2645;
  wire  _EVAL_2646;
  wire  _EVAL_2647;
  wire  _EVAL_2649;
  wire  _EVAL_2652;
  wire  _EVAL_2654;
  wire  _EVAL_2656;
  wire  _EVAL_2657;
  wire  _EVAL_2658;
  wire  _EVAL_2660;
  wire  _EVAL_2661;
  wire  _EVAL_2663;
  wire  _EVAL_2664;
  wire  _EVAL_2665;
  wire  _EVAL_2666;
  wire  _EVAL_2667;
  wire  _EVAL_2669;
  wire  _EVAL_2670;
  wire  _EVAL_2671;
  wire  _EVAL_2672;
  wire  _EVAL_2675;
  wire  _EVAL_2677;
  wire  _EVAL_2678;
  wire  _EVAL_2679;
  wire  _EVAL_2680;
  wire  _EVAL_2681;
  wire  _EVAL_2685;
  wire  _EVAL_2690;
  wire  _EVAL_2692;
  wire  _EVAL_2693;
  wire  _EVAL_2694;
  wire  _EVAL_2696;
  wire  _EVAL_2701;
  wire  _EVAL_2702;
  wire  _EVAL_2708;
  wire  _EVAL_2710;
  wire  _EVAL_2715;
  wire  _EVAL_2717;
  wire  _EVAL_2718;
  wire  _EVAL_2719;
  wire  _EVAL_2722;
  wire  _EVAL_2723;
  wire  _EVAL_2726;
  wire  _EVAL_2728;
  wire  _EVAL_2729;
  wire  _EVAL_2733;
  wire  _EVAL_2734;
  wire  _EVAL_2738;
  wire  _EVAL_2739;
  wire  _EVAL_2740;
  wire  _EVAL_2745;
  wire  _EVAL_2747;
  wire  _EVAL_2748;
  wire  _EVAL_2751;
  wire  _EVAL_2752;
  wire  _EVAL_2753;
  wire  _EVAL_2754;
  wire  _EVAL_2760;
  wire  _EVAL_2762;
  wire  _EVAL_2764;
  wire  _EVAL_2765;
  wire  _EVAL_2766;
  wire  _EVAL_2767;
  wire  _EVAL_2768;
  wire  _EVAL_2772;
  wire  _EVAL_2773;
  wire  _EVAL_2776;
  wire  _EVAL_2778;
  wire  _EVAL_2779;
  wire  _EVAL_2782;
  wire  _EVAL_2783;
  wire  _EVAL_2784;
  wire  _EVAL_2785;
  wire  _EVAL_2787;
  wire  _EVAL_2790;
  wire  _EVAL_2792;
  wire  _EVAL_2793;
  wire  _EVAL_2795;
  wire  _EVAL_2796;
  wire  _EVAL_2798;
  wire  _EVAL_2799;
  wire  _EVAL_2800;
  wire  _EVAL_2802;
  wire  _EVAL_2803;
  wire  _EVAL_2805;
  wire  _EVAL_2806;
  wire  _EVAL_2808;
  wire  _EVAL_2813;
  wire  _EVAL_2814;
  wire  _EVAL_2817;
  wire  _EVAL_2824;
  wire  _EVAL_2825;
  wire  _EVAL_2826;
  wire  _EVAL_2827;
  wire  _EVAL_2830;
  wire  _EVAL_2832;
  wire  _EVAL_2833;
  wire  _EVAL_2834;
  wire  _EVAL_2835;
  wire  _EVAL_2839;
  wire  _EVAL_2844;
  wire  _EVAL_2846;
  wire  _EVAL_2848;
  wire  _EVAL_2849;
  wire  _EVAL_2852;
  wire  _EVAL_2856;
  wire  _EVAL_2857;
  wire  _EVAL_2859;
  wire  _EVAL_2860;
  wire  _EVAL_2863;
  wire  _EVAL_2865;
  wire  _EVAL_2866;
  wire  _EVAL_2867;
  wire  _EVAL_2868;
  wire  _EVAL_2869;
  wire  _EVAL_2872;
  wire  _EVAL_2873;
  wire  _EVAL_2875;
  wire  _EVAL_2876;
  wire  _EVAL_2877;
  wire  _EVAL_2880;
  wire  _EVAL_2884;
  wire  _EVAL_2889;
  wire  _EVAL_2891;
  wire  _EVAL_2892;
  wire  _EVAL_2897;
  wire  _EVAL_2898;
  wire  _EVAL_2900;
  wire  _EVAL_2901;
  wire  _EVAL_2902;
  wire  _EVAL_2903;
  wire  _EVAL_2904;
  wire  _EVAL_2906;
  wire  _EVAL_2907;
  wire  _EVAL_2909;
  wire  _EVAL_2910;
  wire  _EVAL_2912;
  wire  _EVAL_2914;
  wire  _EVAL_2916;
  wire  _EVAL_2917;
  wire  _EVAL_2918;
  wire  _EVAL_2919;
  wire  _EVAL_2922;
  wire  _EVAL_2923;
  wire  _EVAL_2924;
  wire  _EVAL_2925;
  wire  _EVAL_2926;
  wire  _EVAL_2930;
  wire  _EVAL_2931;
  wire  _EVAL_2933;
  wire  _EVAL_2935;
  wire  _EVAL_2936;
  wire  _EVAL_2940;
  wire  _EVAL_2941;
  wire  _EVAL_2942;
  wire  _EVAL_2943;
  wire  _EVAL_2944;
  wire  _EVAL_2946;
  wire  _EVAL_2947;
  wire  _EVAL_2949;
  wire  _EVAL_2950;
  wire  _EVAL_2952;
  wire  _EVAL_2953;
  wire  _EVAL_2954;
  wire  _EVAL_2960;
  wire  _EVAL_2962;
  wire  _EVAL_2963;
  wire  _EVAL_2966;
  wire  _EVAL_2967;
  wire  _EVAL_2968;
  wire  _EVAL_2969;
  wire  _EVAL_2971;
  wire  _EVAL_2972;
  wire  _EVAL_2973;
  wire  _EVAL_2975;
  wire  _EVAL_2976;
  wire  _EVAL_2980;
  wire  _EVAL_2981;
  wire  _EVAL_2982;
  wire  _EVAL_2983;
  wire  _EVAL_2990;
  wire  _EVAL_2991;
  wire  _EVAL_2993;
  wire  _EVAL_2997;
  wire  _EVAL_2998;
  wire [3:0] _EVAL_2999;
  wire  _EVAL_3006;
  wire  _EVAL_3007;
  wire  _EVAL_3008;
  wire  _EVAL_3010;
  wire  _EVAL_3012;
  wire  _EVAL_3014;
  wire  _EVAL_3015;
  wire  _EVAL_3016;
  wire  _EVAL_3018;
  wire  _EVAL_3019;
  wire  _EVAL_3024;
  wire  _EVAL_3028;
  wire  _EVAL_3029;
  wire  _EVAL_3033;
  wire  _EVAL_3034;
  wire  _EVAL_3036;
  wire  _EVAL_3037;
  wire  _EVAL_3040;
  wire  _EVAL_3041;
  wire  _EVAL_3042;
  wire  _EVAL_3044;
  wire  _EVAL_3048;
  wire  _EVAL_3049;
  wire  _EVAL_3051;
  wire  _EVAL_3053;
  wire  _EVAL_3054;
  wire  _EVAL_3055;
  wire  _EVAL_3056;
  wire  _EVAL_3057;
  wire  _EVAL_3058;
  wire  _EVAL_3060;
  wire  _EVAL_3062;
  wire  _EVAL_3063;
  wire  _EVAL_3072;
  wire  _EVAL_3074;
  wire  _EVAL_3075;
  wire  _EVAL_3077;
  wire  _EVAL_3078;
  wire  _EVAL_3079;
  wire  _EVAL_3080;
  wire  _EVAL_3081;
  wire  _EVAL_3082;
  wire  _EVAL_3084;
  wire  _EVAL_3086;
  wire  _EVAL_3091;
  wire  _EVAL_3092;
  wire  _EVAL_3098;
  wire  _EVAL_3099;
  wire  _EVAL_3107;
  wire  _EVAL_3108;
  wire  _EVAL_3110;
  wire  _EVAL_3111;
  wire  _EVAL_3112;
  wire  _EVAL_3114;
  wire  _EVAL_3117;
  wire  _EVAL_3118;
  wire  _EVAL_3120;
  wire  _EVAL_3121;
  wire  _EVAL_3124;
  wire  _EVAL_3125;
  wire  _EVAL_3126;
  wire  _EVAL_3130;
  wire  _EVAL_3131;
  wire  _EVAL_3133;
  wire  _EVAL_3136;
  wire  _EVAL_3137;
  wire  _EVAL_3139;
  wire  _EVAL_3141;
  wire  _EVAL_3142;
  wire  _EVAL_3147;
  wire  _EVAL_3149;
  wire  _EVAL_3150;
  wire  _EVAL_3151;
  wire  _EVAL_3153;
  wire  _EVAL_3156;
  wire  _EVAL_3158;
  wire  _EVAL_3161;
  wire  _EVAL_3162;
  wire  _EVAL_3163;
  wire  _EVAL_3164;
  wire  _EVAL_3166;
  wire  _EVAL_3167;
  wire  _EVAL_3168;
  wire  _EVAL_3170;
  wire  _EVAL_3175;
  wire  _EVAL_3180;
  wire  _EVAL_3181;
  wire  _EVAL_3184;
  wire  _EVAL_3185;
  wire  _EVAL_3186;
  wire  _EVAL_3188;
  wire  _EVAL_3190;
  wire  _EVAL_3191;
  wire  _EVAL_3192;
  wire  _EVAL_3197;
  wire  _EVAL_3198;
  wire  _EVAL_3199;
  wire  _EVAL_3201;
  wire  _EVAL_3202;
  wire  _EVAL_3204;
  wire  _EVAL_3205;
  wire  _EVAL_3208;
  wire  _EVAL_3210;
  wire  _EVAL_3211;
  wire  _EVAL_3213;
  wire  _EVAL_3214;
  wire  _EVAL_3215;
  wire  _EVAL_3216;
  wire  _EVAL_3218;
  wire  _EVAL_3222;
  wire  _EVAL_3224;
  wire  _EVAL_3225;
  wire  _EVAL_3226;
  wire  _EVAL_3229;
  wire  _EVAL_3232;
  wire  _EVAL_3240;
  wire  _EVAL_3242;
  wire  _EVAL_3243;
  wire  _EVAL_3245;
  wire  _EVAL_3253;
  wire  _EVAL_3255;
  wire  _EVAL_3256;
  wire  _EVAL_3257;
  wire  _EVAL_3260;
  wire  _EVAL_3261;
  wire  _EVAL_3263;
  wire  _EVAL_3266;
  wire  _EVAL_3267;
  wire  _EVAL_3269;
  wire  _EVAL_3272;
  wire  _EVAL_3273;
  wire  _EVAL_3274;
  wire  _EVAL_3277;
  wire  _EVAL_3278;
  wire  _EVAL_3282;
  wire  _EVAL_3284;
  wire  _EVAL_3285;
  wire  _EVAL_3286;
  wire  _EVAL_3287;
  wire  _EVAL_3289;
  wire  _EVAL_3291;
  wire  _EVAL_3292;
  wire  _EVAL_3293;
  wire  _EVAL_3294;
  wire  _EVAL_3296;
  wire  _EVAL_3297;
  wire  _EVAL_3300;
  wire  _EVAL_3301;
  wire  _EVAL_3303;
  wire  _EVAL_3304;
  wire  _EVAL_3305;
  wire  _EVAL_3307;
  wire  _EVAL_3308;
  wire  _EVAL_3311;
  wire  _EVAL_3312;
  wire  _EVAL_3313;
  wire  _EVAL_3314;
  wire  _EVAL_3315;
  wire  _EVAL_3317;
  wire  _EVAL_3324;
  wire  _EVAL_3327;
  wire  _EVAL_3330;
  wire  _EVAL_3332;
  wire  _EVAL_3333;
  wire  _EVAL_3334;
  wire  _EVAL_3335;
  wire  _EVAL_3336;
  wire  _EVAL_3340;
  wire  _EVAL_3341;
  wire  _EVAL_3344;
  wire  _EVAL_3345;
  wire  _EVAL_3346;
  wire  _EVAL_3347;
  wire  _EVAL_3350;
  wire  _EVAL_3351;
  wire  _EVAL_3352;
  wire  _EVAL_3353;
  wire  _EVAL_3354;
  wire  _EVAL_3355;
  wire  _EVAL_3357;
  wire  _EVAL_3358;
  wire  _EVAL_3360;
  wire  _EVAL_3361;
  wire  _EVAL_3362;
  wire  _EVAL_3363;
  wire  _EVAL_3364;
  wire  _EVAL_3365;
  wire  _EVAL_3367;
  wire  _EVAL_3368;
  wire  _EVAL_3370;
  wire  _EVAL_3371;
  wire  _EVAL_3373;
  wire  _EVAL_3374;
  wire  _EVAL_3375;
  wire  _EVAL_3376;
  wire  _EVAL_3378;
  wire  _EVAL_3380;
  wire  _EVAL_3381;
  wire  _EVAL_3382;
  wire  _EVAL_3383;
  wire  _EVAL_3384;
  wire  _EVAL_3386;
  wire  _EVAL_3391;
  wire  _EVAL_3392;
  wire  _EVAL_3394;
  wire  _EVAL_3396;
  wire  _EVAL_3397;
  wire  _EVAL_3398;
  wire  _EVAL_3399;
  wire  _EVAL_3400;
  wire  _EVAL_3401;
  wire  _EVAL_3405;
  wire [9:0] _EVAL_3406;
  wire  _EVAL_3407;
  wire  _EVAL_3410;
  wire  _EVAL_3412;
  wire  _EVAL_3413;
  wire  _EVAL_3414;
  wire  _EVAL_3415;
  wire  _EVAL_3416;
  wire  _EVAL_3419;
  wire  _EVAL_3422;
  wire  _EVAL_3424;
  wire  _EVAL_3430;
  wire  _EVAL_3432;
  wire  _EVAL_3434;
  wire  _EVAL_3435;
  wire  _EVAL_3437;
  wire  _EVAL_3438;
  wire  _EVAL_3439;
  wire  _EVAL_3440;
  wire  _EVAL_3441;
  wire  _EVAL_3445;
  wire  _EVAL_3446;
  wire  _EVAL_3449;
  wire  _EVAL_3450;
  wire  _EVAL_3451;
  wire  _EVAL_3453;
  wire  _EVAL_3455;
  wire  _EVAL_3460;
  wire  _EVAL_3462;
  wire  _EVAL_3463;
  wire  _EVAL_3466;
  wire  _EVAL_3467;
  wire  _EVAL_3468;
  wire  _EVAL_3471;
  wire  _EVAL_3473;
  wire  _EVAL_3477;
  wire  _EVAL_3478;
  wire  _EVAL_3479;
  wire  _EVAL_3483;
  wire  _EVAL_3484;
  wire  _EVAL_3486;
  wire  _EVAL_3488;
  wire  _EVAL_3489;
  wire  _EVAL_3491;
  wire  _EVAL_3492;
  wire  _EVAL_3494;
  wire  _EVAL_3497;
  wire  _EVAL_3501;
  wire  _EVAL_3503;
  wire  _EVAL_3505;
  wire  _EVAL_3510;
  wire  _EVAL_3512;
  wire  _EVAL_3514;
  wire  _EVAL_3516;
  wire  _EVAL_3521;
  wire  _EVAL_3522;
  wire  _EVAL_3523;
  wire  _EVAL_3525;
  wire  _EVAL_3527;
  wire  _EVAL_3528;
  wire  _EVAL_3529;
  wire  _EVAL_3532;
  wire  _EVAL_3533;
  wire  _EVAL_3534;
  wire [10:0] _EVAL_3536;
  wire  _EVAL_3538;
  wire  _EVAL_3543;
  wire  _EVAL_3544;
  wire  _EVAL_3546;
  wire  _EVAL_3547;
  wire  _EVAL_3548;
  wire  _EVAL_3550;
  wire  _EVAL_3552;
  wire  _EVAL_3553;
  wire  _EVAL_3554;
  wire  _EVAL_3556;
  wire  _EVAL_3559;
  wire  _EVAL_3560;
  wire  _EVAL_3561;
  wire  _EVAL_3562;
  wire  _EVAL_3563;
  wire  _EVAL_3564;
  wire  _EVAL_3565;
  wire  _EVAL_3570;
  wire  _EVAL_3571;
  wire  _EVAL_3572;
  wire  _EVAL_3573;
  wire  _EVAL_3575;
  wire  _EVAL_3578;
  wire  _EVAL_3579;
  wire  _EVAL_3580;
  wire  _EVAL_3581;
  wire  _EVAL_3582;
  wire  _EVAL_3584;
  wire  _EVAL_3585;
  wire  _EVAL_3587;
  wire  _EVAL_3592;
  wire  _EVAL_3594;
  wire  _EVAL_3597;
  wire  _EVAL_3601;
  wire  _EVAL_3602;
  wire  _EVAL_3605;
  wire  _EVAL_3607;
  wire  _EVAL_3608;
  wire  _EVAL_3611;
  wire  _EVAL_3615;
  wire  _EVAL_3616;
  wire  _EVAL_3617;
  wire  _EVAL_3618;
  wire  _EVAL_3619;
  wire  _EVAL_3620;
  wire  _EVAL_3621;
  wire  _EVAL_3622;
  wire  _EVAL_3624;
  wire  _EVAL_3625;
  wire  _EVAL_3626;
  wire  _EVAL_3627;
  wire  _EVAL_3628;
  wire  _EVAL_3629;
  wire  _EVAL_3630;
  wire  _EVAL_3631;
  wire  _EVAL_3632;
  wire  _EVAL_3635;
  wire  _EVAL_3636;
  wire  _EVAL_3638;
  wire  _EVAL_3639;
  wire  _EVAL_3640;
  wire  _EVAL_3642;
  wire  _EVAL_3643;
  wire  _EVAL_3645;
  wire  _EVAL_3646;
  wire  _EVAL_3648;
  wire  _EVAL_3655;
  wire  _EVAL_3656;
  wire  _EVAL_3658;
  wire  _EVAL_3659;
  wire  _EVAL_3660;
  wire  _EVAL_3664;
  wire  _EVAL_3665;
  wire  _EVAL_3667;
  wire  _EVAL_3673;
  wire  _EVAL_3674;
  wire  _EVAL_3678;
  wire  _EVAL_3679;
  wire  _EVAL_3680;
  wire  _EVAL_3681;
  wire  _EVAL_3683;
  wire  _EVAL_3684;
  wire  _EVAL_3685;
  wire  _EVAL_3690;
  wire  _EVAL_3691;
  wire  _EVAL_3692;
  wire  _EVAL_3693;
  wire  _EVAL_3696;
  wire  _EVAL_3697;
  wire  _EVAL_3699;
  wire  _EVAL_3702;
  wire  _EVAL_3705;
  wire  _EVAL_3706;
  wire  _EVAL_3708;
  wire  _EVAL_3713;
  wire  _EVAL_3715;
  wire  _EVAL_3716;
  wire  _EVAL_3718;
  wire  _EVAL_3719;
  wire  _EVAL_3720;
  wire  _EVAL_3721;
  wire  _EVAL_3726;
  wire  _EVAL_3728;
  wire  _EVAL_3729;
  wire  _EVAL_3730;
  wire  _EVAL_3732;
  wire  _EVAL_3733;
  wire  _EVAL_3734;
  wire  _EVAL_3735;
  wire  _EVAL_3737;
  wire  _EVAL_3740;
  wire  _EVAL_3744;
  wire  _EVAL_3747;
  wire  _EVAL_3749;
  wire  _EVAL_3752;
  wire  _EVAL_3756;
  wire  _EVAL_3757;
  wire  _EVAL_3758;
  wire  _EVAL_3759;
  wire  _EVAL_3760;
  wire  _EVAL_3765;
  wire  _EVAL_3766;
  wire  _EVAL_3767;
  wire  _EVAL_3768;
  wire  _EVAL_3773;
  wire  _EVAL_3778;
  wire  _EVAL_3779;
  wire  _EVAL_3780;
  wire  _EVAL_3781;
  wire  _EVAL_3785;
  wire  _EVAL_3786;
  wire  _EVAL_3787;
  wire  _EVAL_3789;
  wire  _EVAL_3790;
  wire  _EVAL_3792;
  wire  _EVAL_3794;
  wire  _EVAL_3796;
  wire  _EVAL_3797;
  wire  _EVAL_3798;
  wire  _EVAL_3801;
  wire  _EVAL_3802;
  wire  _EVAL_3803;
  wire  _EVAL_3805;
  wire  _EVAL_3808;
  wire  _EVAL_3810;
  wire  _EVAL_3812;
  wire  _EVAL_3817;
  wire  _EVAL_3818;
  wire  _EVAL_3819;
  wire  _EVAL_3820;
  wire  _EVAL_3821;
  wire  _EVAL_3822;
  wire  _EVAL_3827;
  wire  _EVAL_3828;
  wire  _EVAL_3831;
  wire  _EVAL_3833;
  wire  _EVAL_3835;
  wire  _EVAL_3840;
  _EVAL_138_assert TLMonitor_1 (
    ._EVAL(TLMonitor_1__EVAL),
    ._EVAL_0(TLMonitor_1__EVAL_0),
    ._EVAL_1(TLMonitor_1__EVAL_1),
    ._EVAL_2(TLMonitor_1__EVAL_2),
    ._EVAL_3(TLMonitor_1__EVAL_3),
    ._EVAL_4(TLMonitor_1__EVAL_4),
    ._EVAL_5(TLMonitor_1__EVAL_5),
    ._EVAL_6(TLMonitor_1__EVAL_6),
    ._EVAL_7(TLMonitor_1__EVAL_7),
    ._EVAL_8(TLMonitor_1__EVAL_8),
    ._EVAL_9(TLMonitor_1__EVAL_9),
    ._EVAL_10(TLMonitor_1__EVAL_10),
    ._EVAL_11(TLMonitor_1__EVAL_11),
    ._EVAL_12(TLMonitor_1__EVAL_12),
    ._EVAL_13(TLMonitor_1__EVAL_13),
    ._EVAL_14(TLMonitor_1__EVAL_14)
  );
  _EVAL_137_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14)
  );
  assign _EVAL_3126 = _EVAL_678 & _EVAL_3391;
  assign _EVAL_2475 = _EVAL_2743[451];
  assign _EVAL_591 = _EVAL_2028 & _EVAL_3391;
  assign _EVAL_252 = _EVAL_2729 & _EVAL_2692;
  assign _EVAL_1882 = _EVAL_1782 & _EVAL_1808;
  assign _EVAL_2357 = _EVAL_652 & _EVAL_2474;
  assign _EVAL_3544 = _EVAL_177 & _EVAL_3670;
  assign _EVAL_1239 = _EVAL_168 & _EVAL_2474;
  assign _EVAL_3624 = _EVAL_1421 & _EVAL_3673;
  assign _EVAL_1404 = _EVAL_2743[2];
  assign _EVAL_2612 = _EVAL_3285 & _EVAL_2474;
  assign _EVAL_1453 = _EVAL_818 & _EVAL_2909;
  assign _EVAL_3181 = _EVAL_2043 & _EVAL_3673;
  assign _EVAL_142 = _EVAL_1782 & _EVAL_47;
  assign _EVAL_1727 = _EVAL_2743[12];
  assign _EVAL_1644 = _EVAL_1980 & _EVAL_1856;
  assign _EVAL_1980 = _EVAL_1782 & _EVAL_192;
  assign _EVAL_1780 = _EVAL_3794 & _EVAL_1856;
  assign _EVAL_779 = _EVAL_3201 & _EVAL_1856;
  assign _EVAL_1126 = _EVAL_1016 & _EVAL_1856;
  assign _EVAL_1719 = _EVAL_1740 & _EVAL_2909;
  assign _EVAL_593 = _EVAL_1524 & _EVAL_3391;
  assign _EVAL_2745 = _EVAL_2330 & _EVAL_1856;
  assign _EVAL_3242 = _EVAL_2093 & _EVAL_3391;
  assign _EVAL_1354 = _EVAL_575[7];
  assign _EVAL_1455 = _EVAL_2643 & _EVAL_2499;
  assign _EVAL_2375 = _EVAL_1765 & _EVAL_2909;
  assign _EVAL_3324 = _EVAL_2962 & _EVAL_3673;
  assign _EVAL_2427 = _EVAL_1967 & _EVAL_470;
  assign _EVAL_2751 = _EVAL_298 & _EVAL_3391;
  assign _EVAL_1573 = _EVAL_2019 & _EVAL_2474;
  assign _EVAL_1522 = _EVAL_1405 & _EVAL_3673;
  assign _EVAL_1456 = _EVAL_1782 & _EVAL_3484;
  assign _EVAL_2993 = _EVAL_682 & _EVAL_3391;
  assign _EVAL_691 = _EVAL_1644 & _EVAL_2909;
  assign _EVAL_2140 = _EVAL_2743[394];
  assign _EVAL_1614 = _EVAL_1782 & _EVAL_2576;
  assign _EVAL_2296 = _EVAL_2743[434];
  assign _EVAL_1373 = _EVAL_3361 & _EVAL_3391;
  assign _EVAL_1559 = _EVAL_507 & _EVAL_2474;
  assign _EVAL_831 = _EVAL_684 & _EVAL_3673;
  assign _EVAL_595 = _EVAL_2743[409];
  assign _EVAL_3505 = _EVAL_3674 & _EVAL_3673;
  assign _EVAL_1264 = _EVAL_1630 & _EVAL_1856;
  assign _EVAL_1990 = _EVAL_1716 & _EVAL_3673;
  assign _EVAL_2225 = _EVAL_575[22];
  assign _EVAL_2849 = _EVAL_706 & _EVAL_1856;
  assign _EVAL_2505 = _EVAL_850 & _EVAL_2474;
  assign _EVAL_1729 = _EVAL_2998 & _EVAL_2909;
  assign _EVAL_2205 = _EVAL_2059 & _EVAL_3391;
  assign _EVAL_1903 = _EVAL_2743[354];
  assign _EVAL_3263 = _EVAL_681 & _EVAL_120;
  assign _EVAL_3747 = _EVAL_988 & _EVAL_3391;
  assign _EVAL_1197 = _EVAL_1782 & _EVAL_1313;
  assign _EVAL_980 = _EVAL_1782 & _EVAL_1118;
  assign _EVAL_1967 = _EVAL_3485 & _EVAL_294;
  assign _EVAL_2441 = _EVAL_979 & _EVAL_3438;
  assign _EVAL_2112 = _EVAL_3728 & _EVAL_2474;
  assign _EVAL_3186 = _EVAL_1782 & _EVAL_3289;
  assign _EVAL_1670 = _EVAL_2745 & _EVAL_2474;
  assign _EVAL_888 = _EVAL_2743[219];
  assign _EVAL_224 = _EVAL_2743[427];
  assign _EVAL_3391 = _EVAL_3474 != 8'h0;
  assign _EVAL_1199 = _EVAL_1204 & _EVAL_2909;
  assign _EVAL_1868 = _EVAL_2743[280];
  assign _EVAL_718 = _EVAL_2972 & _EVAL_3391;
  assign _EVAL_796 = _EVAL_1246 & _EVAL_3673;
  assign _EVAL_2027 = _EVAL_2743[302];
  assign _EVAL_1385 = _EVAL_1439 & _EVAL_3673;
  assign _EVAL_2536 = _EVAL_100 & _EVAL_2909;
  assign _EVAL_293 = _EVAL_1780 & _EVAL_2474;
  assign _EVAL_2201 = _EVAL_1456 & _EVAL_1856;
  assign _EVAL_3635 = _EVAL_3024 & _EVAL_2474;
  assign _EVAL_446 = _EVAL_3347 & _EVAL_2909;
  assign _EVAL_1282 = _EVAL_1454 & _EVAL_1856;
  assign _EVAL_1491 = _EVAL_2743[408];
  assign _EVAL_1112 = _EVAL_287 & _EVAL_2909;
  assign _EVAL_2663 = _EVAL_2743[441];
  assign _EVAL_2824 = _EVAL_953 & _EVAL_2909;
  assign _EVAL_435 = _EVAL_3287 & _EVAL_3391;
  assign _EVAL_1916 = _EVAL_1094 & _EVAL_2474;
  assign _EVAL_3732 = _EVAL_2649 & _EVAL_2474;
  assign _EVAL_2273 = _EVAL_1272 & _EVAL_3673;
  assign TLMonitor__EVAL_14 = _EVAL_21;
  assign _EVAL_3648 = _EVAL_2093 & _EVAL_2474;
  assign _EVAL_3051 = _EVAL_1102 & _EVAL_2909;
  assign _EVAL_96 = _EVAL_2935 & _EVAL_2474;
  assign _EVAL_424 = _EVAL_1282 & _EVAL_2474;
  assign _EVAL_3450 = _EVAL_2743[492];
  assign _EVAL_2877 = _EVAL_575[17];
  assign _EVAL_1369 = _EVAL_2206 & _EVAL_2909;
  assign _EVAL_3216 = _EVAL_508 & _EVAL_1856;
  assign _EVAL_3016 = _EVAL_1782 & _EVAL_777;
  assign _EVAL_2525 = _EVAL_3186 & _EVAL_1856;
  assign _EVAL_1011 = _EVAL_2743[343];
  assign _EVAL_1777 = _EVAL_3757 & _EVAL_1886;
  assign TLMonitor__EVAL_3 = _EVAL_2;
  assign _EVAL_192 = _EVAL_2743[270];
  assign _EVAL_3150 = _EVAL_2743[363];
  assign _EVAL_3224 = _EVAL_2743[274];
  assign _EVAL_2230 = _EVAL_1165 & _EVAL_2474;
  assign _EVAL_82 = _EVAL_2729 & _EVAL_106;
  assign _EVAL_2661 = _EVAL_2423 & _EVAL_1856;
  assign _EVAL_2327 = _EVAL_979 & _EVAL_292;
  assign _EVAL_3049 = _EVAL_3185 & _EVAL_3673;
  assign _EVAL_885 = _EVAL_2214 | _EVAL_38;
  assign _EVAL_3730 = _EVAL_2743[355];
  assign _EVAL_1306 = _EVAL_3055 & _EVAL_2909;
  assign _EVAL_655 = _EVAL_1782 & _EVAL_1628;
  assign _EVAL_1179 = _EVAL_1794 & _EVAL_3391;
  assign _EVAL_2189 = _EVAL_74 & _EVAL_2474;
  assign _EVAL_3214 = _EVAL_1782 & _EVAL_326;
  assign _EVAL_2409 = _EVAL_140 & _EVAL_2474;
  assign _EVAL_646 = _EVAL_3621 & _EVAL_1856;
  assign _EVAL_427 = _EVAL_2743[337];
  assign _EVAL_2814 = _EVAL_2745 & _EVAL_2909;
  assign _EVAL_449 = _EVAL_575[5];
  assign _EVAL_425 = _EVAL_2743[315];
  assign _EVAL_1317 = _EVAL_575[14];
  assign _EVAL_2099 = _EVAL_2743[346];
  assign _EVAL_2511 = _EVAL_2068 & _EVAL_2909;
  assign TLMonitor_1__EVAL_8 = _EVAL_36;
  assign _EVAL_971 = _EVAL_1780 & _EVAL_3673;
  assign _EVAL_2147 = _EVAL_1189 & _EVAL_2474;
  assign _EVAL_2118 = _EVAL_2743[359];
  assign _EVAL_2778 = _EVAL_1915 & _EVAL_3391;
  assign _EVAL_2293 = _EVAL_623 & _EVAL_3391;
  assign _EVAL_3289 = _EVAL_2743[312];
  assign _EVAL_1464 = _EVAL_1329 & _EVAL_3673;
  assign _EVAL_626 = _EVAL_1782 & _EVAL_680;
  assign _EVAL_1579 = _EVAL_1282 & _EVAL_3391;
  assign _EVAL_673 = _EVAL_575[15:12];
  assign _EVAL_3611 = _EVAL_1309 & _EVAL_2474;
  assign _EVAL_1353 = _EVAL_2743[260];
  assign _EVAL_561 = _EVAL_1064 & _EVAL_2474;
  assign _EVAL_1157 = _EVAL_2743[414];
  assign TLMonitor_1__EVAL_14 = _EVAL_13;
  assign TLMonitor__EVAL_11 = _EVAL_15;
  assign _EVAL_3728 = _EVAL_2114 & _EVAL_1856;
  assign _EVAL_1388 = _EVAL_2743[435];
  assign _EVAL_657 = _EVAL_2743[267];
  assign _EVAL_164 = _EVAL_3245 & _EVAL_3673;
  assign _EVAL_44 = _EVAL_2229 & _EVAL_3673;
  assign _EVAL_3773 = _EVAL_1586 & _EVAL_3673;
  assign TLMonitor_1__EVAL_5 = _EVAL_14;
  assign _EVAL_3357 = _EVAL_3293 & _EVAL_1856;
  assign _EVAL_2234 = _EVAL_1782 & _EVAL_2740;
  assign _EVAL_3054 = _EVAL_2743[297];
  assign _EVAL_2798 = _EVAL_3055 & _EVAL_2474;
  assign _EVAL_1617 = _EVAL_3149 & _EVAL_2909;
  assign _EVAL_1638 = _EVAL_1782 & _EVAL_2003;
  assign _EVAL_2470 = _EVAL_298 & _EVAL_3673;
  assign _EVAL_1607 = _EVAL_2743[455];
  assign _EVAL_3383 = _EVAL_682 & _EVAL_2474;
  assign _EVAL_159 = _EVAL_3734 & _EVAL_3391;
  assign _EVAL_1996 = _EVAL_70 & _EVAL_1337;
  assign _EVAL_3253 = _EVAL_2055 & _EVAL_2474;
  assign _EVAL_226 = _EVAL_376 & _EVAL_2474;
  assign _EVAL_825 = _EVAL_2743[508];
  assign _EVAL_698 = _EVAL_2656 & _EVAL_3673;
  assign _EVAL_3108 = _EVAL_850 & _EVAL_3391;
  assign _EVAL_43 = _EVAL_518 & _EVAL_1856;
  assign _EVAL_523 = _EVAL_1915 & _EVAL_3673;
  assign _EVAL_1070 = _EVAL_2037 & _EVAL_3391;
  assign _EVAL_2846 = _EVAL_2743[424];
  assign _EVAL_1892 = _EVAL_418 & _EVAL_1856;
  assign _EVAL_1663 = _EVAL_2555 & _EVAL_2474;
  assign _EVAL_57 = _EVAL_1498 & _EVAL_3673;
  assign _EVAL_923 = _EVAL_2316 & _EVAL_2909;
  assign _EVAL_2139 = _EVAL_660 & _EVAL_1856;
  assign _EVAL_3401 = _EVAL_3726 & _EVAL_3391;
  assign _EVAL_1148 = _EVAL_2743[292];
  assign _EVAL_919 = _EVAL_2240 & _EVAL_1856;
  assign _EVAL_1908 = _EVAL_3185 & _EVAL_3391;
  assign _EVAL_2263 = _EVAL_2768 & _EVAL_2474;
  assign _EVAL_2267 = _EVAL_575[28:24];
  assign _EVAL_1866 = _EVAL_2043 & _EVAL_2474;
  assign _EVAL_1466 = _EVAL_2643 & _EVAL_1897;
  assign _EVAL_3733 = _EVAL_2743[478];
  assign _EVAL_3398 = _EVAL_575[10];
  assign _EVAL_2715 = _EVAL_1657 & _EVAL_2474;
  assign _EVAL_2723 = _EVAL_3802 & _EVAL_3391;
  assign _EVAL_1137 = _EVAL_3024 & _EVAL_3391;
  assign _EVAL_824 = _EVAL_3620 & _EVAL_2909;
  assign _EVAL_1929 = _EVAL_1391 & _EVAL_2474;
  assign _EVAL_695 = _EVAL_2743[463];
  assign _EVAL_3628 = _EVAL_3360 & _EVAL_2474;
  assign _EVAL_263 = _EVAL_1299 & _EVAL_3673;
  assign _EVAL_2722 = _EVAL_2743[442];
  assign _EVAL_2656 = _EVAL_50 & _EVAL_1856;
  assign _EVAL_582 = _EVAL_1782 & _EVAL_778;
  assign _EVAL_1927 = _EVAL_2738 & _EVAL_3673;
  assign _EVAL_2469 = _EVAL_3368 & _EVAL_2474;
  assign _EVAL_3451 = _EVAL_3361 & _EVAL_2909;
  assign _EVAL_3492 = _EVAL_1327 & _EVAL_2909;
  assign _EVAL_2833 = _EVAL_3780 & _EVAL_2909;
  assign _EVAL_2449 = _EVAL_2743[10];
  assign _EVAL_3056 = _EVAL_2203 & _EVAL_3391;
  assign _EVAL_508 = _EVAL_1782 & _EVAL_3422;
  assign _EVAL_3266 = _EVAL_2743[306];
  assign _EVAL_2983 = _EVAL_69 & _EVAL_3391;
  assign _EVAL_2065 = _EVAL_877 & _EVAL_2474;
  assign _EVAL_1973 = _EVAL_1963 & _EVAL_1856;
  assign _EVAL_521 = _EVAL_1785 & _EVAL_2188;
  assign _EVAL_2832 = _EVAL_3522 & _EVAL_2909;
  assign _EVAL_50 = _EVAL_1782 & _EVAL_3730;
  assign _EVAL_2468 = _EVAL_1782 & _EVAL_3266;
  assign _EVAL_213 = _EVAL_3691 & _EVAL_3391;
  assign _EVAL_811 = _EVAL_286 & _EVAL_3391;
  assign _EVAL_2443 = _EVAL_1986 & _EVAL_2474;
  assign _EVAL_2258 = _EVAL_2352 & _EVAL_3391;
  assign _EVAL_441 = _EVAL_2743[342];
  assign _EVAL_932 = _EVAL_1782 & _EVAL_1060;
  assign _EVAL_1216 = _EVAL_2064 & _EVAL_1856;
  assign _EVAL_678 = _EVAL_345 & _EVAL_1856;
  assign _EVAL_1088 = _EVAL_297 & _EVAL_3391;
  assign _EVAL_1657 = _EVAL_2696 & _EVAL_3670;
  assign _EVAL_1143 = _EVAL_2743[474];
  assign _EVAL_410 = _EVAL_780 & _EVAL_3391;
  assign _EVAL_1952 = _EVAL_2649 & _EVAL_3673;
  assign _EVAL_1848 = _EVAL_1542 & _EVAL_3391;
  assign _EVAL_1534 = _EVAL_1529 & _EVAL_3673;
  assign _EVAL_2071 = _EVAL_2554 & _EVAL_3673;
  assign _EVAL_3015 = _EVAL_1696 & _EVAL_1856;
  assign _EVAL_568 = _EVAL_1782 & _EVAL_2968;
  assign _EVAL_426 = _EVAL_1782 & _EVAL_2739;
  assign _EVAL_603 = _EVAL_2203 & _EVAL_2909;
  assign _EVAL_3394 = _EVAL_1782 & _EVAL_1890;
  assign _EVAL_580 = _EVAL_1782 & _EVAL_2433;
  assign _EVAL_2374 = _EVAL_2677 & _EVAL_897;
  assign _EVAL_105 = _EVAL_455 & _EVAL_3673;
  assign _EVAL_1932 = _EVAL_1188 & _EVAL_3391;
  assign _EVAL_3494 = _EVAL_337 & _EVAL_1856;
  assign _EVAL_3510 = _EVAL_1782 & _EVAL_1560;
  assign _EVAL_2514 = _EVAL_2743[329];
  assign _EVAL_897 = _EVAL_2363 != 32'h0;
  assign _EVAL_3744 = _EVAL_1782 & _EVAL_2465;
  assign _EVAL_3548 = _EVAL_1586 & _EVAL_2474;
  assign _EVAL_356 = _EVAL_83[9];
  assign _EVAL_1255 = _EVAL_1100 & _EVAL_1950;
  assign _EVAL_1686 = _EVAL_1782 & _EVAL_1011;
  assign _EVAL_1316 = _EVAL_1235 & _EVAL_3673;
  assign _EVAL_661 = _EVAL_1043 & _EVAL_2474;
  assign _EVAL_597 = _EVAL_2271 & _EVAL_2474;
  assign _EVAL_2070 = _EVAL_1216 & _EVAL_3391;
  assign _EVAL_294 = ~_EVAL_421;
  assign _EVAL_2933 = _EVAL_1782 & _EVAL_2158;
  assign _EVAL_2559 = _EVAL_99 & _EVAL_1856;
  assign _EVAL_453 = _EVAL_1782 & _EVAL_2839;
  assign _EVAL_2134 = _EVAL_3573 & _EVAL_1856;
  assign _EVAL_3414 = _EVAL_646 & _EVAL_2474;
  assign _EVAL_1708 = _EVAL_1782 & _EVAL_3006;
  assign _EVAL_2765 = _EVAL_3437 & _EVAL_1856;
  assign _EVAL_428 = _EVAL_1102 & _EVAL_2474;
  assign _EVAL_1610 = _EVAL_717 & _EVAL_2474;
  assign _EVAL_1447 = _EVAL_1782 & _EVAL_3137;
  assign _EVAL_947 = _EVAL_1782 & _EVAL_2283;
  assign _EVAL_3086 = _EVAL_646 & _EVAL_3673;
  assign _EVAL_2546 = _EVAL_3696 & _EVAL_3391;
  assign _EVAL_1288 = _EVAL_2555 & _EVAL_3391;
  assign _EVAL_3166 = _EVAL_1529 & _EVAL_2909;
  assign _EVAL_1858 = _EVAL_376 & _EVAL_3673;
  assign _EVAL_3594 = _EVAL_1782 & _EVAL_3033;
  assign _EVAL_2545 = _EVAL_2201 & _EVAL_3391;
  assign _EVAL_2549 = _EVAL_274 & _EVAL_2474;
  assign TLMonitor__EVAL_12 = {{2'd0}, _EVAL_3155};
  assign _EVAL_772 = _EVAL_2628 != 3'h0;
  assign _EVAL_2342 = _EVAL_1782 & _EVAL_676;
  assign _EVAL_2319 = _EVAL_717 & _EVAL_3391;
  assign _EVAL_2935 = _EVAL_1861 & _EVAL_1856;
  assign _EVAL_3024 = _EVAL_1962 & _EVAL_1856;
  assign _EVAL_465 = _EVAL_100 & _EVAL_3391;
  assign _EVAL_2679 = _EVAL_3726 & _EVAL_2474;
  assign _EVAL_2493 = _EVAL_1782 & _EVAL_243;
  assign _EVAL_1971 = _EVAL_575[7:4];
  assign _EVAL_1298 = _EVAL_3370 & _EVAL_3391;
  assign _EVAL_1262 = _EVAL_2352 & _EVAL_2474;
  assign _EVAL_999 = _EVAL_2020 & _EVAL_1856;
  assign _EVAL_3413 = _EVAL_3684 & _EVAL_2474;
  assign _EVAL_1904 = _EVAL_1363 & _EVAL_3391;
  assign _EVAL_3304 = _EVAL_2613 & _EVAL_2909;
  assign _EVAL_893 = _EVAL_235 & _EVAL_3391;
  assign _EVAL_743 = _EVAL_3245 & _EVAL_3391;
  assign _EVAL_136 = _EVAL_1782 & _EVAL_361;
  assign _EVAL_1333 = _EVAL_2119 & _EVAL_3673;
  assign _EVAL_2236 = _EVAL_1122 & _EVAL_1856;
  assign _EVAL_690 = _EVAL_1782 & _EVAL_2186;
  assign _EVAL_100 = _EVAL_1397 & _EVAL_1856;
  assign _EVAL_3308 = _EVAL_2743[485];
  assign _EVAL_3161 = _EVAL_1782 & _EVAL_1582;
  assign _EVAL_671 = _EVAL_2743[345];
  assign _EVAL_3699 = _EVAL_998 & _EVAL_2474;
  assign _EVAL_777 = _EVAL_2743[486];
  assign _EVAL_511 = _EVAL_1017 & _EVAL_1856;
  assign _EVAL_1414 = _EVAL_1882 & _EVAL_1856;
  assign _EVAL_1107 = _EVAL_2613 & _EVAL_3673;
  assign _EVAL_3466 = _EVAL_3594 & _EVAL_3670;
  assign _EVAL_3340 = _EVAL_3592 & _EVAL_2474;
  assign _EVAL_1786 = _EVAL_2743[457];
  assign _EVAL_3646 = _EVAL_720 & _EVAL_2474;
  assign _EVAL_1519 = _EVAL_137 & _EVAL_3391;
  assign _EVAL_1446 = _EVAL_2119 & _EVAL_2474;
  assign _EVAL_2047 = _EVAL_2743[272];
  assign _EVAL_507 = _EVAL_517 & _EVAL_1856;
  assign _EVAL_2825 = _EVAL_953 & _EVAL_3673;
  assign _EVAL_3534 = _EVAL_3416 & _EVAL_1856;
  assign _EVAL_2003 = _EVAL_2743[273];
  assign _EVAL_1053 = _EVAL_2743[382];
  assign _EVAL_1225 = _EVAL_2661 & _EVAL_3391;
  assign _EVAL_1577 = _EVAL_2643 & _EVAL_3836;
  assign _EVAL_515 = _EVAL_2729 & _EVAL_2639;
  assign _EVAL_3501 = _EVAL_3430 & _EVAL_3391;
  assign _EVAL_274 = _EVAL_3435 & _EVAL_1856;
  assign _EVAL_3756 = _EVAL_2765 & _EVAL_2909;
  assign _EVAL_1301 = _EVAL_929 & _EVAL_1856;
  assign _EVAL_918 = _EVAL_2305 & _EVAL_3391;
  assign _EVAL_2316 = _EVAL_932 & _EVAL_1856;
  assign _EVAL_950 = _EVAL_140 & _EVAL_3673;
  assign _EVAL_3820 = _EVAL_2743[446];
  assign _EVAL_3078 = _EVAL_2849 & _EVAL_3673;
  assign _EVAL_1413 = _EVAL_1782 & _EVAL_321;
  assign _EVAL_3716 = _EVAL_1964 & _EVAL_2474;
  assign _EVAL_3311 = _EVAL_2421 & _EVAL_2909;
  assign _EVAL_176 = _EVAL_3204 & _EVAL_1856;
  assign _EVAL_2465 = _EVAL_2743[493];
  assign _EVAL_3715 = _EVAL_3821 & _EVAL_2474;
  assign _EVAL_190 = _EVAL_2743[419];
  assign _EVAL_3605 = _EVAL_948 & _EVAL_3673;
  assign _EVAL_3560 = _EVAL_1165 & _EVAL_2909;
  assign _EVAL_2523 = _EVAL_2180 & _EVAL_2474;
  assign _EVAL_1595 = _EVAL_3151 & _EVAL_2909;
  assign _EVAL_2654 = _EVAL_3536 != 11'h0;
  assign _EVAL_2972 = _EVAL_770 & _EVAL_1856;
  assign _EVAL_3121 = _EVAL_979 & _EVAL_1919;
  assign _EVAL_914 = _EVAL_2743[426];
  assign _EVAL_1389 = _EVAL_1065 & _EVAL_3391;
  assign _EVAL_2936 = _EVAL_2126 & _EVAL_1856;
  assign _EVAL_738 = _EVAL_2953 & _EVAL_2474;
  assign _EVAL_3075 = _EVAL_3718 & _EVAL_3391;
  assign _EVAL_1946 = _EVAL_2119 & _EVAL_2909;
  assign _EVAL_2844 = _EVAL_548 & _EVAL_2474;
  assign _EVAL_3044 = _EVAL_1986 & _EVAL_2909;
  assign _EVAL_77 = _EVAL_1782 & _EVAL_2406;
  assign _EVAL_1997 = _EVAL_2729 & _EVAL_1634;
  assign _EVAL_1961 = _EVAL_447 & _EVAL_1856;
  assign _EVAL_3175 = _EVAL_1782 & _EVAL_1388;
  assign _EVAL_1938 = _EVAL_1457 & _EVAL_1856;
  assign _EVAL_2916 = _EVAL_1973 & _EVAL_2909;
  assign _EVAL_1064 = _EVAL_3744 & _EVAL_1856;
  assign _EVAL_3336 = _EVAL_2600 & _EVAL_3673;
  assign _EVAL_2221 = _EVAL_3080 & _EVAL_2474;
  assign _EVAL_504 = _EVAL_1782 & _EVAL_2664;
  assign _EVAL_3296 = _EVAL_576 & _EVAL_2909;
  assign _EVAL_562 = _EVAL_2478 & _EVAL_3391;
  assign _EVAL_677 = _EVAL_652 & _EVAL_2909;
  assign _EVAL_1310 = _EVAL_3494 & _EVAL_3391;
  assign _EVAL_394 = _EVAL_2316 & _EVAL_3673;
  assign _EVAL_660 = _EVAL_1782 & _EVAL_2717;
  assign _EVAL_1692 = _EVAL_3728 & _EVAL_3673;
  assign _EVAL_3522 = _EVAL_2257 & _EVAL_1856;
  assign _EVAL_2575 = _EVAL_1782 & _EVAL_1607;
  assign _EVAL_1757 = _EVAL_3620 & _EVAL_3391;
  assign _EVAL_1202 = _EVAL_1986 & _EVAL_3391;
  assign _EVAL_1178 = _EVAL_2139 & _EVAL_3673;
  assign _EVAL_3397 = _EVAL_818 & _EVAL_3391;
  assign _EVAL_314 = _EVAL_336 & _EVAL_1856;
  assign _EVAL_2231 = _EVAL_1782 & _EVAL_64;
  assign _EVAL_604 = _EVAL_1782 & _EVAL_1353;
  assign _EVAL_2717 = _EVAL_2743[262];
  assign _EVAL_2467 = _EVAL_1794 & _EVAL_3673;
  assign TLMonitor_1__EVAL_13 = _EVAL;
  assign _EVAL_112 = _EVAL_872 & _EVAL_2909;
  assign _EVAL_2098 = _EVAL_314 & _EVAL_2474;
  assign _EVAL_1094 = _EVAL_2954 & _EVAL_1856;
  assign _EVAL_3625 = _EVAL_3360 & _EVAL_3391;
  assign _EVAL_273 = _EVAL_684 & _EVAL_3391;
  assign _EVAL_2942 = _EVAL_1172 & _EVAL_3391;
  assign _EVAL_974 = _EVAL_3024 & _EVAL_2909;
  assign _EVAL_423 = _EVAL_3368 & _EVAL_3673;
  assign _EVAL_786 = _EVAL_1294 & _EVAL_3391;
  assign _EVAL_3620 = _EVAL_3678 & _EVAL_1856;
  assign _EVAL_3345 = _EVAL_1638 & _EVAL_1856;
  assign _EVAL_3378 = _EVAL_201 & _EVAL_3391;
  assign _EVAL_1207 = _EVAL_1484 & _EVAL_1856;
  assign _EVAL_361 = _EVAL_2743[422];
  assign _EVAL_2779 = _EVAL_2936 & _EVAL_2909;
  assign _EVAL_3690 = _EVAL_1782 & _EVAL_2846;
  assign _EVAL_2796 = _EVAL_3779 & _EVAL_3391;
  assign _EVAL_3405 = _EVAL_550 & _EVAL_2909;
  assign _EVAL_292 = _EVAL_2404 != 12'h0;
  assign _EVAL_2922 = _EVAL_1531 & _EVAL_1856;
  assign _EVAL_1756 = _EVAL_201 & _EVAL_2474;
  assign _EVAL_687 = _EVAL_2729 & _EVAL_1354;
  assign _EVAL_1808 = _EVAL_2743[433];
  assign _EVAL_2603 = _EVAL_3232 & _EVAL_3391;
  assign _EVAL_708 = _EVAL_1782 & _EVAL_3768;
  assign _EVAL_1432 = _EVAL_2342 & _EVAL_3670;
  assign _EVAL_2982 = _EVAL_2743[397];
  assign _EVAL_2947 = _EVAL_2201 & _EVAL_2909;
  assign _EVAL_373 = _EVAL_1299 & _EVAL_3391;
  assign _EVAL_1214 = _EVAL_3370 & _EVAL_2909;
  assign _EVAL_517 = _EVAL_1782 & _EVAL_1945;
  assign TLMonitor__EVAL_13 = _EVAL_41;
  assign _EVAL_839 = _EVAL_1340 & _EVAL_2909;
  assign _EVAL_564 = _EVAL_1782 & _EVAL_1157;
  assign _EVAL_3547 = _EVAL_1126 & _EVAL_2909;
  assign _EVAL_3147 = _EVAL_1782 & _EVAL_2389;
  assign _EVAL_1028 = _EVAL_1189 & _EVAL_3673;
  assign _EVAL_2968 = _EVAL_2743[389];
  assign _EVAL_1811 = _EVAL_988 & _EVAL_2474;
  assign _EVAL_383 = _EVAL_70 & _EVAL_1948;
  assign TLMonitor__EVAL_8 = _EVAL_33;
  assign _EVAL_2338 = _EVAL_1748 & _EVAL_1856;
  assign _EVAL_1074 = _EVAL_2910 & _EVAL_3391;
  assign _EVAL_804 = _EVAL_2236 & _EVAL_2909;
  assign _EVAL_1601 = _EVAL_673 != 4'h0;
  assign _EVAL_3133 = _EVAL_2743[378];
  assign _EVAL_443 = _EVAL_2743[291];
  assign _EVAL_2053 = _EVAL_1100 & _EVAL_2654;
  assign _EVAL_3293 = _EVAL_1782 & _EVAL_2834;
  assign _EVAL_1850 = _EVAL_2743[16];
  assign _EVAL_2863 = _EVAL_548 & _EVAL_3391;
  assign _EVAL_3660 = _EVAL_2935 & _EVAL_2909;
  assign _EVAL_3354 = _EVAL_2401 & _EVAL_2909;
  assign _EVAL_1981 = _EVAL_3587 & _EVAL_3391;
  assign _EVAL_2198 = _EVAL_1782 & _EVAL_3019;
  assign _EVAL_2023 = _EVAL_2799 & _EVAL_3673;
  assign TLMonitor__EVAL_10 = _EVAL_30;
  assign _EVAL_892 = _EVAL_1204 & _EVAL_3391;
  assign _EVAL_3215 = _EVAL_1094 & _EVAL_3391;
  assign _EVAL_2137 = _EVAL_1782 & _EVAL_2204;
  assign _EVAL_245 = _EVAL_2401 & _EVAL_3673;
  assign _EVAL_953 = _EVAL_2760 & _EVAL_1856;
  assign _EVAL_2710 = _EVAL_2743[473];
  assign _EVAL_3618 = _EVAL_3691 & _EVAL_3673;
  assign _EVAL_1524 = _EVAL_2848 & _EVAL_1856;
  assign _EVAL_85 = _EVAL_1765 & _EVAL_3391;
  assign _EVAL_1542 = _EVAL_444 & _EVAL_1856;
  assign _EVAL_1119 = _EVAL_1782 & _EVAL_1379;
  assign _EVAL_1210 = _EVAL_1782 & _EVAL_3042;
  assign _EVAL_3521 = _EVAL_1782 & _EVAL_2802;
  assign _EVAL_3563 = _EVAL_1340 & _EVAL_3391;
  assign _EVAL_2167 = _EVAL_1782 & _EVAL_1818;
  assign _EVAL_2388 = _EVAL_2743[483];
  assign _EVAL_3525 = _EVAL_2201 & _EVAL_2474;
  assign _EVAL_269 = _EVAL_2525 & _EVAL_3673;
  assign _EVAL_155 = _EVAL_322 & _EVAL_2474;
  assign _EVAL_3008 = _EVAL_3608 & _EVAL_3673;
  assign _EVAL_1836 = _EVAL_2738 & _EVAL_2909;
  assign _EVAL_709 = _EVAL_1414 & _EVAL_2909;
  assign _EVAL_681 = _EVAL_1466 & _EVAL_2188;
  assign _EVAL_3019 = _EVAL_2743[319];
  assign _EVAL_2762 = _EVAL_1782 & _EVAL_2382;
  assign _EVAL_712 = _EVAL_2227 & _EVAL_1856;
  assign _EVAL_349 = _EVAL_575[18];
  assign _EVAL_2976 = _EVAL_511 & _EVAL_2909;
  assign _EVAL_70 = _EVAL_1577 & _EVAL_2655;
  assign _EVAL_1349 = _EVAL_1782 & _EVAL_3831;
  assign _EVAL_2792 = _EVAL_2643 & _EVAL_3564;
  assign _EVAL_3592 = _EVAL_3257 & _EVAL_1856;
  assign _EVAL_3817 = _EVAL_1424 & _EVAL_1856;
  assign _EVAL_3484 = _EVAL_2743[410];
  assign _EVAL_1865 = _EVAL_3718 & _EVAL_2909;
  assign _EVAL_1825 = _EVAL_575[13];
  assign _EVAL_240 = _EVAL_2180 & _EVAL_3391;
  assign _EVAL_1323 = _EVAL_1432 & _EVAL_3673;
  assign _EVAL_1711 = _EVAL_3734 & _EVAL_3673;
  assign _EVAL_2868 = _EVAL_3351 & _EVAL_2474;
  assign _EVAL_1582 = _EVAL_2743[509];
  assign _EVAL_1917 = _EVAL_2743[295];
  assign _EVAL_3720 = _EVAL_1235 & _EVAL_3391;
  assign _EVAL_1775 = _EVAL_988 & _EVAL_2909;
  assign _EVAL_812 = _EVAL_1656 & _EVAL_2909;
  assign _EVAL_2719 = _EVAL_2743[313];
  assign _EVAL_770 = _EVAL_1782 & _EVAL_2719;
  assign _EVAL_2785 = _EVAL_3229 & _EVAL_2474;
  assign _EVAL_1371 = _EVAL_3357 & _EVAL_3391;
  assign _EVAL_3471 = _EVAL_1381 & _EVAL_3391;
  assign _EVAL_3229 = _EVAL_1119 & _EVAL_1856;
  assign _EVAL_1828 = _EVAL_646 & _EVAL_2909;
  assign _EVAL_232 = _EVAL_2743[290];
  assign _EVAL_1364 = _EVAL_2525 & _EVAL_3391;
  assign _EVAL_3158 = _EVAL_137 & _EVAL_2909;
  assign _EVAL_693 = _EVAL_1524 & _EVAL_2909;
  assign _EVAL_827 = _EVAL_2953 & _EVAL_3673;
  assign _EVAL_911 = _EVAL_1413 & _EVAL_1856;
  assign _EVAL_3752 = _EVAL_3691 & _EVAL_2474;
  assign _EVAL_1797 = _EVAL_1356 & _EVAL_2474;
  assign _EVAL_2925 = _EVAL_2743[372];
  assign _EVAL_1497 = _EVAL_1782 & _EVAL_1305;
  assign _EVAL_2971 = _EVAL_3817 & _EVAL_2474;
  assign _EVAL_3053 = _EVAL_1783 & _EVAL_3673;
  assign _EVAL_3808 = _EVAL_3802 & _EVAL_3673;
  assign _EVAL_335 = _EVAL_1793 & _EVAL_3673;
  assign _EVAL_2997 = _EVAL_288 & _EVAL_3391;
  assign _EVAL_1829 = _EVAL_878 & _EVAL_2909;
  assign _EVAL_3312 = _EVAL_2743[445];
  assign _EVAL_3225 = _EVAL_2253 & _EVAL_2474;
  assign _EVAL_1382 = _EVAL_201 & _EVAL_2909;
  assign _EVAL_2257 = _EVAL_1782 & _EVAL_3048;
  assign _EVAL_3768 = _EVAL_2743[324];
  assign _EVAL_798 = _EVAL_2743[437];
  assign _EVAL_261 = _EVAL_2922 & _EVAL_2909;
  assign _EVAL_2282 = _EVAL_216 & _EVAL_1856;
  assign _EVAL_3554 = _EVAL_1264 & _EVAL_2909;
  assign _EVAL_684 = _EVAL_3198 & _EVAL_1856;
  assign _EVAL_3664 = _EVAL_2316 & _EVAL_2474;
  assign _EVAL_1781 = _EVAL_3527 & _EVAL_2474;
  assign _EVAL_1924 = _EVAL_1421 & _EVAL_2474;
  assign _EVAL_3422 = _EVAL_2743[400];
  assign _EVAL_1760 = _EVAL_2743[376];
  assign _EVAL_1498 = _EVAL_3510 & _EVAL_1856;
  assign _EVAL_413 = _EVAL_1782 & _EVAL_495;
  assign _EVAL_663 = _EVAL_998 & _EVAL_3391;
  assign _EVAL_2114 = _EVAL_1782 & _EVAL_798;
  assign _EVAL_3313 = _EVAL_1765 & _EVAL_2474;
  assign _EVAL_1976 = _EVAL_2034 & _EVAL_3391;
  assign _EVAL_2278 = _EVAL_2353 & _EVAL_2909;
  assign _EVAL_3412 = _EVAL_726 & _EVAL_2909;
  assign _EVAL_161 = _EVAL_2743[322];
  assign _EVAL_2960 = _EVAL_2743[362];
  assign _EVAL_1203 = _EVAL_596 & _EVAL_3391;
  assign _EVAL_3098 = _EVAL_3361 & _EVAL_2474;
  assign _EVAL_2154 = _EVAL_1782 & _EVAL_1056;
  assign _EVAL_2203 = _EVAL_1500 & _EVAL_1856;
  assign _EVAL_2195 = _EVAL_2972 & _EVAL_2909;
  assign _EVAL_1596 = _EVAL_1782 & _EVAL_3079;
  assign _EVAL_315 = _EVAL_3347 & _EVAL_2474;
  assign _EVAL_1457 = _EVAL_1782 & _EVAL_440;
  assign _EVAL_3386 = _EVAL_140 & _EVAL_2909;
  assign _EVAL_1642 = _EVAL_2743[371];
  assign _EVAL_1840 = _EVAL_2743[220];
  assign _EVAL_2909 = _EVAL_3750 != 8'h0;
  assign _EVAL_3211 = _EVAL_70 & _EVAL_1195;
  assign _EVAL_3486 = _EVAL_2253 & _EVAL_3391;
  assign _EVAL_437 = _EVAL_818 & _EVAL_3673;
  assign _EVAL_731 = _EVAL_2353 & _EVAL_3673;
  assign _EVAL_2026 = _EVAL_2743[387];
  assign _EVAL_3621 = _EVAL_1782 & _EVAL_1868;
  assign _EVAL_2963 = _EVAL_1656 & _EVAL_2474;
  assign _EVAL_1847 = _EVAL_2743[293];
  assign _EVAL_2692 = _EVAL_575[6];
  assign _EVAL_2733 = _EVAL_1782 & _EVAL_1955;
  assign _EVAL_2998 = _EVAL_1090 & _EVAL_1856;
  assign _EVAL_1751 = _EVAL_2743[261];
  assign _EVAL_2283 = _EVAL_2743[370];
  assign _EVAL_2490 = _EVAL_2743[6];
  assign _EVAL_3767 = _EVAL_305 & _EVAL_2909;
  assign _EVAL_609 = _EVAL_717 & _EVAL_2909;
  assign _EVAL_2142 = _EVAL_1740 & _EVAL_3673;
  assign _EVAL_1313 = _EVAL_2743[256];
  assign _EVAL_369 = _EVAL_2559 & _EVAL_3391;
  assign _EVAL_3080 = _EVAL_2991 & _EVAL_1856;
  assign _EVAL_729 = _EVAL_1126 & _EVAL_3391;
  assign _EVAL_2408 = _EVAL_535 & _EVAL_2909;
  assign _EVAL_3114 = _EVAL_2259 & _EVAL_1856;
  assign _EVAL_1118 = _EVAL_2743[341];
  assign _EVAL_253 = _EVAL_3149 & _EVAL_3391;
  assign _EVAL_1634 = _EVAL_575[19];
  assign _EVAL_2425 = _EVAL_582 & _EVAL_1856;
  assign _EVAL_2582 = _EVAL_1235 & _EVAL_2909;
  assign _EVAL_1648 = _EVAL_1782 & _EVAL_1355;
  assign _EVAL_2204 = _EVAL_2743[477];
  assign _EVAL_2675 = _EVAL_1788 & _EVAL_3670;
  assign _EVAL_2678 = _EVAL_3728 & _EVAL_2909;
  assign _EVAL_296 = _EVAL_2962 & _EVAL_2909;
  assign _EVAL_2243 = _EVAL_1065 & _EVAL_3673;
  assign _EVAL_688 = _EVAL_176 & _EVAL_2909;
  assign _EVAL_3432 = _EVAL_2743[468];
  assign _EVAL_2260 = _EVAL_1782 & _EVAL_3308;
  assign _EVAL_462 = _EVAL_1189 & _EVAL_3391;
  assign _EVAL_2181 = _EVAL_322 & _EVAL_3673;
  assign _EVAL_194 = _EVAL_173 & _EVAL_2909;
  assign _EVAL_404 = _EVAL_3561 & _EVAL_2474;
  assign _EVAL_844 = _EVAL_1782 & _EVAL_350;
  assign _EVAL_146 = _EVAL_3466 & _EVAL_2909;
  assign _EVAL_2606 = _EVAL_3345 & _EVAL_2474;
  assign _EVAL_3726 = _EVAL_716 & _EVAL_1856;
  assign _EVAL_2164 = _EVAL_550 & _EVAL_2474;
  assign _EVAL_1560 = _EVAL_2743[497];
  assign _EVAL_3084 = _EVAL_1951 & _EVAL_2474;
  assign _EVAL_3627 = _EVAL_1783 & _EVAL_2474;
  assign _EVAL_3587 = _EVAL_2826 & _EVAL_1856;
  assign _EVAL_1267 = _EVAL_3529 & _EVAL_2909;
  assign _EVAL_1810 = _EVAL_1204 & _EVAL_3673;
  assign _EVAL_2799 = _EVAL_2199 & _EVAL_1856;
  assign _EVAL_1254 = _EVAL_74 & _EVAL_3391;
  assign _EVAL_2038 = _EVAL_2084 & _EVAL_2474;
  assign _EVAL_2752 = _EVAL_2729 & _EVAL_349;
  assign _EVAL_933 = _EVAL_1782 & _EVAL_3729;
  assign _EVAL_478 = _EVAL_977 & _EVAL_3673;
  assign _EVAL_2048 = _EVAL_2743[381];
  assign _EVAL_3333 = _EVAL_3399 & _EVAL_2909;
  assign _EVAL_667 = _EVAL_568 & _EVAL_1856;
  assign _EVAL_1502 = _EVAL_3534 & _EVAL_2474;
  assign _EVAL_3789 = _EVAL_2849 & _EVAL_3391;
  assign _EVAL_500 = _EVAL_2430 & _EVAL_1523;
  assign _EVAL_3167 = _EVAL_513 & _EVAL_1856;
  assign _EVAL_716 = _EVAL_1782 & _EVAL_2047;
  assign _EVAL_1359 = _EVAL_2817 & _EVAL_3673;
  assign _EVAL_2044 = _EVAL_3803 & _EVAL_3391;
  assign _EVAL_2969 = _EVAL_1954 & _EVAL_897;
  assign _EVAL_1381 = _EVAL_1295 & _EVAL_1856;
  assign _EVAL_305 = _EVAL_2349 & _EVAL_3670;
  assign _EVAL_3130 = _EVAL_1794 & _EVAL_2909;
  assign _EVAL_3445 = _EVAL_2729 & _EVAL_2877;
  assign _EVAL_3060 = _EVAL_1405 & _EVAL_2909;
  assign _EVAL_199 = _EVAL_286 & _EVAL_2474;
  assign _EVAL_1309 = _EVAL_855 & _EVAL_1856;
  assign _EVAL_2498 = _EVAL_2743[286];
  assign _EVAL_1059 = _EVAL_2743[265];
  assign _EVAL_2576 = _EVAL_2743[271];
  assign _EVAL_778 = _EVAL_2743[404];
  assign _EVAL_2638 = _EVAL_2880 & _EVAL_3391;
  assign _EVAL_1060 = _EVAL_2743[309];
  assign _EVAL_2685 = _EVAL_717 & _EVAL_3673;
  assign _EVAL_3616 = _EVAL_2953 & _EVAL_3391;
  assign _EVAL_1061 = _EVAL_575[15:1];
  assign _EVAL_3491 = _EVAL_3760 & _EVAL_3673;
  assign _EVAL_3327 = _EVAL_1679 & _EVAL_1856;
  assign _EVAL_2341 = _EVAL_1172 & _EVAL_3673;
  assign _EVAL_2903 = _EVAL_445 & _EVAL_2909;
  assign _EVAL_714 = _EVAL_2555 & _EVAL_2909;
  assign _EVAL_1111 = _EVAL_2743[436];
  assign _EVAL_1398 = _EVAL_3734 & _EVAL_2909;
  assign _EVAL_1526 = _EVAL_3726 & _EVAL_2909;
  assign _EVAL_3255 = _EVAL_235 & _EVAL_2909;
  assign _EVAL_838 = _EVAL_2046 & _EVAL_3391;
  assign _EVAL_641 = _EVAL_877 & _EVAL_3673;
  assign _EVAL_3260 = _EVAL_3527 & _EVAL_3673;
  assign _EVAL_227 = _EVAL_999 & _EVAL_2474;
  assign _EVAL_3693 = _EVAL_3696 & _EVAL_2909;
  assign _EVAL_3168 = _EVAL_1782 & _EVAL_1847;
  assign _EVAL_3455 = _EVAL_2559 & _EVAL_3673;
  assign _EVAL_2187 = _EVAL_3494 & _EVAL_2474;
  assign _EVAL_2170 = _EVAL_2568 & _EVAL_2909;
  assign _EVAL_2953 = _EVAL_3840 & _EVAL_1856;
  assign _EVAL_2244 = _EVAL_2765 & _EVAL_3673;
  assign _EVAL_2592 = _EVAL_2743[498];
  assign _EVAL_2370 = _EVAL_2743[461];
  assign _EVAL_1600 = _EVAL_2729 & _EVAL_1940;
  assign _EVAL_2671 = _EVAL_2743[304];
  assign _EVAL_1055 = _EVAL_3532 & _EVAL_3391;
  assign _EVAL_3350 = _EVAL_2428 & _EVAL_3673;
  assign _EVAL_287 = _EVAL_3758 & _EVAL_1856;
  assign _EVAL_2530 = _EVAL_1503 & _EVAL_2474;
  assign _EVAL_3673 = _EVAL_2662 != 8'h0;
  assign _EVAL_553 = _EVAL_1782 & _EVAL_1048;
  assign _EVAL_2690 = _EVAL_1656 & _EVAL_3391;
  assign _EVAL_3284 = ~_EVAL_3425;
  assign _EVAL_2739 = _EVAL_2743[411];
  assign _EVAL_834 = _EVAL_3365 & _EVAL_3673;
  assign _EVAL_2856 = _EVAL_2743[503];
  assign _EVAL_2902 = _EVAL_3358 & _EVAL_2474;
  assign _EVAL_826 = _EVAL_1782 & _EVAL_746;
  assign _EVAL_1042 = _EVAL_1414 & _EVAL_2474;
  assign _EVAL_86 = _EVAL_507 & _EVAL_2909;
  assign _EVAL_1649 = _EVAL_3351 & _EVAL_2909;
  assign _EVAL_352 = _EVAL_2743[504];
  assign _EVAL_1444 = _EVAL_1782 & _EVAL_357;
  assign _EVAL_535 = _EVAL_262 & _EVAL_1856;
  assign _EVAL_973 = _EVAL_2743[489];
  assign _EVAL_3528 = _EVAL_305 & _EVAL_2474;
  assign _EVAL_1428 = _EVAL_1782 & _EVAL_3450;
  assign _EVAL_2767 = _EVAL_3597 & _EVAL_3673;
  assign _EVAL_1995 = ~_EVAL_470;
  assign _EVAL_1346 = _EVAL_208 & _EVAL_2909;
  assign _EVAL_706 = _EVAL_1782 & _EVAL_3579;
  assign _EVAL_1168 = _EVAL_3327 & _EVAL_2909;
  assign _EVAL_2784 = _EVAL_398 & _EVAL_2909;
  assign _EVAL_1308 = _EVAL_3527 & _EVAL_2909;
  assign _EVAL_2639 = _EVAL_575[11];
  assign _EVAL_2835 = _EVAL_3645 & _EVAL_2909;
  assign _EVAL_1776 = _EVAL_550 & _EVAL_3673;
  assign _EVAL_2869 = _EVAL_1272 & _EVAL_2474;
  assign _EVAL_438 = _EVAL_2743[502];
  assign _EVAL_1907 = _EVAL_1586 & _EVAL_2909;
  assign _EVAL_1918 = _EVAL_2303 & _EVAL_2909;
  assign _EVAL_3136 = _EVAL_3532 & _EVAL_3673;
  assign _EVAL_983 = _EVAL_3216 & _EVAL_2909;
  assign _EVAL_3582 = _EVAL_2718 & _EVAL_3391;
  assign _EVAL_1764 = _EVAL_2661 & _EVAL_2474;
  assign _EVAL_939 = _EVAL_3285 & _EVAL_3673;
  assign _EVAL_3137 = _EVAL_2743[479];
  assign _EVAL_531 = _EVAL_2059 & _EVAL_2909;
  assign _EVAL_1802 = _EVAL_2525 & _EVAL_2909;
  assign _EVAL_2133 = _EVAL_1938 & _EVAL_3673;
  assign _EVAL_3396 = _EVAL_1782 & _EVAL_3410;
  assign _EVAL_2640 = _EVAL_850 & _EVAL_3673;
  assign _EVAL_2105 = _EVAL_3608 & _EVAL_2909;
  assign _EVAL_80 = _EVAL_2743[278];
  assign _EVAL_2652 = _EVAL_2028 & _EVAL_2909;
  assign _EVAL_3697 = _EVAL_2396 & _EVAL_3673;
  assign _EVAL_2473 = _EVAL_1329 & _EVAL_3391;
  assign _EVAL_2696 = _EVAL_1782 & _EVAL_1372;
  assign _EVAL_3012 = _EVAL_1782 & _EVAL_1300;
  assign _EVAL_3347 = _EVAL_1342 & _EVAL_3670;
  assign _EVAL_1733 = _EVAL_3821 & _EVAL_3673;
  assign _EVAL_1726 = _EVAL_1188 & _EVAL_3673;
  assign _EVAL_3821 = _EVAL_3164 & _EVAL_1856;
  assign _EVAL_2259 = _EVAL_1782 & _EVAL_2241;
  assign _EVAL_2492 = _EVAL_2743[448];
  assign _EVAL_466 = _EVAL_2059 & _EVAL_3673;
  assign _EVAL_289 = _EVAL_2305 & _EVAL_3673;
  assign _EVAL_2918 = _EVAL_1614 & _EVAL_1856;
  assign _EVAL_3665 = _EVAL_1782 & _EVAL_166;
  assign _EVAL_1703 = _EVAL_1782 & _EVAL_2622;
  assign _EVAL_2999 = _EVAL_575[23:20];
  assign _EVAL_1361 = _EVAL_2019 & _EVAL_3391;
  assign _EVAL_2007 = _EVAL_3494 & _EVAL_2909;
  assign _EVAL_2304 = _EVAL_3835 & _EVAL_3673;
  assign _EVAL_221 = _EVAL_3684 & _EVAL_3673;
  assign _EVAL_1623 = _EVAL_1782 & _EVAL_438;
  assign _EVAL_652 = _EVAL_1956 & _EVAL_3670;
  assign _EVAL_2323 = _EVAL_3370 & _EVAL_2474;
  assign _EVAL_2515 = _EVAL_1782 & _EVAL_1548;
  assign _EVAL_3082 = _EVAL_3812 & _EVAL_3673;
  assign _EVAL_3243 = _EVAL_1783 & _EVAL_3391;
  assign _EVAL_2889 = _EVAL_89 & _EVAL_2474;
  assign _EVAL_355 = _EVAL_2790 & _EVAL_1856;
  assign _EVAL_1253 = _EVAL_1780 & _EVAL_3391;
  assign _EVAL_3696 = _EVAL_3665 & _EVAL_1856;
  assign _EVAL_2239 = _EVAL_2134 & _EVAL_2474;
  assign _EVAL_2380 = _EVAL_1524 & _EVAL_2474;
  assign _EVAL_3584 = _EVAL_1635 & _EVAL_2474;
  assign _EVAL_1801 = _EVAL_2729 & _EVAL_3681;
  assign _EVAL_2068 = _EVAL_2122 & _EVAL_1856;
  assign _EVAL_1005 = _EVAL_1421 & _EVAL_2909;
  assign _EVAL_3208 = _EVAL_2046 & _EVAL_2909;
  assign _EVAL_1195 = _EVAL_612 != 2'h0;
  assign _EVAL_1550 = _EVAL_2743[276];
  assign _EVAL_1065 = _EVAL_2941 & _EVAL_1856;
  assign _EVAL_2561 = _EVAL_3780 & _EVAL_3391;
  assign _EVAL_2657 = _EVAL_1782 & _EVAL_1212;
  assign _EVAL_1879 = _EVAL_2656 & _EVAL_2474;
  assign _EVAL_3640 = _EVAL_1782 & _EVAL_2926;
  assign _EVAL_1511 = _EVAL_2743[413];
  assign _EVAL_1092 = _EVAL_1043 & _EVAL_3391;
  assign _EVAL_457 = _EVAL_1246 & _EVAL_3391;
  assign _EVAL_970 = _EVAL_2667 & _EVAL_2909;
  assign _EVAL_2962 = _EVAL_2827 & _EVAL_1856;
  assign _EVAL_3523 = _EVAL_2117 & _EVAL_1856;
  assign _EVAL_1315 = _EVAL_168 & _EVAL_3673;
  assign _EVAL_1481 = _EVAL_1207 & _EVAL_3673;
  assign _EVAL_1033 = _EVAL_2055 & _EVAL_2909;
  assign _EVAL_2226 = _EVAL_1542 & _EVAL_2474;
  assign _EVAL_2553 = _EVAL_1782 & _EVAL_2345;
  assign _EVAL_1283 = _EVAL_1961 & _EVAL_2909;
  assign _EVAL_2667 = _EVAL_2198 & _EVAL_1856;
  assign _EVAL_107 = _EVAL_1782 & _EVAL_1386;
  assign _EVAL_3575 = _EVAL_1542 & _EVAL_2909;
  assign _EVAL_2622 = _EVAL_2743[406];
  assign _EVAL_166 = _EVAL_2743[428];
  assign _EVAL_297 = _EVAL_2734 & _EVAL_1856;
  assign _EVAL_122 = _EVAL_1961 & _EVAL_3673;
  assign _EVAL_3780 = _EVAL_3016 & _EVAL_1856;
  assign _EVAL_1584 = _EVAL_1529 & _EVAL_3391;
  assign _EVAL_1984 = _EVAL_1782 & _EVAL_1278;
  assign _EVAL_2345 = _EVAL_2743[281];
  assign _EVAL_853 = _EVAL_2981 & _EVAL_2474;
  assign _EVAL_720 = _EVAL_2260 & _EVAL_1856;
  assign _EVAL_3802 = _EVAL_1393 & _EVAL_3670;
  assign _EVAL_2372 = _EVAL_2743[458];
  assign _EVAL_2087 = _EVAL_720 & _EVAL_3673;
  assign _EVAL_3503 = _EVAL_2559 & _EVAL_2474;
  assign _EVAL_1241 = _EVAL_1782 & _EVAL_3679;
  assign _EVAL_3141 = _EVAL_2743[19];
  assign _EVAL_903 = _EVAL_3167 & _EVAL_3391;
  assign _EVAL_2753 = _EVAL_2600 & _EVAL_3391;
  assign _EVAL_2180 = _EVAL_2154 & _EVAL_1856;
  assign _EVAL_1855 = _EVAL_2743[365];
  assign _EVAL_1817 = _EVAL_2180 & _EVAL_2909;
  assign _EVAL_2064 = _EVAL_1782 & _EVAL_1898;
  assign _EVAL_532 = _EVAL_2981 & _EVAL_3391;
  assign _EVAL_764 = _EVAL_2745 & _EVAL_3673;
  assign _EVAL_328 = _EVAL_1782 & _EVAL_188;
  assign _EVAL_1188 = _EVAL_220 & _EVAL_3670;
  assign _EVAL_3018 = _EVAL_1782 & _EVAL_2541;
  assign _EVAL_3256 = _EVAL_3718 & _EVAL_3673;
  assign _EVAL_2404 = _EVAL_575[11:0];
  assign _EVAL_319 = _EVAL_1381 & _EVAL_3673;
  assign _EVAL_1816 = _EVAL_2203 & _EVAL_3673;
  assign _EVAL_2618 = _EVAL_2743[494];
  assign _EVAL_3734 = _EVAL_1623 & _EVAL_1856;
  assign _EVAL_1700 = _EVAL_1197 & _EVAL_1856;
  assign _EVAL_3462 = _EVAL_877 & _EVAL_3391;
  assign _EVAL_3210 = _EVAL_3817 & _EVAL_3673;
  assign _EVAL_1716 = _EVAL_1444 & _EVAL_3670;
  assign _EVAL_1609 = _EVAL_3287 & _EVAL_2474;
  assign _EVAL_1636 = _EVAL_1915 & _EVAL_2909;
  assign _EVAL_929 = _EVAL_1782 & _EVAL_2856;
  assign _EVAL_2521 = _EVAL_2729 & _EVAL_1843;
  assign _EVAL_456 = _EVAL_69 & _EVAL_3673;
  assign _EVAL_1247 = _EVAL_999 & _EVAL_2909;
  assign _EVAL_873 = _EVAL_580 & _EVAL_1856;
  assign _EVAL_627 = _EVAL_2139 & _EVAL_3391;
  assign _EVAL_255 = _EVAL_1782 & _EVAL_962;
  assign _EVAL_3400 = _EVAL_3430 & _EVAL_2474;
  assign _EVAL_2931 = _EVAL_297 & _EVAL_2909;
  assign _EVAL_1586 = _EVAL_3175 & _EVAL_1856;
  assign _EVAL_2621 = _EVAL_1381 & _EVAL_2474;
  assign _EVAL_1627 = _EVAL_2743[415];
  assign _EVAL_3269 = _EVAL_310 & _EVAL_1856;
  assign _EVAL_704 = _EVAL_2743[480];
  assign _EVAL_1766 = _EVAL_1543 & _EVAL_1856;
  assign _EVAL_2430 = _EVAL_3284 & _EVAL_749;
  assign _EVAL_574 = _EVAL_1216 & _EVAL_2909;
  assign _EVAL_3303 = _EVAL_69 & _EVAL_2909;
  assign _EVAL_1122 = _EVAL_1782 & _EVAL_860;
  assign _EVAL_137 = _EVAL_367 & _EVAL_1856;
  assign _EVAL_3180 = _EVAL_2307 & _EVAL_2474;
  assign _EVAL_2580 = _EVAL_1782 & _EVAL_1143;
  assign _EVAL_3149 = _EVAL_2245 & _EVAL_1856;
  assign _EVAL_3488 = _EVAL_2016 & _EVAL_3673;
  assign _EVAL_2625 = _EVAL_3332 & _EVAL_3391;
  assign _EVAL_3553 = _EVAL_2123 & _EVAL_1856;
  assign _EVAL_3041 = _EVAL_3521 & _EVAL_1856;
  assign _EVAL_848 = _EVAL_850 & _EVAL_2909;
  assign _EVAL_396 = _EVAL_2425 & _EVAL_3391;
  assign _EVAL_925 = _EVAL_2743[339];
  assign _EVAL_2109 = _EVAL_2431 & _EVAL_3673;
  assign _EVAL_2510 = _EVAL_2551 & _EVAL_3673;
  assign _EVAL_3449 = _EVAL_1782 & _EVAL_524;
  assign _EVAL_302 = _EVAL_3817 & _EVAL_3391;
  assign _EVAL_3570 = _EVAL_977 & _EVAL_2909;
  assign _EVAL_2859 = _EVAL_2055 & _EVAL_3673;
  assign _EVAL_3601 = _EVAL_1100 & _EVAL_772;
  assign _EVAL_1966 = _EVAL_1782 & _EVAL_1850;
  assign _EVAL_3131 = _EVAL_2935 & _EVAL_3673;
  assign _EVAL_1605 = _EVAL_1743 & _EVAL_3673;
  assign _EVAL_3828 = _EVAL_2424 & _EVAL_3391;
  assign _EVAL_1637 = _EVAL_2743[420];
  assign _EVAL_2502 = _EVAL_2666 & _EVAL_3673;
  assign _EVAL_2135 = _EVAL_1782 & _EVAL_427;
  assign _EVAL_543 = _EVAL_1782 & _EVAL_1550;
  assign _EVAL_1862 = _EVAL_3151 & _EVAL_3673;
  assign _EVAL_668 = _EVAL_2972 & _EVAL_2474;
  assign _EVAL_2548 = _EVAL_1782 & _EVAL_1232;
  assign _EVAL_295 = _EVAL_2743[13];
  assign _EVAL_3786 = _EVAL_1782 & _EVAL_750;
  assign _EVAL_896 = _EVAL_3080 & _EVAL_3673;
  assign _EVAL_2212 = _EVAL_1100 & _EVAL_3681;
  assign _EVAL_3392 = _EVAL_1452 & _EVAL_2474;
  assign _EVAL_358 = _EVAL_2729 & _EVAL_1317;
  assign _EVAL_1619 = _EVAL_3638 & _EVAL_3391;
  assign _EVAL_1554 = _EVAL_2551 & _EVAL_2909;
  assign _EVAL_2754 = _EVAL_2675 & _EVAL_3673;
  assign _EVAL_189 = _EVAL_977 & _EVAL_3391;
  assign _EVAL_1172 = _EVAL_961 & _EVAL_1856;
  assign _EVAL_2702 = _EVAL_3261 & _EVAL_2909;
  assign _EVAL_3483 = _EVAL_3232 & _EVAL_3673;
  assign _EVAL_1134 = _EVAL_3527 & _EVAL_3391;
  assign _EVAL_3674 = _EVAL_2364 & _EVAL_1856;
  assign _EVAL_3273 = _EVAL_100 & _EVAL_2474;
  assign _EVAL_210 = _EVAL_2037 & _EVAL_2909;
  assign _EVAL_1411 = _EVAL_2743[417];
  assign _EVAL_782 = _EVAL_3114 & _EVAL_2474;
  assign _EVAL_1479 = _EVAL_3425 | _EVAL_1164;
  assign _EVAL_1535 = _EVAL_2787 & _EVAL_3673;
  assign _EVAL_490 = _EVAL_712 & _EVAL_3673;
  assign _EVAL_733 = _EVAL_173 & _EVAL_3673;
  assign _EVAL_749 = ~_EVAL_1681;
  assign _EVAL_631 = _EVAL_2307 & _EVAL_2909;
  assign _EVAL_3779 = _EVAL_53 & _EVAL_1856;
  assign _EVAL_2377 = _EVAL_2936 & _EVAL_3673;
  assign _EVAL_816 = _EVAL_2649 & _EVAL_2909;
  assign _EVAL_3197 = _EVAL_1766 & _EVAL_2909;
  assign _EVAL_3564 = _EVAL_83[10];
  assign _EVAL_1120 = _EVAL_1246 & _EVAL_2909;
  assign _EVAL_2100 = _EVAL_3055 & _EVAL_3673;
  assign TLMonitor_1__EVAL_6 = {{2'd0}, _EVAL_2004};
  assign _EVAL_3057 = _EVAL_2180 & _EVAL_3673;
  assign _EVAL_1696 = _EVAL_1782 & _EVAL_3054;
  assign _EVAL_3638 = _EVAL_1520 & _EVAL_1856;
  assign _EVAL_1024 = _EVAL_780 & _EVAL_2909;
  assign _EVAL_2122 = _EVAL_1782 & _EVAL_1618;
  assign _EVAL_173 = _EVAL_1378 & _EVAL_1856;
  assign _EVAL_3232 = _EVAL_2657 & _EVAL_1856;
  assign _EVAL_1661 = _EVAL_176 & _EVAL_2474;
  assign _EVAL_1001 = _EVAL_1043 & _EVAL_2909;
  assign _EVAL_2454 = _EVAL_1352 & _EVAL_3391;
  assign _EVAL_3382 = _EVAL_1782 & _EVAL_1242;
  assign _EVAL_588 = _EVAL_176 & _EVAL_3391;
  assign _EVAL_856 = _EVAL_780 & _EVAL_2474;
  assign _EVAL_2633 = _EVAL_1782 & _EVAL_925;
  assign _EVAL_904 = _EVAL_1414 & _EVAL_3673;
  assign _EVAL_2539 = _EVAL_2743[402];
  assign _EVAL_1870 = _EVAL_1309 & _EVAL_2909;
  assign _EVAL_1857 = _EVAL_2034 & _EVAL_2909;
  assign _EVAL_1705 = _EVAL_2425 & _EVAL_2909;
  assign _EVAL_3201 = _EVAL_1782 & _EVAL_3267;
  assign _EVAL_1585 = _EVAL_1782 & _EVAL_2388;
  assign _EVAL_495 = _EVAL_2743[300];
  assign _EVAL_1679 = _EVAL_1782 & _EVAL_1075;
  assign _EVAL_3142 = _EVAL_2743[330];
  assign _EVAL_871 = _EVAL_3015 & _EVAL_2474;
  assign _EVAL_140 = _EVAL_157 & _EVAL_1856;
  assign _EVAL_2245 = _EVAL_1782 & _EVAL_1831;
  assign _EVAL_1259 = _EVAL_712 & _EVAL_2474;
  assign _EVAL_801 = _EVAL_2743[323];
  assign _EVAL_3033 = _EVAL_2743[14];
  assign _EVAL_2644 = _EVAL_3370 & _EVAL_3673;
  assign _EVAL_594 = _EVAL_2425 & _EVAL_3673;
  assign _EVAL_2322 = _EVAL_2743[507];
  assign _EVAL_3222 = _EVAL_1264 & _EVAL_3673;
  assign _EVAL_2637 = _EVAL_1782 & _EVAL_3424;
  assign _EVAL_1424 = _EVAL_1782 & _EVAL_3150;
  assign _EVAL_3352 = _EVAL_999 & _EVAL_3391;
  assign _EVAL_380 = _EVAL_2936 & _EVAL_2474;
  assign _EVAL_2228 = _EVAL_1391 & _EVAL_2909;
  assign _EVAL_2760 = _EVAL_1782 & _EVAL_2270;
  assign _EVAL_246 = _EVAL_1782 & _EVAL_2310;
  assign _EVAL_2013 = _EVAL_3040 & _EVAL_3673;
  assign _EVAL_2912 = _EVAL_1782 & _EVAL_823;
  assign _EVAL_2693 = _EVAL_3317 & _EVAL_1856;
  assign _EVAL_1289 = _EVAL_2922 & _EVAL_3391;
  assign _EVAL_880 = _EVAL_2718 & _EVAL_3673;
  assign _EVAL_1877 = _EVAL_74 & _EVAL_3673;
  assign _EVAL_1409 = _EVAL_1439 & _EVAL_3391;
  assign _EVAL_2670 = _EVAL_1657 & _EVAL_2909;
  assign _EVAL_528 = _EVAL_3216 & _EVAL_2474;
  assign _EVAL_2599 = _EVAL_3399 & _EVAL_3673;
  assign _EVAL_992 = _EVAL_1782 & _EVAL_2027;
  assign _EVAL_2950 = _EVAL_2282 & _EVAL_2909;
  assign _EVAL_3578 = _EVAL_3216 & _EVAL_3673;
  assign _EVAL_3267 = _EVAL_2743[314];
  assign _EVAL_2034 = _EVAL_2852 & _EVAL_1856;
  assign _EVAL_330 = _EVAL_89 & _EVAL_3391;
  assign _EVAL_1162 = _EVAL_878 & _EVAL_3673;
  assign _EVAL_1500 = _EVAL_1782 & _EVAL_2372;
  assign _EVAL_913 = _EVAL_2743[303];
  assign _EVAL_852 = _EVAL_445 & _EVAL_2474;
  assign _EVAL_1305 = _EVAL_2743[331];
  assign _EVAL_2202 = _EVAL_1782 & _EVAL_3376;
  assign _EVAL_299 = _EVAL_2316 & _EVAL_3391;
  assign _EVAL_944 = _EVAL_2745 & _EVAL_3391;
  assign _EVAL_670 = _EVAL_2743[269];
  assign _EVAL_1489 = _EVAL_535 & _EVAL_2474;
  assign _EVAL_1920 = _EVAL_1301 & _EVAL_3673;
  assign _EVAL_1431 = _EVAL_43 & _EVAL_2909;
  assign _EVAL_1434 = _EVAL_2019 & _EVAL_3673;
  assign _EVAL_746 = _EVAL_2743[484];
  assign _EVAL_496 = _EVAL_1782 & _EVAL_828;
  assign _EVAL_2718 = _EVAL_980 & _EVAL_1856;
  assign _EVAL_3758 = _EVAL_1782 & _EVAL_2492;
  assign _EVAL_621 = _EVAL_2918 & _EVAL_2474;
  assign _EVAL_1485 = _EVAL_3245 & _EVAL_2909;
  assign _EVAL_1260 = _EVAL_2424 & _EVAL_2474;
  assign _EVAL_2839 = _EVAL_2743[348];
  assign _EVAL_1645 = _EVAL_355 & _EVAL_3673;
  assign _EVAL_1794 = _EVAL_301 & _EVAL_1856;
  assign _EVAL_625 = _EVAL_3149 & _EVAL_2474;
  assign _EVAL_937 = _EVAL_3780 & _EVAL_3673;
  assign _EVAL_3286 = _EVAL_2139 & _EVAL_2474;
  assign _EVAL_2300 = _EVAL_2743[352];
  assign _EVAL_3037 = _EVAL_2693 & _EVAL_2474;
  assign _EVAL_2906 = _EVAL_2435 & _EVAL_2474;
  assign _EVAL_2782 = _EVAL_287 & _EVAL_2474;
  assign _EVAL_303 = _EVAL_1782 & _EVAL_1626;
  assign _EVAL_321 = _EVAL_2743[393];
  assign _EVAL_1956 = _EVAL_1782 & _EVAL_534;
  assign _EVAL_2132 = _EVAL_623 & _EVAL_3673;
  assign _EVAL_2030 = _EVAL_1043 & _EVAL_3673;
  assign _EVAL_447 = _EVAL_1782 & _EVAL_2498;
  assign _EVAL_1294 = _EVAL_553 & _EVAL_1856;
  assign _EVAL_1164 = ~_EVAL_2400;
  assign _EVAL_2946 = _EVAL_3778 & _EVAL_3391;
  assign _EVAL_1266 = _EVAL_3802 & _EVAL_2474;
  assign _EVAL_1029 = _EVAL_163 & _EVAL_3673;
  assign _EVAL_2148 = _EVAL_314 & _EVAL_3391;
  assign _EVAL_1281 = _EVAL_173 & _EVAL_2474;
  assign _EVAL_250 = _EVAL_60 & _EVAL_1856;
  assign _EVAL_1263 = _EVAL_2799 & _EVAL_2909;
  assign TLMonitor_1__EVAL_0 = _EVAL_20;
  assign _EVAL_2748 = _EVAL_2743[305];
  assign _EVAL_1652 = _EVAL_1715 & _EVAL_2909;
  assign _EVAL_2153 = _EVAL_740 & _EVAL_3673;
  assign _EVAL_3643 = _EVAL_3261 & _EVAL_2474;
  assign _EVAL_3330 = _EVAL_3592 & _EVAL_2909;
  assign _EVAL_483 = _EVAL_2421 & _EVAL_3391;
  assign _EVAL_1521 = _EVAL_2729 & _EVAL_1430;
  assign _EVAL_1712 = _EVAL_3358 & _EVAL_2909;
  assign _EVAL_2069 = _EVAL_1498 & _EVAL_2909;
  assign _EVAL_2949 = _EVAL_2743[466];
  assign _EVAL_3355 = _EVAL_684 & _EVAL_2909;
  assign _EVAL_2329 = _EVAL_2768 & _EVAL_2909;
  assign _EVAL_3351 = _EVAL_3640 & _EVAL_1856;
  assign _EVAL_3218 = _EVAL_3780 & _EVAL_2474;
  assign _EVAL_2649 = _EVAL_1428 & _EVAL_1856;
  assign _EVAL_281 = _EVAL_1006 & _EVAL_3391;
  assign _EVAL_2664 = _EVAL_2743[462];
  assign _EVAL_2331 = _EVAL_2253 & _EVAL_3673;
  assign _EVAL_2281 = _EVAL_818 & _EVAL_2474;
  assign _EVAL_3705 = _EVAL_1322 & _EVAL_2474;
  assign _EVAL_3798 = _EVAL_2743[326];
  assign _EVAL_2897 = _EVAL_3494 & _EVAL_3673;
  assign _EVAL_2000 = _EVAL_173 & _EVAL_3391;
  assign _EVAL_120 = _EVAL_575 != 32'h0;
  assign _EVAL_286 = _EVAL_1440 & _EVAL_1856;
  assign _EVAL_3835 = _EVAL_1533 & _EVAL_1856;
  assign _EVAL_1501 = _EVAL_2787 & _EVAL_2909;
  assign _EVAL_2666 = _EVAL_2058 & _EVAL_1856;
  assign _EVAL_2940 = _EVAL_548 & _EVAL_3673;
  assign _EVAL_2541 = _EVAL_2743[385];
  assign _EVAL_2292 = _EVAL_1503 & _EVAL_2909;
  assign _EVAL_2943 = _EVAL_1961 & _EVAL_3391;
  assign _EVAL_525 = _EVAL_414 & _EVAL_2909;
  assign _EVAL_260 = _EVAL_2431 & _EVAL_3391;
  assign _EVAL_550 = _EVAL_2468 & _EVAL_1856;
  assign _EVAL_2240 = _EVAL_1782 & _EVAL_430;
  assign _EVAL_978 = _EVAL_3620 & _EVAL_3673;
  assign _EVAL_2093 = _EVAL_2022 & _EVAL_1856;
  assign _EVAL_643 = _EVAL_1340 & _EVAL_3673;
  assign _EVAL_1898 = _EVAL_2743[431];
  assign _EVAL_1536 = _EVAL_2743[321];
  assign _EVAL_1890 = _EVAL_2743[307];
  assign _EVAL_211 = _EVAL_1503 & _EVAL_3673;
  assign _EVAL_3274 = _EVAL_2693 & _EVAL_2909;
  assign _EVAL_843 = _EVAL_2236 & _EVAL_3391;
  assign _EVAL_2607 = _EVAL_414 & _EVAL_3673;
  assign _EVAL_472 = _EVAL_780 & _EVAL_3673;
  assign _EVAL_475 = _EVAL_274 & _EVAL_3391;
  assign _EVAL_534 = _EVAL_2743[0];
  assign _EVAL_3749 = _EVAL_678 & _EVAL_3673;
  assign _EVAL_2297 = _EVAL_2981 & _EVAL_2909;
  assign _EVAL_701 = _EVAL_2055 & _EVAL_3391;
  assign _EVAL_2303 = _EVAL_3120 & _EVAL_3670;
  assign _EVAL_2386 = _EVAL_667 & _EVAL_2909;
  assign _EVAL_927 = _EVAL_2028 & _EVAL_2474;
  assign _EVAL_2681 = _EVAL_1299 & _EVAL_2909;
  assign _EVAL_1715 = _EVAL_1648 & _EVAL_1856;
  assign _EVAL_1630 = _EVAL_1782 & _EVAL_2710;
  assign _EVAL_3617 = _EVAL_1783 & _EVAL_2909;
  assign _EVAL_3757 = _EVAL_1967 & _EVAL_1995;
  assign _EVAL_75 = _EVAL_1782 & _EVAL_2448;
  assign _EVAL_1063 = _EVAL_3347 & _EVAL_3673;
  assign _EVAL_894 = _EVAL_2282 & _EVAL_2474;
  assign _EVAL_3112 = _EVAL_2743[259];
  assign _EVAL_388 = _EVAL_2849 & _EVAL_2474;
  assign _EVAL_579 = _EVAL_1782 & _EVAL_161;
  assign _EVAL_2337 = _EVAL_1964 & _EVAL_2909;
  assign _EVAL_3538 = _EVAL_3803 & _EVAL_2909;
  assign _EVAL_3117 = _EVAL_1715 & _EVAL_3391;
  assign _EVAL_3565 = _EVAL_3261 & _EVAL_3673;
  assign _EVAL_818 = _EVAL_1667 & _EVAL_1856;
  assign _EVAL_2407 = _EVAL_2743[390];
  assign _EVAL_278 = _EVAL_168 & _EVAL_3391;
  assign _EVAL_1551 = _EVAL_1782 & _EVAL_411;
  assign _EVAL_3631 = _EVAL_3821 & _EVAL_2909;
  assign _EVAL_1440 = _EVAL_1782 & _EVAL_2944;
  assign _EVAL_864 = _EVAL_3285 & _EVAL_3391;
  assign _EVAL_267 = _EVAL_2817 & _EVAL_2474;
  assign _EVAL_2910 = _EVAL_107 & _EVAL_1856;
  assign _EVAL_2954 = _EVAL_1782 & _EVAL_476;
  assign _EVAL_2876 = _EVAL_1986 & _EVAL_3673;
  assign _EVAL_408 = _EVAL_3778 & _EVAL_2474;
  assign _EVAL_1032 = _EVAL_1479 | _EVAL_470;
  assign _EVAL_452 = _EVAL_2910 & _EVAL_2909;
  assign _EVAL_3619 = _EVAL_2743[505];
  assign _EVAL_3573 = _EVAL_1782 & _EVAL_3820;
  assign _EVAL_2966 = _EVAL_1363 & _EVAL_2909;
  assign _EVAL_3362 = _EVAL_1635 & _EVAL_3673;
  assign _EVAL_3344 = _EVAL_1356 & _EVAL_2909;
  assign _EVAL_2632 = _EVAL_2729 & _EVAL_3438;
  assign _EVAL_1537 = _EVAL_2435 & _EVAL_2909;
  assign _EVAL_3803 = _EVAL_3373 & _EVAL_1856;
  assign _EVAL_1750 = _EVAL_1356 & _EVAL_3391;
  assign _EVAL_1022 = _EVAL_1782 & _EVAL_1714;
  assign _EVAL_2346 = _EVAL_1301 & _EVAL_2474;
  assign _EVAL_637 = _EVAL_2743[456];
  assign _EVAL_2152 = _EVAL_1094 & _EVAL_2909;
  assign _EVAL_2614 = _EVAL_2743[491];
  assign _EVAL_1058 = _EVAL_445 & _EVAL_3391;
  assign _EVAL_780 = _EVAL_142 & _EVAL_1856;
  assign _EVAL_2082 = _EVAL_2161 & _EVAL_2909;
  assign _EVAL_889 = _EVAL_3466 & _EVAL_3391;
  assign _EVAL_1762 = _EVAL_1715 & _EVAL_3673;
  assign _EVAL_2172 = _EVAL_3835 & _EVAL_3391;
  assign _EVAL_2349 = _EVAL_1782 & _EVAL_101;
  assign _EVAL_3048 = _EVAL_2743[495];
  assign _EVAL_1800 = _EVAL_1294 & _EVAL_2909;
  assign _EVAL_2269 = _EVAL_550 & _EVAL_3391;
  assign _EVAL_800 = _EVAL_3229 & _EVAL_3673;
  assign _EVAL_1048 = _EVAL_2743[412];
  assign _EVAL_845 = _EVAL_3332 & _EVAL_2474;
  assign _EVAL_742 = _EVAL_2799 & _EVAL_3391;
  assign _EVAL_899 = _EVAL_2303 & _EVAL_3673;
  assign _EVAL_1443 = _EVAL_3532 & _EVAL_2474;
  assign _EVAL_2534 = _EVAL_1782 & _EVAL_914;
  assign _EVAL_3579 = _EVAL_2743[391];
  assign _EVAL_3812 = _EVAL_1091 & _EVAL_1856;
  assign _EVAL_1208 = _EVAL_1782 & _EVAL_3512;
  assign _EVAL_1454 = _EVAL_1782 & _EVAL_1917;
  assign _EVAL_1919 = _EVAL_2999 != 4'h0;
  assign _EVAL_1144 = _EVAL_1329 & _EVAL_2909;
  assign _EVAL_1964 = _EVAL_604 & _EVAL_1856;
  assign _EVAL_3375 = _EVAL_2554 & _EVAL_2474;
  assign _EVAL_1621 = _EVAL_3285 & _EVAL_2909;
  assign _EVAL_1901 = _EVAL_779 & _EVAL_2474;
  assign _EVAL_2904 = _EVAL_355 & _EVAL_2474;
  assign _EVAL_917 = _EVAL_3040 & _EVAL_2474;
  assign _EVAL_3729 = _EVAL_2743[257];
  assign _EVAL_2518 = _EVAL_2229 & _EVAL_3391;
  assign _EVAL_2550 = _EVAL_2743[7];
  assign _EVAL_672 = _EVAL_2229 & _EVAL_2474;
  assign _EVAL_1384 = _EVAL_1782 & _EVAL_190;
  assign _EVAL_2991 = _EVAL_1782 & _EVAL_2722;
  assign _EVAL_2646 = _EVAL_740 & _EVAL_2474;
  assign _EVAL_518 = _EVAL_1782 & _EVAL_2475;
  assign _EVAL_247 = _EVAL_1452 & _EVAL_2909;
  assign _EVAL_633 = _EVAL_3608 & _EVAL_3391;
  assign _EVAL_2155 = _EVAL_652 & _EVAL_3673;
  assign _EVAL_1233 = _EVAL_3587 & _EVAL_2909;
  assign _EVAL_2764 = _EVAL_3229 & _EVAL_2909;
  assign _EVAL_576 = _EVAL_579 & _EVAL_1856;
  assign _EVAL_1974 = _EVAL_2743[366];
  assign _EVAL_2123 = _EVAL_1782 & _EVAL_657;
  assign _EVAL_359 = _EVAL_1327 & _EVAL_3673;
  assign _EVAL_2266 = _EVAL_3287 & _EVAL_2909;
  assign _EVAL_821 = _EVAL_1782 & _EVAL_1078;
  assign _EVAL_874 = _EVAL_2037 & _EVAL_2474;
  assign _EVAL_2179 = _EVAL_3368 & _EVAL_3391;
  assign _EVAL_3213 = _EVAL_1782 & _EVAL_1840;
  assign _EVAL_813 = _EVAL_3523 & _EVAL_3673;
  assign _EVAL_3479 = _EVAL_455 & _EVAL_2474;
  assign _EVAL_3079 = _EVAL_2743[282];
  assign _EVAL_3365 = _EVAL_3786 & _EVAL_1856;
  assign _EVAL_197 = _EVAL_1766 & _EVAL_3673;
  assign _EVAL_3272 = _EVAL_2743[405];
  assign _EVAL_887 = _EVAL_511 & _EVAL_2474;
  assign _EVAL_1943 = _EVAL_740 & _EVAL_3391;
  assign _EVAL_3440 = _EVAL_3466 & _EVAL_3673;
  assign _EVAL_3245 = _EVAL_1966 & _EVAL_3670;
  assign _EVAL_2669 = _EVAL_979 & _EVAL_3639;
  assign _EVAL_2270 = _EVAL_2743[317];
  assign _EVAL_2124 = _EVAL_1782 & _EVAL_2296;
  assign _EVAL_157 = _EVAL_1782 & _EVAL_2925;
  assign _EVAL_1784 = _EVAL_2613 & _EVAL_3391;
  assign _EVAL_750 = _EVAL_2743[358];
  assign _EVAL_1250 = _EVAL_2743[454];
  assign _EVAL_1748 = _EVAL_1782 & _EVAL_2276;
  assign _EVAL_1949 = _EVAL_2068 & _EVAL_2474;
  assign TLMonitor__EVAL_2 = _EVAL_38;
  assign _EVAL_3622 = _EVAL_2203 & _EVAL_2474;
  assign _EVAL_262 = _EVAL_1782 & _EVAL_1627;
  assign _EVAL_218 = _EVAL_305 & _EVAL_3391;
  assign _EVAL_3514 = _EVAL_1892 & _EVAL_2474;
  assign _EVAL_1356 = _EVAL_2146 & _EVAL_1856;
  assign _EVAL_1223 = _EVAL_1201 & _EVAL_2909;
  assign _EVAL_1158 = _EVAL_3803 & _EVAL_2474;
  assign _EVAL_1430 = _EVAL_575[9];
  assign _EVAL_3801 = _EVAL_250 & _EVAL_2474;
  assign _EVAL_3406 = _EVAL_26[9:0];
  assign _EVAL_2446 = _EVAL_2271 & _EVAL_3673;
  assign _EVAL_629 = _EVAL_3532 & _EVAL_2909;
  assign _EVAL_2442 = _EVAL_2743[11];
  assign _EVAL_3358 = _EVAL_413 & _EVAL_1856;
  assign _EVAL_2787 = _EVAL_3226 & _EVAL_1856;
  assign _EVAL_1788 = _EVAL_1782 & _EVAL_503;
  assign _EVAL_114 = _EVAL_1782 & _EVAL_2197;
  assign _EVAL_2289 = _EVAL_3674 & _EVAL_3391;
  assign _EVAL_2011 = _EVAL_1542 & _EVAL_3673;
  assign _EVAL_1442 = _EVAL_1282 & _EVAL_3673;
  assign _EVAL_1852 = _EVAL_576 & _EVAL_3391;
  assign _EVAL_828 = _EVAL_2743[488];
  assign _EVAL_1355 = _EVAL_2743[356];
  assign _EVAL_3376 = _EVAL_2743[377];
  assign _EVAL_1416 = _EVAL_2016 & _EVAL_2909;
  assign _EVAL_1272 = _EVAL_690 & _EVAL_1856;
  assign _EVAL_830 = _EVAL_1938 & _EVAL_2909;
  assign _EVAL_1520 = _EVAL_1782 & _EVAL_3477;
  assign _EVAL_3831 = _EVAL_2743[395];
  assign _EVAL_3819 = _EVAL_2043 & _EVAL_3391;
  assign _EVAL_3301 = _EVAL_999 & _EVAL_3673;
  assign _EVAL_635 = _EVAL_3080 & _EVAL_2909;
  assign _EVAL_814 = _EVAL_1743 & _EVAL_2909;
  assign _EVAL_644 = _EVAL_3357 & _EVAL_2909;
  assign _EVAL_2577 = _EVAL_2435 & _EVAL_3673;
  assign _EVAL_300 = _EVAL_2656 & _EVAL_2909;
  assign _EVAL_3718 = _EVAL_371 & _EVAL_1856;
  assign _EVAL_1533 = _EVAL_1782 & _EVAL_560;
  assign _EVAL_1293 = _EVAL_1793 & _EVAL_3391;
  assign _EVAL_1608 = _EVAL_3597 & _EVAL_2474;
  assign _EVAL_3162 = _EVAL_2743[380];
  assign _EVAL_371 = _EVAL_1782 & _EVAL_2048;
  assign _EVAL_3721 = _EVAL_398 & _EVAL_3391;
  assign _EVAL_1915 = _EVAL_2980 & _EVAL_1856;
  assign _EVAL_2941 = _EVAL_1782 & _EVAL_1642;
  assign _EVAL_1505 = _EVAL_3114 & _EVAL_3673;
  assign _EVAL_3040 = _EVAL_1702 & _EVAL_1856;
  assign _EVAL_3118 = _EVAL_2743[467];
  assign _EVAL_3562 = _EVAL_1782 & _EVAL_704;
  assign _EVAL_46 = _EVAL_2743[373];
  assign _EVAL_1837 = _EVAL_1782 & _EVAL_2634;
  assign _EVAL_850 = _EVAL_134 & _EVAL_1856;
  assign _EVAL_2310 = _EVAL_2743[334];
  assign _EVAL_2062 = _EVAL_2675 & _EVAL_3391;
  assign _EVAL_3516 = _EVAL_3760 & _EVAL_3391;
  assign _EVAL_47 = _EVAL_2743[423];
  assign _EVAL_310 = _EVAL_1782 & _EVAL_888;
  assign _EVAL_3381 = _EVAL_873 & _EVAL_2474;
  assign _EVAL_1265 = _EVAL_3534 & _EVAL_3673;
  assign _EVAL_1284 = _EVAL_2667 & _EVAL_3391;
  assign _EVAL_2975 = _EVAL_3779 & _EVAL_2474;
  assign _EVAL_1452 = _EVAL_1384 & _EVAL_1856;
  assign _EVAL_1189 = _EVAL_2772 & _EVAL_3670;
  assign _EVAL_2772 = _EVAL_1782 & _EVAL_1727;
  assign _EVAL_1278 = _EVAL_2743[481];
  assign _EVAL_2860 = _EVAL_1065 & _EVAL_2474;
  assign _EVAL_3410 = _EVAL_2743[476];
  assign _EVAL_2543 = _EVAL_1189 & _EVAL_2909;
  assign _EVAL_48 = _EVAL_1064 & _EVAL_2909;
  assign _EVAL_803 = _EVAL_1165 & _EVAL_3673;
  assign _EVAL_3437 = _EVAL_1782 & _EVAL_2748;
  assign _EVAL_1484 = _EVAL_1782 & _EVAL_2960;
  assign _EVAL_665 = _EVAL_2134 & _EVAL_2909;
  assign _EVAL_3407 = _EVAL_1381 & _EVAL_2909;
  assign _EVAL_1449 = _EVAL_1782 & _EVAL_2490;
  assign _EVAL_3546 = _EVAL_3544 & _EVAL_2909;
  assign _EVAL_2645 = _EVAL_2229 & _EVAL_2909;
  assign _EVAL_2045 = _EVAL_2743[349];
  assign _EVAL_3300 = _EVAL_2165 & _EVAL_2909;
  assign _EVAL_2483 = _EVAL_1793 & _EVAL_2909;
  assign _EVAL_1951 = _EVAL_3394 & _EVAL_1856;
  assign _EVAL_3441 = _EVAL_3327 & _EVAL_3673;
  assign _EVAL_1574 = _EVAL_1782 & _EVAL_1250;
  assign _EVAL_1749 = _EVAL_596 & _EVAL_3673;
  assign _EVAL_337 = _EVAL_1782 & _EVAL_2949;
  assign _EVAL_2926 = _EVAL_2743[368];
  assign _EVAL_1765 = _EVAL_246 & _EVAL_1856;
  assign _EVAL_283 = _EVAL_720 & _EVAL_3391;
  assign _EVAL_1689 = _EVAL_2743[452];
  assign _EVAL_648 = _EVAL_3040 & _EVAL_2909;
  assign _EVAL_1205 = _EVAL_2743[438];
  assign _EVAL_2206 = _EVAL_2202 & _EVAL_1856;
  assign _EVAL_2728 = _EVAL_1740 & _EVAL_2474;
  assign _EVAL_1504 = _EVAL_2253 & _EVAL_2909;
  assign _EVAL_3285 = _EVAL_3562 & _EVAL_1856;
  assign _EVAL_2738 = _EVAL_708 & _EVAL_1856;
  assign _EVAL_1730 = ~_EVAL_885;
  assign _EVAL_1473 = _EVAL_1439 & _EVAL_2474;
  assign _EVAL_2900 = _EVAL_2093 & _EVAL_3673;
  assign _EVAL_3559 = _EVAL_168 & _EVAL_2909;
  assign _EVAL_342 = _EVAL_2880 & _EVAL_3673;
  assign _EVAL_400 = _EVAL_1657 & _EVAL_3391;
  assign _EVAL_1809 = _EVAL_1973 & _EVAL_3673;
  assign _EVAL_3792 = _EVAL_1309 & _EVAL_3673;
  assign _EVAL_2766 = _EVAL_1743 & _EVAL_3391;
  assign _EVAL_966 = _EVAL_1782 & _EVAL_224;
  assign _EVAL_3708 = _EVAL_355 & _EVAL_3391;
  assign _EVAL_2197 = _EVAL_2743[285];
  assign _EVAL_761 = _EVAL_3269 & _EVAL_897;
  assign _EVAL_1141 = _EVAL_376 & _EVAL_3391;
  assign _EVAL_2084 = _EVAL_2553 & _EVAL_1856;
  assign _EVAL_2450 = _EVAL_3332 & _EVAL_3673;
  assign _EVAL_2564 = _EVAL_1414 & _EVAL_3391;
  assign _EVAL_2271 = _EVAL_2231 & _EVAL_3670;
  assign _EVAL_2694 = _EVAL_1782 & _EVAL_3112;
  assign _EVAL_3489 = _EVAL_2161 & _EVAL_2474;
  assign _EVAL_2033 = _EVAL_2743[308];
  assign _EVAL_3373 = _EVAL_1782 & _EVAL_1053;
  assign _EVAL_1922 = ~_EVAL_38;
  assign _EVAL_3833 = _EVAL_286 & _EVAL_2909;
  assign _EVAL_2562 = _EVAL_2525 & _EVAL_2474;
  assign _EVAL_640 = _EVAL_2338 & _EVAL_2474;
  assign _EVAL_2287 = _EVAL_3167 & _EVAL_2909;
  assign _EVAL_68 = _EVAL_1327 & _EVAL_2474;
  assign TLMonitor__EVAL_4 = _EVAL_2;
  assign _EVAL_618 = _EVAL_1782 & _EVAL_2127;
  assign _EVAL_791 = _EVAL_2666 & _EVAL_2909;
  assign _EVAL_1796 = _EVAL_610 & _EVAL_2909;
  assign _EVAL_3278 = _EVAL_548 & _EVAL_2909;
  assign _EVAL_3678 = _EVAL_1782 & _EVAL_3133;
  assign _EVAL_2597 = _EVAL_2743[490];
  assign _EVAL_2182 = _EVAL_2206 & _EVAL_2474;
  assign _EVAL_1451 = _EVAL_3151 & _EVAL_2474;
  assign _EVAL_69 = _EVAL_3396 & _EVAL_1856;
  assign _EVAL_135 = _EVAL_740 & _EVAL_2909;
  assign _EVAL_3760 = _EVAL_1574 & _EVAL_1856;
  assign _EVAL_3787 = _EVAL_1782 & _EVAL_2449;
  assign _EVAL_3810 = _EVAL_2743[332];
  assign _EVAL_1336 = _EVAL_414 & _EVAL_3391;
  assign _EVAL_1492 = _EVAL_1094 & _EVAL_3673;
  assign _EVAL_2557 = _EVAL_1405 & _EVAL_2474;
  assign _EVAL_2802 = _EVAL_2743[320];
  assign _EVAL_3805 = _EVAL_2918 & _EVAL_3391;
  assign _EVAL_2396 = _EVAL_2933 & _EVAL_1856;
  assign _EVAL_3363 = _EVAL_286 & _EVAL_3673;
  assign _EVAL_350 = _EVAL_2743[347];
  assign _EVAL_183 = _EVAL_2396 & _EVAL_2909;
  assign _EVAL_3124 = _EVAL_1782 & _EVAL_2407;
  assign _EVAL_2914 = _EVAL_2019 & _EVAL_2909;
  assign _EVAL_998 = _EVAL_1241 & _EVAL_1856;
  assign _EVAL_2516 = _EVAL_414 & _EVAL_2474;
  assign _EVAL_1814 = _EVAL_288 & _EVAL_2909;
  assign _EVAL_1655 = _EVAL_1782 & _EVAL_2597;
  assign _EVAL_823 = _EVAL_2743[17];
  assign _EVAL_3074 = _EVAL_3779 & _EVAL_2909;
  assign _EVAL_1192 = _EVAL_2428 & _EVAL_2909;
  assign _EVAL_1482 = _EVAL_3229 & _EVAL_3391;
  assign _EVAL_1651 = _EVAL_3645 & _EVAL_3673;
  assign _EVAL_2773 = _EVAL_779 & _EVAL_3673;
  assign _EVAL_2119 = _EVAL_3091 & _EVAL_1856;
  assign _EVAL_476 = _EVAL_2743[266];
  assign _EVAL_2184 = _EVAL_1794 & _EVAL_2474;
  assign _EVAL_3533 = _EVAL_1782 & _EVAL_1193;
  assign _EVAL_994 = _EVAL_2743[447];
  assign _EVAL_3785 = _EVAL_1352 & _EVAL_3673;
  assign _EVAL_2884 = _EVAL_3151 & _EVAL_3391;
  assign _EVAL_1102 = _EVAL_618 & _EVAL_1856;
  assign _EVAL_2032 = _EVAL_3534 & _EVAL_3391;
  assign _EVAL_981 = _EVAL_2935 & _EVAL_3391;
  assign _EVAL_338 = _EVAL_287 & _EVAL_3673;
  assign _EVAL_2660 = _EVAL_1782 & _EVAL_3224;
  assign _EVAL_717 = _EVAL_1708 & _EVAL_1856;
  assign _EVAL_732 = _EVAL_2743[499];
  assign _EVAL_2321 = _EVAL_3779 & _EVAL_3673;
  assign _EVAL_2200 = _EVAL_2428 & _EVAL_3391;
  assign _EVAL_1190 = _EVAL_3167 & _EVAL_3673;
  assign _EVAL_1565 = _EVAL_137 & _EVAL_2474;
  assign _EVAL_494 = _EVAL_535 & _EVAL_3391;
  assign _EVAL_2609 = _EVAL_1782 & _EVAL_3822;
  assign _EVAL_3120 = _EVAL_1782 & _EVAL_1404;
  assign _EVAL_2776 = _EVAL_2282 & _EVAL_3391;
  assign _EVAL_806 = _EVAL_176 & _EVAL_3673;
  assign _EVAL_460 = _EVAL_3015 & _EVAL_2909;
  assign _EVAL_307 = _EVAL_575[19:17];
  assign _EVAL_3840 = _EVAL_1782 & _EVAL_1760;
  assign _EVAL_2866 = _EVAL_1973 & _EVAL_2474;
  assign _EVAL_2952 = _EVAL_1782 & _EVAL_3170;
  assign _EVAL_878 = _EVAL_2701 & _EVAL_1856;
  assign _EVAL_767 = _EVAL_3232 & _EVAL_2474;
  assign _EVAL_2416 = _EVAL_2729 & _EVAL_145;
  assign _EVAL_1393 = _EVAL_1782 & _EVAL_2442;
  assign _EVAL_524 = _EVAL_2743[418];
  assign _EVAL_418 = _EVAL_1782 & _EVAL_3432;
  assign _EVAL_445 = _EVAL_303 & _EVAL_1856;
  assign _EVAL_2919 = _EVAL_610 & _EVAL_3673;
  assign _EVAL_1171 = _EVAL_2998 & _EVAL_3673;
  assign _EVAL_2852 = _EVAL_1782 & _EVAL_390;
  assign _EVAL_276 = _EVAL_1282 & _EVAL_2909;
  assign _EVAL_1722 = _EVAL_1782 & _EVAL_3453;
  assign _EVAL_74 = _EVAL_2025 & _EVAL_1856;
  assign _EVAL_682 = _EVAL_3371 & _EVAL_1856;
  assign _EVAL_3827 = _EVAL_3149 & _EVAL_3673;
  assign _EVAL_1899 = _EVAL_1635 & _EVAL_2909;
  assign _EVAL_3107 = _EVAL_2649 & _EVAL_3391;
  assign _EVAL_584 = _EVAL_2765 & _EVAL_2474;
  assign _EVAL_2587 = _EVAL_1716 & _EVAL_3391;
  assign _EVAL_3317 = _EVAL_1782 & _EVAL_2539;
  assign _EVAL_1292 = _EVAL_2643 & _EVAL_138;
  assign _EVAL_1629 = _EVAL_1782 & _EVAL_671;
  assign _EVAL_1406 = _EVAL_140 & _EVAL_3391;
  assign _EVAL_1002 = _EVAL_3041 & _EVAL_2909;
  assign _EVAL_3467 = _EVAL_2600 & _EVAL_2474;
  assign _EVAL_3042 = _EVAL_2743[388];
  assign _EVAL_222 = _EVAL_3638 & _EVAL_2474;
  assign _EVAL_1674 = _EVAL_1432 & _EVAL_3391;
  assign _EVAL_3341 = _EVAL_726 & _EVAL_2474;
  assign _EVAL_1782 = _EVAL_624 & _EVAL_2004;
  assign _EVAL_364 = _EVAL_1644 & _EVAL_3673;
  assign _EVAL_2795 = _EVAL_1782 & _EVAL_232;
  assign _EVAL_2305 = _EVAL_231 & _EVAL_1856;
  assign _EVAL_1930 = _EVAL_1272 & _EVAL_3391;
  assign _EVAL_1204 = _EVAL_1447 & _EVAL_1856;
  assign _EVAL_3655 = _EVAL_2068 & _EVAL_3673;
  assign _EVAL_2535 = _EVAL_2981 & _EVAL_3673;
  assign _EVAL_3185 = _EVAL_1570 & _EVAL_1856;
  assign _EVAL_231 = _EVAL_1782 & _EVAL_2370;
  assign _EVAL_2567 = _EVAL_726 & _EVAL_3673;
  assign _EVAL_491 = _EVAL_507 & _EVAL_3673;
  assign _EVAL_2813 = _EVAL_1272 & _EVAL_2909;
  assign _EVAL_2250 = _EVAL_2787 & _EVAL_2474;
  assign _EVAL_322 = _EVAL_1551 & _EVAL_1856;
  assign _EVAL_2848 = _EVAL_1782 & _EVAL_2322;
  assign _EVAL_920 = _EVAL_83[11];
  assign _EVAL_676 = _EVAL_2743[15];
  assign _EVAL_570 = _EVAL_235 & _EVAL_2474;
  assign TLMonitor__EVAL_0 = _EVAL_33;
  assign _EVAL_1318 = _EVAL_1782 & _EVAL_1691;
  assign _EVAL_2747 = _EVAL_911 & _EVAL_2909;
  assign _EVAL_1043 = _EVAL_1960 & _EVAL_1856;
  assign _EVAL_1647 = _EVAL_948 & _EVAL_3391;
  assign _EVAL_3261 = _EVAL_1655 & _EVAL_1856;
  assign _EVAL_3063 = _EVAL_298 & _EVAL_2909;
  assign _EVAL_2898 = _EVAL_2478 & _EVAL_2474;
  assign _EVAL_586 = _EVAL_1207 & _EVAL_3391;
  assign _EVAL_1673 = _EVAL_3216 & _EVAL_3391;
  assign _EVAL_2478 = _EVAL_947 & _EVAL_1856;
  assign _EVAL_3477 = _EVAL_2743[399];
  assign _EVAL_116 = _EVAL_1006 & _EVAL_2909;
  assign _EVAL_2126 = _EVAL_1782 & _EVAL_1169;
  assign _EVAL_2805 = _EVAL_1700 & _EVAL_2909;
  assign _EVAL_385 = _EVAL_2068 & _EVAL_3391;
  assign _EVAL_1632 = _EVAL_3638 & _EVAL_2909;
  assign _EVAL_2551 = _EVAL_933 & _EVAL_1856;
  assign _EVAL_1277 = _EVAL_1782 & _EVAL_1205;
  assign _EVAL_1129 = _EVAL_1126 & _EVAL_2474;
  assign _EVAL_3371 = _EVAL_1782 & _EVAL_2118;
  assign _EVAL_2307 = _EVAL_1318 & _EVAL_1856;
  assign _EVAL_544 = _EVAL_712 & _EVAL_2909;
  assign _EVAL_1016 = _EVAL_1782 & _EVAL_1998;
  assign _EVAL_1861 = _EVAL_1782 & _EVAL_2099;
  assign _EVAL_2568 = _EVAL_3740 & _EVAL_1856;
  assign _EVAL_455 = _EVAL_75 & _EVAL_1856;
  assign _EVAL_2037 = _EVAL_1662 & _EVAL_1856;
  assign _EVAL_2444 = _EVAL_1006 & _EVAL_3673;
  assign _EVAL_3419 = _EVAL_2768 & _EVAL_3391;
  assign _EVAL_1340 = _EVAL_3473 & _EVAL_1856;
  assign _EVAL_2019 = _EVAL_656 & _EVAL_1856;
  assign _EVAL_440 = _EVAL_2743[263];
  assign _EVAL_1963 = _EVAL_1782 & _EVAL_758;
  assign _EVAL_3581 = _EVAL_3561 & _EVAL_3673;
  assign _EVAL_623 = _EVAL_578 & _EVAL_1856;
  assign _EVAL_318 = _EVAL_3674 & _EVAL_2474;
  assign _EVAL_429 = _EVAL_667 & _EVAL_3391;
  assign _EVAL_2448 = _EVAL_2743[432];
  assign _EVAL_411 = _EVAL_2743[299];
  assign _EVAL_2875 = _EVAL_3638 & _EVAL_3673;
  assign _EVAL_1025 = _EVAL_646 & _EVAL_3391;
  assign _EVAL_2232 = _EVAL_1586 & _EVAL_3391;
  assign _EVAL_3818 = _EVAL_3365 & _EVAL_3391;
  assign _EVAL_1299 = _EVAL_3382 & _EVAL_1856;
  assign _EVAL_1763 = _EVAL_3287 & _EVAL_3673;
  assign _EVAL_2613 = _EVAL_2439 & _EVAL_1856;
  assign _EVAL_2356 = _EVAL_3041 & _EVAL_3391;
  assign _EVAL_3532 = _EVAL_2795 & _EVAL_1856;
  assign _EVAL_2826 = _EVAL_1782 & _EVAL_1128;
  assign _EVAL_3765 = _EVAL_3645 & _EVAL_2474;
  assign _EVAL_2526 = _EVAL_1782 & _EVAL_1751;
  assign _EVAL_2924 = _EVAL_1766 & _EVAL_3391;
  assign _EVAL_2423 = _EVAL_1782 & _EVAL_1234;
  assign _EVAL_3277 = _EVAL_3630 & _EVAL_2474;
  assign _EVAL_1691 = _EVAL_2743[268];
  assign _EVAL_52 = _EVAL_2165 & _EVAL_3673;
  assign _EVAL_1006 = _EVAL_1277 & _EVAL_1856;
  assign _EVAL_2531 = _EVAL_2134 & _EVAL_3391;
  assign _EVAL_1743 = _EVAL_1703 & _EVAL_1856;
  assign _EVAL_1612 = _EVAL_2693 & _EVAL_3391;
  assign _EVAL_1923 = _EVAL_3817 & _EVAL_2909;
  assign _EVAL_1843 = _EVAL_575[4];
  assign _EVAL_2617 = _EVAL_3114 & _EVAL_2909;
  assign _EVAL_489 = _EVAL_2962 & _EVAL_2474;
  assign _EVAL_144 = _EVAL_2675 & _EVAL_2474;
  assign _EVAL_2171 = _EVAL_2880 & _EVAL_2909;
  assign _EVAL_2439 = _EVAL_1782 & _EVAL_2793;
  assign _EVAL_2431 = _EVAL_3124 & _EVAL_1856;
  assign _EVAL_1156 = _EVAL_3347 & _EVAL_3391;
  assign _EVAL_988 = _EVAL_3690 & _EVAL_1856;
  assign _EVAL_1671 = _EVAL_3778 & _EVAL_2909;
  assign _EVAL_2880 = _EVAL_1566 & _EVAL_1856;
  assign _EVAL_3607 = _EVAL_1100 & _EVAL_128;
  assign _EVAL_148 = _EVAL_1964 & _EVAL_3391;
  assign _EVAL_2192 = _EVAL_3368 & _EVAL_2909;
  assign _EVAL_2401 = _EVAL_3214 & _EVAL_1856;
  assign _EVAL_1072 = _EVAL_507 & _EVAL_3391;
  assign _EVAL_2923 = _EVAL_1452 & _EVAL_3391;
  assign _EVAL_3007 = _EVAL_2922 & _EVAL_2474;
  assign _EVAL_598 = _EVAL_1656 & _EVAL_3673;
  assign _EVAL_2783 = _EVAL_2765 & _EVAL_3391;
  assign _EVAL_128 = _EVAL_2267 != 5'h0;
  assign _EVAL_2389 = _EVAL_2743[416];
  assign _EVAL_773 = _EVAL_596 & _EVAL_2909;
  assign _EVAL_3360 = _EVAL_1837 & _EVAL_1856;
  assign _EVAL_1791 = _EVAL_948 & _EVAL_2909;
  assign _EVAL_758 = _EVAL_2743[453];
  assign _EVAL_536 = _EVAL_1294 & _EVAL_3673;
  assign _EVAL_1602 = _EVAL_1322 & _EVAL_3391;
  assign _EVAL_658 = _EVAL_201 & _EVAL_3673;
  assign _EVAL_2830 = _EVAL_3674 & _EVAL_2909;
  assign _EVAL_2677 = _EVAL_3213 & _EVAL_1856;
  assign _EVAL_1745 = _EVAL_610 & _EVAL_2474;
  assign _EVAL_865 = _EVAL_3760 & _EVAL_2474;
  assign _EVAL_1256 = _EVAL_575[8];
  assign _EVAL_291 = _EVAL_3041 & _EVAL_3673;
  assign _EVAL_1625 = _EVAL_1644 & _EVAL_2474;
  assign _EVAL_862 = _EVAL_1498 & _EVAL_2474;
  assign _EVAL_940 = _EVAL_2165 & _EVAL_2474;
  assign _EVAL_3163 = _EVAL_3630 & _EVAL_2909;
  assign _EVAL_3029 = _EVAL_3645 & _EVAL_3391;
  assign _EVAL_1954 = _EVAL_328 & _EVAL_1856;
  assign _EVAL_1688 = _EVAL_2271 & _EVAL_2909;
  assign _EVAL_1818 = _EVAL_2743[506];
  assign _EVAL_1792 = _EVAL_3630 & _EVAL_3673;
  assign _EVAL_3571 = _EVAL_2743[379];
  assign _EVAL_3204 = _EVAL_1782 & _EVAL_3810;
  assign _EVAL_1146 = _EVAL_1352 & _EVAL_2474;
  assign _EVAL_2740 = _EVAL_2743[496];
  assign _EVAL_1998 = _EVAL_2743[364];
  assign _EVAL_165 = _EVAL_2435 & _EVAL_3391;
  assign _EVAL_2165 = _EVAL_564 & _EVAL_1856;
  assign _EVAL_3307 = _EVAL_3024 & _EVAL_3673;
  assign _EVAL_1017 = _EVAL_1782 & _EVAL_1491;
  assign _EVAL_1626 = _EVAL_2743[327];
  assign _EVAL_196 = _EVAL_1421 & _EVAL_3391;
  assign _EVAL_560 = _EVAL_2743[425];
  assign _EVAL_1581 = _EVAL_2743[264];
  assign _EVAL_208 = _EVAL_2694 & _EVAL_1856;
  assign _EVAL_2355 = _EVAL_2743[301];
  assign _EVAL_1635 = _EVAL_1596 & _EVAL_1856;
  assign _EVAL_1421 = _EVAL_2234 & _EVAL_1856;
  assign _EVAL_2406 = _EVAL_2743[318];
  assign _EVAL_2973 = _EVAL_3080 & _EVAL_3391;
  assign _EVAL_2680 = _EVAL_2424 & _EVAL_3673;
  assign _EVAL_201 = _EVAL_1187 & _EVAL_1856;
  assign _EVAL_3656 = _EVAL_623 & _EVAL_2474;
  assign _EVAL_391 = _EVAL_2743[5];
  assign _EVAL_1391 = _EVAL_2901 & _EVAL_1856;
  assign _EVAL_3585 = _EVAL_2282 & _EVAL_3673;
  assign _EVAL_170 = _EVAL_2431 & _EVAL_2909;
  assign _EVAL_264 = _EVAL_2428 & _EVAL_2474;
  assign _EVAL_186 = _EVAL_2478 & _EVAL_3673;
  assign _EVAL_2808 = _EVAL_3232 & _EVAL_2909;
  assign _EVAL_3353 = _EVAL_2910 & _EVAL_2474;
  assign _EVAL_235 = _EVAL_2169 & _EVAL_1856;
  assign _EVAL_2108 = _EVAL_1766 & _EVAL_2474;
  assign _EVAL_2320 = _EVAL_873 & _EVAL_3391;
  assign _EVAL_1100 = _EVAL_1455 & _EVAL_2188;
  assign _EVAL_1327 = _EVAL_2167 & _EVAL_1856;
  assign _EVAL_1604 = _EVAL_1309 & _EVAL_3391;
  assign _EVAL_1543 = _EVAL_1782 & _EVAL_2033;
  assign _EVAL_1227 = _EVAL_2743[398];
  assign _EVAL_3639 = _EVAL_307 != 3'h0;
  assign _EVAL_243 = _EVAL_2743[450];
  assign _EVAL_1412 = _EVAL_1700 & _EVAL_3391;
  assign _EVAL_2817 = _EVAL_3147 & _EVAL_1856;
  assign _EVAL_1386 = _EVAL_2743[277];
  assign _EVAL_924 = _EVAL_1327 & _EVAL_3391;
  assign _EVAL_3364 = _EVAL_2236 & _EVAL_3673;
  assign _EVAL_1212 = _EVAL_2743[287];
  assign _EVAL_2213 = _EVAL_43 & _EVAL_3391;
  assign _EVAL_2528 = _EVAL_455 & _EVAL_3391;
  assign _EVAL_2672 = _EVAL_2817 & _EVAL_3391;
  assign _EVAL_2020 = _EVAL_1782 & _EVAL_2140;
  assign _EVAL_3282 = _EVAL_2401 & _EVAL_3391;
  assign _EVAL_2460 = _EVAL_2787 & _EVAL_3391;
  assign _EVAL_581 = _EVAL_873 & _EVAL_2909;
  assign _EVAL_3536 = _EVAL_575[23:13];
  assign _EVAL_1396 = _EVAL_3522 & _EVAL_3391;
  assign _EVAL_976 = _EVAL_2139 & _EVAL_2909;
  assign _EVAL_1704 = _EVAL_355 & _EVAL_2909;
  assign _EVAL_840 = _EVAL_2743[429];
  assign _EVAL_444 = _EVAL_1782 & _EVAL_2592;
  assign _EVAL_2790 = _EVAL_1782 & _EVAL_441;
  assign _EVAL_1222 = _EVAL_1715 & _EVAL_2474;
  assign _EVAL_195 = _EVAL_3040 & _EVAL_3391;
  assign _EVAL_3439 = _EVAL_2303 & _EVAL_2474;
  assign _EVAL_2626 = _EVAL_2656 & _EVAL_3391;
  assign _EVAL_2397 = _EVAL_1740 & _EVAL_3391;
  assign _EVAL_901 = _EVAL_1216 & _EVAL_2474;
  assign _EVAL_2025 = _EVAL_1782 & _EVAL_425;
  assign _EVAL_3010 = _EVAL_3523 & _EVAL_2474;
  assign _EVAL_1986 = _EVAL_2124 & _EVAL_1856;
  assign _EVAL_2072 = _EVAL_2034 & _EVAL_2474;
  assign _EVAL_2827 = _EVAL_1782 & _EVAL_1786;
  assign _EVAL_1458 = _EVAL_288 & _EVAL_2474;
  assign _EVAL_60 = _EVAL_1782 & _EVAL_3142;
  assign _EVAL_2043 = _EVAL_966 & _EVAL_1856;
  assign _EVAL_433 = _EVAL_2555 & _EVAL_3673;
  assign _EVAL_1906 = _EVAL_2551 & _EVAL_2474;
  assign _EVAL_3632 = _EVAL_1782 & _EVAL_3162;
  assign _EVAL_3550 = _EVAL_2551 & _EVAL_3391;
  assign _EVAL_1378 = _EVAL_1782 & _EVAL_973;
  assign _EVAL_905 = _EVAL_2161 & _EVAL_3391;
  assign _EVAL_2186 = _EVAL_2743[482];
  assign _EVAL_1886 = _EVAL_1987 == 2'h3;
  assign _EVAL_390 = _EVAL_2743[350];
  assign _EVAL_1548 = _EVAL_2743[510];
  assign _EVAL_2433 = _EVAL_2743[501];
  assign _EVAL_216 = _EVAL_1782 & _EVAL_3719;
  assign _EVAL_3561 = _EVAL_3735 & _EVAL_1856;
  assign _EVAL_3077 = _EVAL_726 & _EVAL_3391;
  assign _EVAL_2085 = _EVAL_2559 & _EVAL_2909;
  assign _EVAL_2176 = _EVAL_1938 & _EVAL_2474;
  assign _EVAL_3735 = _EVAL_1782 & _EVAL_316;
  assign _EVAL_3608 = _EVAL_255 & _EVAL_1856;
  assign _EVAL_2315 = _EVAL_1782 & _EVAL_1227;
  assign _EVAL_3691 = _EVAL_2660 & _EVAL_1856;
  assign _EVAL_398 = _EVAL_3449 & _EVAL_1856;
  assign _EVAL_3629 = _EVAL_288 & _EVAL_3673;
  assign _EVAL_430 = _EVAL_2743[223];
  assign _EVAL_3702 = _EVAL_376 & _EVAL_2909;
  assign _EVAL_610 = _EVAL_2137 & _EVAL_1856;
  assign _EVAL_2981 = _EVAL_254 & _EVAL_1856;
  assign _EVAL_589 = _EVAL_1294 & _EVAL_2474;
  assign _EVAL_1345 = _EVAL_1782 & _EVAL_2614;
  assign _EVAL_2620 = _EVAL_3015 & _EVAL_3673;
  assign _EVAL_2353 = _EVAL_1153 & _EVAL_1856;
  assign _EVAL_129 = _EVAL_2743[469];
  assign _EVAL_755 = _EVAL_2600 & _EVAL_2909;
  assign TLMonitor_1__EVAL_10 = _EVAL_5;
  assign _EVAL_149 = _EVAL_1964 & _EVAL_3673;
  assign _EVAL_1624 = _EVAL_3592 & _EVAL_3391;
  assign _EVAL_2572 = _EVAL_1165 & _EVAL_3391;
  assign _EVAL_316 = _EVAL_2743[500];
  assign _EVAL_1793 = _EVAL_1984 & _EVAL_1856;
  assign _EVAL_2634 = _EVAL_2743[439];
  assign _EVAL_2393 = _EVAL_1216 & _EVAL_3673;
  assign _EVAL_3191 = _EVAL_2568 & _EVAL_2474;
  assign _EVAL_405 = _EVAL_398 & _EVAL_2474;
  assign _EVAL_1338 = _EVAL_712 & _EVAL_3391;
  assign _EVAL_3240 = _EVAL_2613 & _EVAL_2474;
  assign _EVAL_188 = _EVAL_2743[192];
  assign _EVAL_1438 = _EVAL_1301 & _EVAL_2909;
  assign _EVAL_1695 = _EVAL_2743[464];
  assign TLMonitor__EVAL_9 = _EVAL_41;
  assign _EVAL_2901 = _EVAL_1782 & _EVAL_1093;
  assign _EVAL_1329 = _EVAL_2952 & _EVAL_1856;
  assign _EVAL_1483 = _EVAL_2643 & _EVAL_356;
  assign _EVAL_1252 = _EVAL_305 & _EVAL_3673;
  assign _EVAL_3192 = _EVAL_3835 & _EVAL_2909;
  assign _EVAL_2413 = _EVAL_298 & _EVAL_2474;
  assign _EVAL_615 = _EVAL_2084 & _EVAL_2909;
  assign _EVAL_326 = _EVAL_2743[360];
  assign _EVAL_1768 = _EVAL_100 & _EVAL_3673;
  assign _EVAL_666 = _EVAL_2661 & _EVAL_3673;
  assign _EVAL_1103 = _EVAL_3734 & _EVAL_2474;
  assign _EVAL_3205 = _EVAL_872 & _EVAL_3673;
  assign _EVAL_2049 = _EVAL_1301 & _EVAL_3391;
  assign _EVAL_1142 = _EVAL_1892 & _EVAL_3673;
  assign _EVAL_1714 = _EVAL_2743[357];
  assign _EVAL_3766 = _EVAL_3185 & _EVAL_2474;
  assign _EVAL_3297 = _EVAL_948 & _EVAL_2474;
  assign _EVAL_548 = _EVAL_77 & _EVAL_1856;
  assign _EVAL_1405 = _EVAL_992 & _EVAL_1856;
  assign _EVAL_3794 = _EVAL_1782 & _EVAL_2355;
  assign _EVAL_632 = _EVAL_2478 & _EVAL_2909;
  assign _EVAL_1054 = _EVAL_3466 & _EVAL_2474;
  assign _EVAL_1352 = _EVAL_2526 & _EVAL_1856;
  assign _EVAL_2768 = _EVAL_2633 & _EVAL_1856;
  assign _EVAL_1588 = _EVAL_1765 & _EVAL_3673;
  assign _EVAL_341 = _EVAL_3803 & _EVAL_3673;
  assign _EVAL_3460 = _EVAL_2352 & _EVAL_2909;
  assign _EVAL_1300 = _EVAL_2743[383];
  assign _EVAL_1566 = _EVAL_1782 & _EVAL_2665;
  assign _EVAL_2350 = _EVAL_667 & _EVAL_3673;
  assign _EVAL_1580 = _EVAL_2568 & _EVAL_3391;
  assign _EVAL_1397 = _EVAL_1782 & _EVAL_539;
  assign _EVAL_1912 = _EVAL_610 & _EVAL_3391;
  assign _EVAL_3790 = _EVAL_3544 & _EVAL_3391;
  assign _EVAL_2462 = _EVAL_2667 & _EVAL_2474;
  assign _EVAL_103 = _EVAL_3018 & _EVAL_1856;
  assign _EVAL_2803 = _EVAL_3696 & _EVAL_3673;
  assign _EVAL_3202 = _EVAL_274 & _EVAL_3673;
  assign TLMonitor_1__EVAL_11 = _EVAL_39;
  assign _EVAL_3198 = _EVAL_1782 & _EVAL_129;
  assign _EVAL_1668 = _EVAL_1951 & _EVAL_3673;
  assign _EVAL_2158 = _EVAL_2743[258];
  assign _EVAL_2917 = _EVAL_3351 & _EVAL_3673;
  assign _EVAL_503 = _EVAL_2743[4];
  assign _EVAL_2466 = _EVAL_2743[298];
  assign _EVAL_2542 = _EVAL_3327 & _EVAL_3391;
  assign _EVAL_2088 = _EVAL_1102 & _EVAL_3673;
  assign _EVAL_2701 = _EVAL_1782 & _EVAL_1068;
  assign _EVAL_3463 = _EVAL_2421 & _EVAL_2474;
  assign _EVAL_3332 = _EVAL_2580 & _EVAL_1856;
  assign _EVAL_2474 = _EVAL_2864 != 8'h0;
  assign _EVAL_3713 = _EVAL_3597 & _EVAL_3391;
  assign _EVAL_954 = _EVAL_1126 & _EVAL_3673;
  assign _EVAL_1660 = _EVAL_2554 & _EVAL_3391;
  assign _EVAL_2586 = _EVAL_1782 & _EVAL_1111;
  assign _EVAL_3125 = _EVAL_2768 & _EVAL_3673;
  assign _EVAL_1940 = _EVAL_575[15];
  assign TLMonitor_1__EVAL_9 = _EVAL_14;
  assign _EVAL_138 = _EVAL_83[16];
  assign _EVAL_1640 = _EVAL_2918 & _EVAL_3673;
  assign _EVAL_1286 = _EVAL_3630 & _EVAL_3391;
  assign _EVAL_902 = _EVAL_1246 & _EVAL_2474;
  assign _EVAL_529 = _EVAL_2799 & _EVAL_2474;
  assign _EVAL_1854 = _EVAL_3587 & _EVAL_3673;
  assign _EVAL_288 = _EVAL_2548 & _EVAL_1856;
  assign _EVAL_2364 = _EVAL_1782 & _EVAL_1903;
  assign _EVAL_1570 = _EVAL_1782 & _EVAL_2262;
  assign _EVAL_2658 = _EVAL_1657 & _EVAL_3673;
  assign _EVAL_1161 = _EVAL_2743[328];
  assign _EVAL_414 = _EVAL_2537 & _EVAL_1856;
  assign TLMonitor_1__EVAL_7 = _EVAL_32;
  assign _EVAL_1459 = _EVAL_2046 & _EVAL_3673;
  assign _EVAL_1229 = _EVAL_1951 & _EVAL_3391;
  assign _EVAL_1628 = _EVAL_2743[465];
  assign _EVAL_883 = _EVAL_314 & _EVAL_3673;
  assign _EVAL_1826 = _EVAL_287 & _EVAL_3391;
  assign _EVAL_2596 = _EVAL_1432 & _EVAL_2909;
  assign _EVAL_1427 = _EVAL_3245 & _EVAL_2474;
  assign _EVAL_2301 = _EVAL_1006 & _EVAL_2474;
  assign _EVAL_898 = _EVAL_3691 & _EVAL_2909;
  assign _EVAL_1707 = _EVAL_2059 & _EVAL_2474;
  assign TLMonitor_1__EVAL_1 = _EVAL_38;
  assign _EVAL_3552 = _EVAL_2922 & _EVAL_3673;
  assign _EVAL_2352 = _EVAL_3161 & _EVAL_1856;
  assign _EVAL_346 = _EVAL_235 & _EVAL_3673;
  assign _EVAL_854 = _EVAL_2743[351];
  assign _EVAL_348 = _EVAL_1973 & _EVAL_3391;
  assign _EVAL_2161 = _EVAL_3533 & _EVAL_1856;
  assign _EVAL_938 = _EVAL_1201 & _EVAL_3673;
  assign _EVAL_907 = _EVAL_998 & _EVAL_2909;
  assign _EVAL_1245 = _EVAL_3544 & _EVAL_2474;
  assign _EVAL_2241 = _EVAL_2743[333];
  assign _EVAL_2734 = _EVAL_1782 & _EVAL_1895;
  assign _EVAL_2229 = _EVAL_3468 & _EVAL_1856;
  assign _EVAL_1193 = _EVAL_2743[367];
  assign _EVAL_2556 = _EVAL_1188 & _EVAL_2474;
  assign _EVAL_1960 = _EVAL_1782 & _EVAL_737;
  assign _EVAL_948 = _EVAL_821 & _EVAL_1856;
  assign _EVAL_1079 = _EVAL_2119 & _EVAL_3391;
  assign _EVAL_2276 = _EVAL_2743[396];
  assign _EVAL_1785 = _EVAL_2643 & _EVAL_920;
  assign _EVAL_694 = _EVAL_3802 & _EVAL_2909;
  assign _EVAL_2477 = _EVAL_1782 & _EVAL_1402;
  assign _EVAL_961 = _EVAL_1782 & _EVAL_1511;
  assign _EVAL_2382 = _EVAL_2743[375];
  assign _EVAL_2601 = _EVAL_455 & _EVAL_2909;
  assign _EVAL_3685 = _EVAL_103 & _EVAL_2909;
  assign _EVAL_2873 = _EVAL_2743[325];
  assign _EVAL_2361 = _EVAL_3015 & _EVAL_3391;
  assign _EVAL_501 = _EVAL_3718 & _EVAL_2474;
  assign _EVAL_3368 = _EVAL_2586 & _EVAL_1856;
  assign _EVAL_1656 = _EVAL_1210 & _EVAL_1856;
  assign _EVAL_134 = _EVAL_1782 & _EVAL_801;
  assign TLMonitor__EVAL = _EVAL_40;
  assign _EVAL_1165 = _EVAL_2315 & _EVAL_1856;
  assign _EVAL_3645 = _EVAL_426 & _EVAL_1856;
  assign _EVAL_1717 = _EVAL_297 & _EVAL_2474;
  assign _EVAL_2600 = _EVAL_2912 & _EVAL_3670;
  assign _EVAL_3430 = _EVAL_504 & _EVAL_1856;
  assign _EVAL_1117 = _EVAL_3529 & _EVAL_3673;
  assign _EVAL_2391 = _EVAL_1439 & _EVAL_2909;
  assign _EVAL_3110 = _EVAL_137 & _EVAL_3673;
  assign _EVAL_3572 = _EVAL_2661 & _EVAL_2909;
  assign _EVAL_2058 = _EVAL_1782 & _EVAL_994;
  assign _EVAL_1322 = _EVAL_3632 & _EVAL_1856;
  assign _EVAL_3091 = _EVAL_1782 & _EVAL_2466;
  assign _EVAL_787 = _EVAL_2037 & _EVAL_3673;
  assign _EVAL_2529 = _EVAL_2303 & _EVAL_3391;
  assign _EVAL_2107 = _EVAL_3561 & _EVAL_3391;
  assign _EVAL_776 = _EVAL_878 & _EVAL_3391;
  assign _EVAL_345 = _EVAL_1782 & _EVAL_1855;
  assign _EVAL_3415 = _EVAL_3821 & _EVAL_3391;
  assign _EVAL_855 = _EVAL_1782 & _EVAL_46;
  assign _EVAL_3642 = _EVAL_1782 & _EVAL_242;
  assign _EVAL_1013 = _EVAL_1782 & _EVAL_825;
  assign _EVAL_647 = _EVAL_1782 & _EVAL_2873;
  assign _EVAL_3446 = _EVAL_2165 & _EVAL_3391;
  assign _EVAL_2313 = _EVAL_208 & _EVAL_3673;
  assign _EVAL_2574 = _EVAL_3553 & _EVAL_3673;
  assign _EVAL_2094 = _EVAL_103 & _EVAL_3391;
  assign _EVAL_805 = _EVAL_1700 & _EVAL_2474;
  assign _EVAL_1926 = _EVAL_2693 & _EVAL_3673;
  assign _EVAL_2605 = _EVAL_2743[18];
  assign _EVAL_3797 = _EVAL_2849 & _EVAL_2909;
  assign TLMonitor_1__EVAL_3 = _EVAL_28;
  assign _EVAL_3737 = _EVAL_1700 & _EVAL_3673;
  assign _EVAL_340 = _EVAL_1299 & _EVAL_2474;
  assign _EVAL_1709 = _EVAL_919 & _EVAL_897;
  assign _EVAL_740 = _EVAL_783 & _EVAL_1856;
  assign _EVAL_3796 = _EVAL_2093 & _EVAL_2909;
  assign _EVAL_2834 = _EVAL_2743[294];
  assign _EVAL_2362 = _EVAL_2427 & _EVAL_2400;
  assign _EVAL_203 = _EVAL_1204 & _EVAL_2474;
  assign _EVAL_807 = _EVAL_2016 & _EVAL_2474;
  assign _EVAL_89 = _EVAL_1022 & _EVAL_1856;
  assign _EVAL_1387 = _EVAL_511 & _EVAL_3391;
  assign _EVAL_2159 = _EVAL_2305 & _EVAL_2474;
  assign _EVAL_3315 = _EVAL_1782 & _EVAL_391;
  assign _EVAL_884 = _EVAL_988 & _EVAL_3673;
  assign _EVAL_1234 = _EVAL_2743[384];
  assign _EVAL_2009 = _EVAL_576 & _EVAL_2474;
  assign _EVAL_3434 = _EVAL_1405 & _EVAL_3391;
  assign _EVAL_741 = _EVAL_3055 & _EVAL_3391;
  assign _EVAL_977 = _EVAL_1208 & _EVAL_1856;
  assign _EVAL_2060 = _EVAL_2817 & _EVAL_2909;
  assign _EVAL_2424 = _EVAL_844 & _EVAL_1856;
  assign _EVAL_2930 = _EVAL_911 & _EVAL_2474;
  assign _EVAL_2016 = _EVAL_2647 & _EVAL_3670;
  assign _EVAL_2369 = _EVAL_3345 & _EVAL_2909;
  assign _EVAL_1702 = _EVAL_1782 & _EVAL_840;
  assign _EVAL_781 = _EVAL_1782 & _EVAL_595;
  assign _EVAL_3151 = _EVAL_2477 & _EVAL_1856;
  assign _EVAL_3822 = _EVAL_2743[361];
  assign _EVAL_2394 = _EVAL_2206 & _EVAL_3673;
  assign _EVAL_3529 = _EVAL_2733 & _EVAL_1856;
  assign _EVAL_1737 = _EVAL_1100 & _EVAL_2639;
  assign _EVAL_1209 = _EVAL_575[21:20];
  assign _EVAL_1068 = _EVAL_2743[401];
  assign _EVAL_1735 = _EVAL_511 & _EVAL_3673;
  assign _EVAL_1770 = _EVAL_2034 & _EVAL_3673;
  assign _EVAL_3680 = _EVAL_43 & _EVAL_3673;
  assign _EVAL_1248 = _EVAL_979 & _EVAL_1601;
  assign _EVAL_747 = _EVAL_2910 & _EVAL_3673;
  assign _EVAL_3719 = _EVAL_2743[374];
  assign _EVAL_357 = _EVAL_2743[3];
  assign _EVAL_928 = _EVAL_678 & _EVAL_2909;
  assign _EVAL_2421 = _EVAL_626 & _EVAL_1856;
  assign _EVAL_1509 = _EVAL_2271 & _EVAL_3391;
  assign TLMonitor_1__EVAL = _EVAL_20;
  assign _EVAL_309 = _EVAL_575[3:0];
  assign _EVAL_64 = _EVAL_2743[8];
  assign _EVAL_3287 = _EVAL_3642 & _EVAL_3670;
  assign _EVAL_2865 = _EVAL_1322 & _EVAL_3673;
  assign _EVAL_3170 = _EVAL_2743[289];
  assign _EVAL_2010 = _EVAL_322 & _EVAL_2909;
  assign _EVAL_2980 = _EVAL_1782 & _EVAL_2514;
  assign _EVAL_3335 = _EVAL_2554 & _EVAL_2909;
  assign _EVAL_2191 = _EVAL_3553 & _EVAL_3391;
  assign _EVAL_3468 = _EVAL_1782 & _EVAL_3798;
  assign _EVAL_3380 = _EVAL_163 & _EVAL_3391;
  assign _EVAL_1962 = _EVAL_1782 & _EVAL_732;
  assign _EVAL_1889 = _EVAL_89 & _EVAL_3673;
  assign _EVAL_469 = _EVAL_2998 & _EVAL_2474;
  assign _EVAL_2242 = _EVAL_2236 & _EVAL_2474;
  assign _EVAL_454 = _EVAL_1782 & _EVAL_854;
  assign TLMonitor_1__EVAL_2 = _EVAL_34;
  assign _EVAL_3291 = _EVAL_3522 & _EVAL_2474;
  assign _EVAL_3659 = _EVAL_1064 & _EVAL_3673;
  assign _EVAL_1246 = _EVAL_2493 & _EVAL_1856;
  assign _EVAL_794 = _EVAL_2743[487];
  assign _EVAL_1531 = _EVAL_1782 & _EVAL_637;
  assign _EVAL_2857 = _EVAL_1793 & _EVAL_2474;
  assign _EVAL_381 = _EVAL_2396 & _EVAL_2474;
  assign _EVAL_162 = _EVAL_1264 & _EVAL_3391;
  assign _EVAL_1093 = _EVAL_2743[511];
  assign _EVAL_1076 = _EVAL_2667 & _EVAL_3673;
  assign _EVAL_2141 = _EVAL_1503 & _EVAL_3391;
  assign _EVAL_3679 = _EVAL_2743[275];
  assign _EVAL_101 = _EVAL_2743[20];
  assign _EVAL_703 = _EVAL_3430 & _EVAL_3673;
  assign _EVAL_168 = _EVAL_1349 & _EVAL_1856;
  assign _EVAL_2208 = _EVAL_2431 & _EVAL_2474;
  assign _EVAL_1009 = _EVAL_1782 & _EVAL_3733;
  assign _EVAL_775 = _EVAL_2568 & _EVAL_3673;
  assign _EVAL_2381 = _EVAL_779 & _EVAL_3391;
  assign _EVAL_3497 = _EVAL_3553 & _EVAL_2474;
  assign _EVAL_2513 = _EVAL_250 & _EVAL_3391;
  assign _EVAL_578 = _EVAL_1782 & _EVAL_1689;
  assign _EVAL_387 = _EVAL_1100 & _EVAL_145;
  assign _EVAL_2800 = _EVAL_535 & _EVAL_3673;
  assign _EVAL_3626 = _EVAL_872 & _EVAL_2474;
  assign _EVAL_1056 = _EVAL_2743[459];
  assign _EVAL_1394 = _EVAL_2918 & _EVAL_2909;
  assign _EVAL_2055 = _EVAL_136 & _EVAL_1856;
  assign _EVAL_2227 = _EVAL_1782 & _EVAL_3312;
  assign _EVAL_1895 = _EVAL_2743[311];
  assign _EVAL_989 = _EVAL_3114 & _EVAL_3391;
  assign _EVAL_756 = _EVAL_3190 & _EVAL_120;
  assign _EVAL_2461 = _EVAL_998 & _EVAL_3673;
  assign _EVAL_3597 = _EVAL_2135 & _EVAL_1856;
  assign _EVAL_1295 = _EVAL_1782 & _EVAL_1536;
  assign _EVAL_2146 = _EVAL_1782 & _EVAL_1974;
  assign _EVAL_3367 = _EVAL_2738 & _EVAL_2474;
  assign _EVAL_1618 = _EVAL_2743[471];
  assign _EVAL_979 = _EVAL_2792 & _EVAL_2188;
  assign TLMonitor__EVAL_5 = _EVAL_40;
  assign _EVAL_1539 = _EVAL_3365 & _EVAL_2909;
  assign _EVAL_298 = _EVAL_2609 & _EVAL_1856;
  assign _EVAL_1187 = _EVAL_1782 & _EVAL_80;
  assign _EVAL_2435 = _EVAL_496 & _EVAL_1856;
  assign _EVAL_945 = _EVAL_1201 & _EVAL_3391;
  assign _EVAL_3602 = _EVAL_3522 & _EVAL_3673;
  assign _EVAL_2036 = _EVAL_1644 & _EVAL_3391;
  assign _EVAL_936 = _EVAL_1892 & _EVAL_2909;
  assign _EVAL_42 = _EVAL_576 & _EVAL_3673;
  assign _EVAL_2990 = _EVAL_1780 & _EVAL_2909;
  assign _EVAL_3512 = _EVAL_2743[279];
  assign _EVAL_2067 = _EVAL_445 & _EVAL_3673;
  assign _EVAL_2647 = _EVAL_1782 & _EVAL_2605;
  assign _EVAL_1947 = _EVAL_1915 & _EVAL_2474;
  assign _EVAL_1999 = _EVAL_1432 & _EVAL_2474;
  assign _EVAL_1236 = _EVAL_103 & _EVAL_3673;
  assign _EVAL_1062 = _EVAL_2421 & _EVAL_3673;
  assign _EVAL_2129 = _EVAL_2953 & _EVAL_2909;
  assign _EVAL_2028 = _EVAL_1345 & _EVAL_1856;
  assign _EVAL_3188 = _EVAL_1102 & _EVAL_3391;
  assign _EVAL_1296 = _EVAL_3561 & _EVAL_2909;
  assign _EVAL_91 = _EVAL_398 & _EVAL_3673;
  assign _EVAL_1510 = _EVAL_3529 & _EVAL_3391;
  assign _EVAL_1662 = _EVAL_1782 & _EVAL_1411;
  assign _EVAL_2944 = _EVAL_2743[472];
  assign _EVAL_2507 = _EVAL_2666 & _EVAL_2474;
  assign _EVAL_872 = _EVAL_647 & _EVAL_1856;
  assign _EVAL_2509 = _EVAL_3592 & _EVAL_3673;
  assign _EVAL_3164 = _EVAL_1782 & _EVAL_695;
  assign _EVAL_81 = _EVAL_1207 & _EVAL_2909;
  assign _EVAL_3190 = _EVAL_1292 & _EVAL_2188;
  assign _EVAL_1555 = _EVAL_521 & _EVAL_120;
  assign _EVAL_3370 = _EVAL_3168 & _EVAL_1856;
  assign _EVAL_975 = _EVAL_3597 & _EVAL_2909;
  assign _EVAL_3684 = _EVAL_1722 & _EVAL_1856;
  assign _EVAL_3580 = _EVAL_2962 & _EVAL_3391;
  assign _EVAL_2563 = _EVAL_3608 & _EVAL_2474;
  assign _EVAL_163 = _EVAL_1686 & _EVAL_1856;
  assign _EVAL_3667 = _EVAL_3812 & _EVAL_2909;
  assign _EVAL_1279 = _EVAL_2666 & _EVAL_3391;
  assign _EVAL_3658 = _EVAL_2206 & _EVAL_3391;
  assign _EVAL_379 = _EVAL_1172 & _EVAL_2909;
  assign _EVAL_1910 = _EVAL_2743[443];
  assign _EVAL_1249 = _EVAL_3553 & _EVAL_2909;
  assign _EVAL_1676 = _EVAL_3620 & _EVAL_2474;
  assign _EVAL_2151 = _EVAL_3358 & _EVAL_3673;
  assign _EVAL_1242 = _EVAL_2743[386];
  assign _EVAL_1529 = _EVAL_3315 & _EVAL_3670;
  assign _EVAL_3346 = _EVAL_2338 & _EVAL_2909;
  assign _EVAL_3435 = _EVAL_1782 & _EVAL_675;
  assign _EVAL_1363 = _EVAL_655 & _EVAL_1856;
  assign _EVAL_3092 = _EVAL_1235 & _EVAL_2474;
  assign _EVAL_3636 = _EVAL_2424 & _EVAL_2909;
  assign _EVAL_1320 = _EVAL_2307 & _EVAL_3391;
  assign _EVAL_3384 = _EVAL_877 & _EVAL_2909;
  assign _EVAL_3292 = _EVAL_2743[449];
  assign TLMonitor__EVAL_6 = _EVAL_0;
  assign _EVAL_3778 = _EVAL_1013 & _EVAL_1856;
  assign _EVAL_1128 = _EVAL_2743[475];
  assign _EVAL_573 = _EVAL_3167 & _EVAL_2474;
  assign _EVAL_2585 = _EVAL_1524 & _EVAL_3673;
  assign _EVAL_1851 = _EVAL_2743[392];
  assign _EVAL_3226 = _EVAL_1782 & _EVAL_1148;
  assign _EVAL_664 = _EVAL_2729 & _EVAL_1256;
  assign _EVAL_53 = _EVAL_1782 & _EVAL_2300;
  assign _EVAL_1372 = _EVAL_2743[1];
  assign _EVAL_2608 = _EVAL_1065 & _EVAL_2909;
  assign _EVAL_1698 = _EVAL_652 & _EVAL_3391;
  assign _EVAL_2253 = _EVAL_2637 & _EVAL_1856;
  assign _EVAL_3139 = _EVAL_1264 & _EVAL_2474;
  assign _EVAL_639 = _EVAL_1064 & _EVAL_3391;
  assign _EVAL_1643 = _EVAL_3345 & _EVAL_3673;
  assign _EVAL_108 = _EVAL_2084 & _EVAL_3391;
  assign _EVAL_1955 = _EVAL_2743[338];
  assign _EVAL_556 = _EVAL_1452 & _EVAL_3673;
  assign _EVAL_986 = _EVAL_2084 & _EVAL_3673;
  assign _EVAL_422 = _EVAL_43 & _EVAL_2474;
  assign _EVAL_2131 = _EVAL_3261 & _EVAL_3391;
  assign _EVAL_3692 = _EVAL_1743 & _EVAL_2474;
  assign _EVAL_1463 = _EVAL_2729 & _EVAL_3398;
  assign _EVAL_513 = _EVAL_1782 & _EVAL_1059;
  assign _EVAL_482 = _EVAL_3523 & _EVAL_3391;
  assign _EVAL_1342 = _EVAL_1782 & _EVAL_3141;
  assign _EVAL_2252 = _EVAL_911 & _EVAL_3673;
  assign _EVAL_3416 = _EVAL_1782 & _EVAL_1637;
  assign _EVAL_1515 = _EVAL_1329 & _EVAL_2474;
  assign _EVAL_1680 = _EVAL_3544 & _EVAL_3673;
  assign _EVAL_1105 = _EVAL_3332 & _EVAL_2909;
  assign _EVAL_1169 = _EVAL_2743[353];
  assign _EVAL_810 = _EVAL_1352 & _EVAL_2909;
  assign _EVAL_656 = _EVAL_1782 & _EVAL_3619;
  assign _EVAL_2415 = _EVAL_3351 & _EVAL_3391;
  assign _EVAL_1075 = _EVAL_2743[369];
  assign _EVAL_3006 = _EVAL_2743[340];
  assign _EVAL_2867 = _EVAL_2353 & _EVAL_2474;
  assign _EVAL_745 = _EVAL_3684 & _EVAL_2909;
  assign _EVAL_783 = _EVAL_1782 & _EVAL_461;
  assign _EVAL_726 = _EVAL_1009 & _EVAL_1856;
  assign _EVAL_62 = _EVAL_720 & _EVAL_2909;
  assign _EVAL_962 = _EVAL_2743[407];
  assign _EVAL_1988 = _EVAL_3361 & _EVAL_3673;
  assign _EVAL_2335 = _EVAL_684 & _EVAL_2474;
  assign _EVAL_2046 = _EVAL_1108 & _EVAL_1856;
  assign _EVAL_1827 = _EVAL_3399 & _EVAL_3391;
  assign _EVAL_1616 = _EVAL_250 & _EVAL_3673;
  assign _EVAL_2376 = _EVAL_1529 & _EVAL_2474;
  assign _EVAL_1783 = _EVAL_2515 & _EVAL_1856;
  assign _EVAL_336 = _EVAL_1782 & _EVAL_794;
  assign _EVAL_2426 = ~_EVAL_2500;
  assign _EVAL_1291 = _EVAL_1207 & _EVAL_2474;
  assign _EVAL_2428 = _EVAL_2534 & _EVAL_1856;
  assign _EVAL_3706 = _EVAL_274 & _EVAL_2909;
  assign _EVAL_1831 = _EVAL_2743[310];
  assign _EVAL_1067 = _EVAL_2738 & _EVAL_3391;
  assign _EVAL_1085 = _EVAL_3357 & _EVAL_3673;
  assign _EVAL_1083 = _EVAL_2201 & _EVAL_3673;
  assign _EVAL_1667 = _EVAL_1782 & _EVAL_2663;
  assign _EVAL_2555 = _EVAL_1772 & _EVAL_1856;
  assign _EVAL_1415 = _EVAL_1188 & _EVAL_2909;
  assign _EVAL_301 = _EVAL_1782 & _EVAL_2982;
  assign _EVAL_2330 = _EVAL_1782 & _EVAL_2026;
  assign _EVAL_3099 = _EVAL_911 & _EVAL_3391;
  assign _EVAL_2537 = _EVAL_1782 & _EVAL_1910;
  assign _EVAL_3781 = _EVAL_2675 & _EVAL_2909;
  assign _EVAL_2500 = _EVAL_1032 | _EVAL_38;
  assign _EVAL_1330 = _EVAL_2729 & _EVAL_449;
  assign _EVAL_3055 = _EVAL_826 & _EVAL_1856;
  assign _EVAL_3199 = _EVAL_3684 & _EVAL_3391;
  assign _EVAL_3683 = _EVAL_74 & _EVAL_2909;
  assign _EVAL_1108 = _EVAL_1782 & _EVAL_1851;
  assign _EVAL_1690 = _EVAL_1340 & _EVAL_2474;
  assign _EVAL_2309 = _EVAL_1938 & _EVAL_3391;
  assign _EVAL_1909 = _EVAL_2880 & _EVAL_2474;
  assign _EVAL_2436 = _EVAL_3360 & _EVAL_3673;
  assign _EVAL_3438 = _EVAL_575[16];
  assign _EVAL_1091 = _EVAL_1782 & _EVAL_1581;
  assign _EVAL_1753 = _EVAL_1716 & _EVAL_2474;
  assign _EVAL_2127 = _EVAL_2743[284];
  assign _EVAL_2209 = _EVAL_779 & _EVAL_2909;
  assign _EVAL_3681 = _EVAL_575[12];
  assign _EVAL_2434 = _EVAL_2338 & _EVAL_3391;
  assign _EVAL_376 = _EVAL_543 & _EVAL_1856;
  assign _EVAL_3058 = _EVAL_3185 & _EVAL_2909;
  assign _EVAL_2665 = _EVAL_2743[335];
  assign _EVAL_1402 = _EVAL_2743[316];
  assign _EVAL_242 = _EVAL_2743[9];
  assign _EVAL_1344 = _EVAL_2718 & _EVAL_2474;
  assign _EVAL_1417 = _EVAL_623 & _EVAL_2909;
  assign _EVAL_1683 = _EVAL_3812 & _EVAL_3391;
  assign _EVAL_3334 = _EVAL_878 & _EVAL_2474;
  assign _EVAL_3374 = _EVAL_3365 & _EVAL_2474;
  assign _EVAL_3556 = _EVAL_1201 & _EVAL_2474;
  assign _EVAL_3036 = _EVAL_3696 & _EVAL_2474;
  assign _EVAL_119 = _EVAL_3778 & _EVAL_3673;
  assign _EVAL_3111 = _EVAL_297 & _EVAL_3673;
  assign _EVAL_3314 = _EVAL_678 & _EVAL_2474;
  assign _EVAL_600 = _EVAL_3430 & _EVAL_2909;
  assign _EVAL_3014 = _EVAL_1363 & _EVAL_3673;
  assign _EVAL_877 = _EVAL_2575 & _EVAL_1856;
  assign _EVAL_539 = _EVAL_2743[283];
  assign _EVAL_2288 = _EVAL_977 & _EVAL_2474;
  assign _EVAL_3527 = _EVAL_1585 & _EVAL_1856;
  assign _EVAL_3062 = _EVAL_1391 & _EVAL_3673;
  assign _EVAL_675 = _EVAL_2743[444];
  assign _EVAL_3028 = _EVAL_3357 & _EVAL_2474;
  assign _EVAL_106 = _EVAL_1209 != 2'h0;
  assign _EVAL_3424 = _EVAL_2743[421];
  assign _EVAL_2726 = _EVAL_953 & _EVAL_3391;
  assign _EVAL_2967 = _EVAL_1356 & _EVAL_3673;
  assign _EVAL_1563 = _EVAL_872 & _EVAL_3391;
  assign _EVAL_193 = _EVAL_2046 & _EVAL_2474;
  assign _EVAL_3740 = _EVAL_1782 & _EVAL_3118;
  assign _EVAL_254 = _EVAL_1782 & _EVAL_2045;
  assign _EVAL_3156 = _EVAL_1172 & _EVAL_2474;
  assign _EVAL_2793 = _EVAL_2743[403];
  assign _EVAL_3759 = _EVAL_873 & _EVAL_3673;
  assign _EVAL_2554 = _EVAL_454 & _EVAL_1856;
  assign _EVAL_1201 = _EVAL_1969 & _EVAL_1856;
  assign _EVAL_1090 = _EVAL_1782 & _EVAL_3292;
  assign TLMonitor_1__EVAL_12 = _EVAL_34;
  assign _EVAL_2405 = _EVAL_3534 & _EVAL_2909;
  assign _EVAL_715 = _EVAL_208 & _EVAL_2474;
  assign _EVAL_1739 = _EVAL_953 & _EVAL_2474;
  assign _EVAL_1130 = _EVAL_3345 & _EVAL_3391;
  assign _EVAL_2059 = _EVAL_3012 & _EVAL_1856;
  assign _EVAL_3305 = _EVAL_3358 & _EVAL_3391;
  assign _EVAL_3543 = _EVAL_2718 & _EVAL_2909;
  assign _EVAL_1969 = _EVAL_1782 & _EVAL_913;
  assign _EVAL_1740 = _EVAL_781 & _EVAL_1856;
  assign _EVAL_2022 = _EVAL_1782 & _EVAL_3571;
  assign _EVAL_2117 = _EVAL_1782 & _EVAL_1161;
  assign _EVAL_1287 = _EVAL_314 & _EVAL_2909;
  assign _EVAL_935 = _EVAL_2043 & _EVAL_2909;
  assign _EVAL_1078 = _EVAL_2743[344];
  assign _EVAL_84 = _EVAL_2016 & _EVAL_3391;
  assign _EVAL_3478 = _EVAL_163 & _EVAL_2474;
  assign _EVAL_2199 = _EVAL_1782 & _EVAL_443;
  assign _EVAL_1558 = _EVAL_3327 & _EVAL_2474;
  assign _EVAL_3081 = _EVAL_1322 & _EVAL_2909;
  assign _EVAL_680 = _EVAL_2743[460];
  assign _EVAL_1864 = _EVAL_667 & _EVAL_2474;
  assign _EVAL_416 = _EVAL_2307 & _EVAL_3673;
  assign _EVAL_1080 = _EVAL_3360 & _EVAL_2909;
  assign _EVAL_3034 = _EVAL_2425 & _EVAL_2474;
  assign _EVAL_2891 = _EVAL_3399 & _EVAL_2474;
  assign _EVAL_1499 = _EVAL_163 & _EVAL_2909;
  assign _EVAL_3153 = _EVAL_250 & _EVAL_2909;
  assign _EVAL_3184 = _EVAL_69 & _EVAL_2474;
  assign _EVAL_104 = _EVAL_208 & _EVAL_3391;
  assign _EVAL_557 = _EVAL_2134 & _EVAL_3673;
  assign _EVAL_596 = _EVAL_453 & _EVAL_1856;
  assign _EVAL_3473 = _EVAL_1782 & _EVAL_670;
  assign _EVAL_461 = _EVAL_2743[336];
  assign _EVAL_1379 = _EVAL_2743[440];
  assign _EVAL_177 = _EVAL_1782 & _EVAL_2550;
  assign _EVAL_2907 = _EVAL_2936 & _EVAL_3391;
  assign _EVAL_1885 = _EVAL_1635 & _EVAL_3391;
  assign _EVAL_2579 = _EVAL_2729 & _EVAL_1825;
  assign _EVAL_2214 = _EVAL_3406 == 10'h0;
  assign _EVAL_2169 = _EVAL_1782 & _EVAL_2488;
  assign _EVAL_2729 = _EVAL_1483 & _EVAL_2188;
  assign _EVAL_160 = _EVAL_322 & _EVAL_3391;
  assign _EVAL_367 = _EVAL_1782 & _EVAL_352;
  assign _EVAL_1664 = _EVAL_3728 & _EVAL_3391;
  assign TLMonitor__EVAL_7 = _EVAL_29;
  assign _EVAL_1772 = _EVAL_1782 & _EVAL_2618;
  assign _EVAL_520 = _EVAL_1363 & _EVAL_2474;
  assign _EVAL_3361 = _EVAL_3787 & _EVAL_3670;
  assign _EVAL_1820 = _EVAL_3041 & _EVAL_2474;
  assign _EVAL_1744 = _EVAL_2972 & _EVAL_3673;
  assign _EVAL_277 = _EVAL_103 & _EVAL_2474;
  assign _EVAL_1302 = _EVAL_1716 & _EVAL_2909;
  assign _EVAL_1232 = _EVAL_2743[288];
  assign _EVAL_3615 = _EVAL_682 & _EVAL_3673;
  assign _EVAL_2872 = _EVAL_3760 & _EVAL_2909;
  assign _EVAL_2150 = _EVAL_3812 & _EVAL_2474;
  assign _EVAL_99 = _EVAL_1782 & _EVAL_2671;
  assign _EVAL_1153 = _EVAL_1782 & _EVAL_3272;
  assign _EVAL_3453 = _EVAL_2743[430];
  assign _EVAL_2042 = _EVAL_596 & _EVAL_2474;
  assign _EVAL_220 = _EVAL_1782 & _EVAL_295;
  assign _EVAL_3399 = _EVAL_1449 & _EVAL_3670;
  assign _EVAL_1503 = _EVAL_114 & _EVAL_1856;
  assign _EVAL_145 = _EVAL_309 != 4'h0;
  assign _EVAL_1235 = _EVAL_1497 & _EVAL_1856;
  assign _EVAL_1113 = _EVAL_2305 & _EVAL_2909;
  assign _EVAL_59 = _EVAL_2401 & _EVAL_2474;
  assign TLMonitor_1__EVAL_4 = _EVAL_39;
  assign _EVAL_2348 = _EVAL_1391 & _EVAL_3391;
  assign _EVAL_537 = _EVAL_2352 & _EVAL_3673;
  assign _EVAL_1280 = _EVAL_682 & _EVAL_2909;
  assign _EVAL_185 = _EVAL_1892 & _EVAL_3391;
  assign _EVAL_3630 = _EVAL_1629 & _EVAL_1856;
  assign _EVAL_1948 = _EVAL_1061 != 15'h0;
  assign _EVAL_587 = _EVAL_2729 & _EVAL_2225;
  assign _EVAL_1819 = _EVAL_1961 & _EVAL_2474;
  assign _EVAL_3294 = _EVAL_1498 & _EVAL_3391;
  assign _EVAL_3257 = _EVAL_1782 & _EVAL_1695;
  assign _EVAL_1874 = _EVAL_2161 & _EVAL_3673;
  assign _EVAL_737 = _EVAL_2743[296];
  assign TLMonitor__EVAL_1 = _EVAL;
  assign _EVAL_1876 = _EVAL_2338 & _EVAL_3673;
  assign _EVAL_73 = _EVAL_3835 & _EVAL_2474;
  assign _EVAL_1439 = _EVAL_2762 & _EVAL_1856;
  assign _EVAL_1950 = _EVAL_1971 != 4'h0;
  assign _EVAL_860 = _EVAL_2743[470];
  assign _EVAL_1173 = _EVAL_2353 & _EVAL_3391;
  assign _EVAL_1970 = _EVAL_89 & _EVAL_2909;
  assign _EVAL_2806 = _EVAL_3726 & _EVAL_3673;
  assign _EVAL_955 = _EVAL_3523 & _EVAL_2909;
  assign _EVAL_3072 = _EVAL_3529 & _EVAL_2474;
  assign _EVAL_2708 = _EVAL_1951 & _EVAL_2909;
  assign _EVAL_2630 = _EVAL_3587 & _EVAL_2474;
  assign _EVAL_1106 = _EVAL_2396 & _EVAL_3391;
  assign _EVAL_2892 = _EVAL_2998 & _EVAL_3391;
  assign _EVAL_1741 = _EVAL_2028 & _EVAL_3673;
  always @(posedge _EVAL) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_661 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d2ed226)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1908 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16278090)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2898 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aed753ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3693 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4915705a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3767 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e727ef5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3808 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d1e6d16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3383 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f03ad585)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1908 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fc8b05f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50c258f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3344 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(601a88a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2278 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f378d0ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1534 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae219800)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3685 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94d143ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31bafece)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3446 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d64faec1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2109 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3f6e589)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1105 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b1ac503)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cef41338)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3584 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d00f1f7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2176 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18ecf1da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2859 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edb03d14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2258 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43090dfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1062 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc5b06c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3034 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2da89380)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1142 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69c3fc1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1604 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa77b8cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2405 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f716356a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_693 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcb0fb67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3082 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c38dab45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3110 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee2c0053)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2543 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6be4c2bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1453 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5725c169)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2436 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d683499)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_668 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fe6f9de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2907 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ff30c91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f521c099)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3667 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a6c8ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2394 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afe8d38c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2505 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7dcbe113)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_904 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8fcdfbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_810 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(285421cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2287 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e5a6332)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1584 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5b0ea0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3cf2b5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2184 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57f221ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2069 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4c3db99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2195 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d15a20b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1920 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(440ccf78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2205 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53193dee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_635 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e380e28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2189 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39733ffe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1683 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69dc5047)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79890528)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3375 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74b08141)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76cae664)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3693 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3d5e0b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2105 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(772758a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2030 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72fab1a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3765 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c758fab7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3153 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60c8f8f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2281 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(370f0fd2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2608 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c50bc70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1762 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ff4bc67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1074 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2c15944)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2107 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c509462)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2321 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9a34ede)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3773 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc467747)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3833 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e5df03e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3626 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c86fb4b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2690 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ede34785)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1505 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72a2c3ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1323 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bb74454)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3362 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f94108c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3622 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d2447e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3218 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48c49218)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1284 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e36371df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b386d515)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_831 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faac9c54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1924 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f37edaa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1482 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(923afab7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2331 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(218cfc26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_410 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(797bced6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1612 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22a2364f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1862 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c16aade5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_887 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32623653)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3205 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(603724bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3384 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c25065c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1768 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd39716b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2361 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(830d2d74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8aed861)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_923 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b12f899d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_894 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0abdd6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1688 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8129c218)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2000 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b53dcaff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1558 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a263f2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2335 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5d17aac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84ff05d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2930 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7852c708)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_687 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5646fda6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1434 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65d4d2ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a3ba6be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2950 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f24c9cf3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3264 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1efaa62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1396 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(562b7e29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3685 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74dc8eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2007 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fc851ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1907 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27e3298e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1775 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b5b5ad2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1763 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d1e0375)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3781 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f42e0fef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1214 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4272bcb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1504 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bb9367d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1338 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20a09ba4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1283 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(923c0996)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1049 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32fac9be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1889 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65aeb668)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1509 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fe040d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2523 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7100c2e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1820 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ad9b590)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1737 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_586 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(488a611)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1647 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10b84bc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2919 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2be872f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3548 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67b3789a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2606 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de93e0a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3136 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a159ae2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2556 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba79ad6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3260 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60d59a1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efc1b1b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1762 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7b5f53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2470 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f77e9fad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1005 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f31d9e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_500 & _EVAL_1730) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2582 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30030cf0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2608 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da55166c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1076 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa159f57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1739 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b95a05cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3253 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80e65368)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3053 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e4d9e9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1848 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d94068d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_446 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d8b99ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1504 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(336f1f5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1604 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2264fa65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2250 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f930c846)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2782 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f84ab731)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2189 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55a2b21f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1049 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(286dd099)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2112 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15ec5859)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1692 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f45e700)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2179 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac74cf6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1899 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f62540a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1451 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81a7ea77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3058 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f188cc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1434 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a1cf361)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3440 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edfd380d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1389 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ace3e18c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3243 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(249db102)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_574 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(553791b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2376 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(874d31c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3667 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c20f363)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2557 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a53e327)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1827 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44bbd901)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2088 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(499bef64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3400 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b22c5cf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27f57a65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2919 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f9992a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2171 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b344a1a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_924 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c584d00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2380 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bc02c7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27199d5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1416 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15f38142)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3439 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28b641a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1398 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ec8f706)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1999 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f14a5184)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3057 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94cc06c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3098 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff76f956)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1190 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0bf7740)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_665 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba67e20e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1371 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c4e40f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bfd1b4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2530 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d092b9aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(199ddf55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2824 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79454ee5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1289 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fe94915)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1141 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66067a21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1168 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e76b5f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2263 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45419b14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3554 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d00e14c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1712 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85efdef0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3505 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adb733c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_747 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f7a578e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2061 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69653ddd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1223 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe526d02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_600 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a14aa44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2071 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b8a9986)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c104532)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_986 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6a0e721)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1112 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6b8cb2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_724 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eeda8606)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1130 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e15280e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2181 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4a342d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69bb54e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3062 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc4fa9a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1584 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e12a2c05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2546 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fdc32a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1888 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b3f1379)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2507 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c5dcc77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2301 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1de137e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1406 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e41f034)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3130 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cd95a79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_981 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce4cc976)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2007 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbe6c76a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_918 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2512cf25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c626b58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1930 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aafbe2a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_672 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53c315f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1442 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40795063)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2917 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7145246e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2380 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(968f9825)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3636 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b04908e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3333 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7ac9266)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2924 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d636a0dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_632 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9e75c6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1617 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d3beecf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_905 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d42bb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1999 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1010464)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1063 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f493d17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2521 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fea9d23a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2348 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(288f7100)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_813 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e03ec398)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1810 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9aa153b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0d6047f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2824 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6edcd5a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2164 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92c176fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_904 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b0cc871)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2950 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(865aeb7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1588 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27fa59e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3828 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15fc6ccd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2651 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1faf3b4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1482 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fc3303b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1539 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5c41874)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8ba0464)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_641 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68ab1330)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_469 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f17b780)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_537 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2991db92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2976 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99af5f22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_369 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d2eee14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1841 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c038648e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1113 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a32bfa45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2931 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d9d9492)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecdeae69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3136 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75c00446)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3084 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab2dac91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3628 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd549325)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3346 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae2b9ff2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a5cd0ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1070 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bed335d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd5b34a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1879 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d6dc48d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2579 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fb4d758)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2835 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(912d8ce3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1280 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(368c2aad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2320 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dec278aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1885 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b95369e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c2d2c97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3060 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df0af0a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_491 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71916590)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3492 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(296c53bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1874 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c29dc58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f118de1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1854 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d8694d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1534 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5516a738)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2678 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e152cf8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_561 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f78bc2fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3628 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d86cb2a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2212 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5fcdf1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1025 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2208f41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5203b04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_556 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91320039)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2531 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ac5f027)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3617 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9c51683)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2400 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9af2409c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3805 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1ddf71c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_400 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23d81408)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1770 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93f2c3bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_341 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bbe4d57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2632 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66290cc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1717 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(476e2183)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1263 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a271bdc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2304 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6770e4d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2966 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a021a1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(372ee302)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_812 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12975a8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2860 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de8df35e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2187 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8154fa3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2863 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b56499c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_955 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(868a5438)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2142 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eeeac095)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3007 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54cdc503)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1485 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21713f2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3303 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94e9eeb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2109 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d76161fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b024ca0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1776 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(136c1122)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1947 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0983911)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3706 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c86e123e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e279fa6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_983 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1855e2de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_633 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad915e93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1676 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b0cdee8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3380 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43b0a421)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3721 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab338576)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1438 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f6c190f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2753 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d6808ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_581 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6253a7a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2327 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fe4a9e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1485 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd72811)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1416 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f8f7bec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3184 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53bb0664)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2523 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c010b467)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_807 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de059ee9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_917 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faf81e58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2374 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9778e839)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2796 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90a27898)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1385 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68e2113b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1829 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dde002c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1255 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1750 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6bcc3c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1387 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(852ce6a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e85cbed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1719 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d3fc8c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_466 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb23204f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2278 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa6c9438)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2252 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97edf677)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_970 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4eda693)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2889 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(871d7ab5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_806 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26859ebd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1827 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37499369)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2651 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a456ee1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1296 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5c1d626)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_703 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dcff9cb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2997 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6c38d24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_950 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d79a8fa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1816 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98e5215a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3605 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a10ebe4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3483 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(785e9622)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2273 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0f02cd9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2906 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(806dca9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2930 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a7a8738)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1499 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afdd5f29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_742 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c57b856)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3683 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3517313)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1673 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f5a7388)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2191 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e12488f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1028 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20afbfd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2038 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2369ab2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb763d9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1042 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bfc9319)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2845 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f087d24e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3796 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cc40d24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3617 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21505d66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a8f9055)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1184 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a05c477)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_335 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27f6992e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_698 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9faf9332)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1680 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(277496ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1741 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d66bd1ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d70de368)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1733 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(717e1c5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1874 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c075680c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_839 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9781e6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1621 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b178d7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2640 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d2ee7f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2585 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c98c9a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_348 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5ab0c80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2767 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d99c9c07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2405 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(facf7cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_358 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b502119)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3419 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3cc340)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_478 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb57e62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba7e736c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2946 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d3d8993)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2728 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7740aa3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1510 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a72bf482)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3034 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ba1f52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2832 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b572aef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_615 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e06da1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2297 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64bc632a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2778 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc9b3a8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1559 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf6ad315)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1415 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5f71a55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_593 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c799de2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3560 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e44f2c91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1797 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c3abfc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2208 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44afc13d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1834 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ea75109)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3607 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efdd0dd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3297 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd3bb686)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_954 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a9c37ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1884b4ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a02dd7e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2796 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d99f8a6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_318 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(686d2cf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3086 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(594e324c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_806 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(419881cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2583 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63647cac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1173 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d955cee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2612 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5890abfd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2393 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cc11ba6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1580 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b77c6a5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3556 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e309257e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_939 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0b300af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3796 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5846ad1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2993 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33398d75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2975 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c20333f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3037 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a83b0b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_924 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e052ba77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1946 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5585f399)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3324 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8037ad1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1316 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5c5aa11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2053 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2990 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e00b8fe3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2997 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab0b7e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1333 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3398942b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2023 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36e5c3f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2728 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8aac3c0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_416 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9f618f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1643 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a25d4886)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_341 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(670aed60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3519 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3366922b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2011 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec8b06f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fa36137)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42bec6fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1711 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9266617)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1373 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b016416)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1214 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4a068a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac639998)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2969 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ed469fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_902 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d130d78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_955 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5077e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a13ce7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2061 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8eb14e5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_557 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c86ebd3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3629 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76f7d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3314 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e57761f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_812 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50107deb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2155 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65fafc0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ec7d002)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3790 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f97b0349)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2200 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14109640)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_621 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b82e1108)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3611 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29bcf696)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1609 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31867662)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_591 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23b7baaa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1625 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7dc22f15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3222 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2e49466)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2098 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb64f2b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3367 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f45b41f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1079 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abedcb17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_581 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(303b6ee3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2971 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8366f0cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3374 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a28f50c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3240 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd2ce8ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1359 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec3dc6eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2645 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(250a3c96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3773 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2e759ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2754 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec1189a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_848 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e06e91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3655 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2261378)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2869 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76c58e8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3405 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ceccc119)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3575 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(932d15f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1862 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd8bb548)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1085 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56826251)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_773 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dcab0a98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_936 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2aec4935)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1870 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4f4c7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1836 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6627358f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_561 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96f20f0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_688 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1917660e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_529 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f9eb898)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3341 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4638e404)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1692 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce167e0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1523 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f0638f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3818 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98e892f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3386 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1c060f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2585 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce2b93fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3350 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6851d82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2362 & _EVAL_1730) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_629 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b13acc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2971 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f55217f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3790 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca4afcfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2072 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9de7cb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2764 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7422c5c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_385 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50304a12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3581 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd76c89d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1970 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(501aa11f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3455 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9765b794)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1559 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3221d74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1168 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e729d42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18598083)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bbf793d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3218 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47da72b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2131 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73a3f2f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3827 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a5e1d33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1088 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fb5fc9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1298 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4323bb6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3286 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63b8c319)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2644 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9eea4af4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1602 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc6c690)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3516 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea47eb2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1266 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fea4ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1811 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af4d7b68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2060 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d66b979d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca58fd05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2571 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47f1b9de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2010 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6178eaf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2408 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1303fad6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_359 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cbe3d94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1192 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8127d78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2426) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_864 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a101562a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2865 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2755bbc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1137 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cdefe04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3602 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c485e063)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1373 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f12f1ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1764 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf78ebb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3556 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68957c1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2876 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e478c93b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(548494a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_880 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edc436ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_971 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36338e54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3708 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfbd2ebb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3819 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19172043)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2032 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf480232)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1791 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b508331f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3180 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cde91c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_658 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f835f14c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2319 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f10c3039)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_884 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e129feb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1609 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(695ad193)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2292 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aec36b0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1364 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cd4f2a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2374 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b20573f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1595 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c698354)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1819 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6116042c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2010 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(657cb508)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2897 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(796d0894)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2309 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a393b55e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2556 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ea6356e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2632 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7194eb96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3405 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ae60cc4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1680 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f575a9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(897ff25c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1796 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9d1d34b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1002 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29d5f4a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1054 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8a77d39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3737 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1ed2b24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1924 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b1b371e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2884 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63ef459d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3501 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4eec1f54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1489 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b049f0fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3051 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5970934)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_791 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4836b1c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2450 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c1f1b8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3503 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b30c933)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3225 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f22cf5d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3386 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfcdea85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2289 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(496fb642)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3648 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bbd29f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1083 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c66f431)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_532 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(730241c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1361 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2b55de6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_433 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a143b42e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2108 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a62ef85c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1539 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19d6feff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1784 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53e50846)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(193ee034)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2903 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b79337)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(778bfebb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2377 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c8de7c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_761 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54a7da53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3626 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2562a73f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_494 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec07027)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2029 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74cf78f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfae3f4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2866 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67b04393)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2859 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(743b2698)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3278 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bca4497)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1463 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fda7b68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1664 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c691a0bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2644 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19522494)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1409 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e60060cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1726 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96d4cc2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2067 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39291646)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1291 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d7b4c75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27057bba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1222 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bf0b2ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1394 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27b7f303)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3546 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16c3e75a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3759 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7da92b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1293 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32474f98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1120 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(beb90d96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf0a6503)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3060 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3828089b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1191 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c410a270)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_845 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e50e3409)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2230 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99acec43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(770ede7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3478 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80618598)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3547 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91344635)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1949 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec27dfe4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_764 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c2738c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2082 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e493c08f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3202 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d05a11be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_589 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(699487e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_871 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(310c12f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(767204d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2232 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be03a944)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2924 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b413a8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2289 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80f5bfd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3037 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b6e3725)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a73c409f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2779 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be45205f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3335 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e083f1ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3205 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2a620c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6578824c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2381 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9b36374)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1768 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4af86d89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_829 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8b0ab00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2751 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(951b48dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae89edd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1134 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74b762b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3062 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0359bfd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3049 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c9f1abb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_615 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8160e6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2947 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f0715b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3479 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b130bf7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3721 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f97044f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2293 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36e51b8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3166 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4592b804)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3099 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4574955)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1287 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58265ee6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_747 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2115a5b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1752 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21cd900e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1315 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7048f65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1252 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e42ebaf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2509 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(841e4d65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1671 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c6bd0fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2672 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7f8597a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2806 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ad02190)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3550 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b1f6bb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1400 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3a58065)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3029 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35485a9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2195 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3afd552)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2535 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15c12314)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3699 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(608103f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f30c1c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_625 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e378ebb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1865 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1b733d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3341 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efe24b79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1320 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a94dc059)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3489 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd57736b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1233 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23dc048a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0f492bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3291 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47d13ec0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_852 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5b42932)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_632 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3e1f010)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2518 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1249facc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2549 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c704424)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1756 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be2f3b63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1744 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(684987aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3503 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a1b116b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_709 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bca6116)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce8fc42e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2906 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ecd896a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2446 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce174912)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4f08558)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3352 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6aa752b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1857 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f706036a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1595 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25b2647e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3158 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(819b5ce7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1563 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b73f4f6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1112 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce0b2364)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2337 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a471bf87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3797 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f72b61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3074 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2799c6a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_862 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(309fefe2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_761 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99381c11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_342 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea99d53b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1866 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fd1d445)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3346 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d051781)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_907 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27e9d0e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1676 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7938b751)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1055 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4990819)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3664 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a16c61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1876 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ae8b5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2369 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9489addd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3255 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86084e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_594 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c45c9589)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_483 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13a3972c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1673 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca9ad26a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3344 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4cd7c19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2798 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d889c17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1830 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e858dde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_387 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c317513)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1222 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f399a7ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2507 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e891190a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1302 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ac4dabe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_648 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2075f3f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1981 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(989fe799)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1072 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76c99811)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3364 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2cda2ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_755 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89500857)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1729 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9db334)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3126 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c688bb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80bcd4ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2891 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9c4a876)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_385 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbd5184b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_691 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(487d46f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_457 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfa45272)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2825 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a7c0337)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2652 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a13b221c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_388 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67c4ae3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61156cc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2832 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(551a2431)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1645 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74d77558)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_738 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37a8ad2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1589 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec8a645)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2062 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2b578d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1481 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae9b7924)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2669 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3307 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(770143d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_570 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c63dc7aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d30d120)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2669 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3601 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8307a869)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2904 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fce52149)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_428 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2df57d3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2797668)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3063 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc648fb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1298 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da46a8ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3210 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1c4fa9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2545 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(373560f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1976 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c95c9f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1286 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bcac078)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2708 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81fa1767)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_603 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dab6cbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_741 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(130fc79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2042 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49bcbcf6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3363 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e23b697)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3658 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5851579)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2179 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbc43327)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2557 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd5fb65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3789 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62531b5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2375 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d382160)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2946 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15475d9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2715 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12f8a8cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_621 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff959615)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_936 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7baca4f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3313 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94d8aaa4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1876 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ff80421)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2785 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3925536f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2866 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35b65ced)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2542 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c0d88b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3350 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c38c2c33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1579 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(508a6369)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1811 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa521e9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36aed0e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3036 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(352b8b9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1247 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24f1a311)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2564 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37df3fca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1346 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20eb02dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1711 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c3662a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c14ef92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_472 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(656106ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2356 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1dd9a27a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3488 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(941a813f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19952183)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_469 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6dbb04a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3305 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95f4346b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3801 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f96fc4ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3078 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41058a2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1105 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21d89ae2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1864 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d6e008b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_944 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(612f99c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4875e202)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3705 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97fc8f3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1916 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d5b831b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2182 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b50c9a2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1719 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(160ae5fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2511 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a944682)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2348 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1dc74fb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1459 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93ff502d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3354 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a29b4317)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3202 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(412d5f6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1996 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c19274b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1660 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bf4dc97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_691 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9f52c48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82537556)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3805 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2af4ad8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_834 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(151f869d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1335 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(186825c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1877 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67b538c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2032 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a73d66d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1a3d7d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0255ceb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2467 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3dfd3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2942 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b192772c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_845 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4636693)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1443 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5685f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_379 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dc5f206)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2513 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66a3f8c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3273 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d06a1f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2607 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35b2c21b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1308 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0145eff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1254 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31ea30ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_400 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9df7bb87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3268 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ff181c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2685 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6d4d908)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1146 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8eb1285)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1865 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8ff6395)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1698 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47d90ed7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1920 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9dce0c0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2546 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73f9eb93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_807 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4550a5e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2857 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1653997)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_677 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c12de8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_523 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a0c5756)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_557 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d92dc1e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(423d6809)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3622 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddedc3d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_889 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5361908)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2187 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa5af8e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2813 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb0932e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1745 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c938a4a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2536 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8751f624)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1565 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ccc26ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3471 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca8d8c89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb636356)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1643 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7df024d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3008 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30ce5bc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2723 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5fe62c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2603 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3de8d19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2212 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbdc9c3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a1fd0a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_531 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7680c878)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2148 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d75d6a79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3303 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c712625e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1990 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5d6bebe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_491 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67f81420)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ce771c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_834 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27c2f899)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3419 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e013e572)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_587 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc39fcb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3643 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d71033b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_600 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d091deed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2205 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdbe36e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2100 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(460dffc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1141 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8a4342c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2226 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13cc43ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2931 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18ab0a68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_918 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8c9298d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3489 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16b55b63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_814 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c13cdf4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1864 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c78e9ee9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3701 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52960974)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_460 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0e8b7c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2460 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5474dff2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3305 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(531f17c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2621 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f6e7827)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2963 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdb73cb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3635 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4358dba1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2319 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c951147)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2023 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4384160)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1777 & _EVAL_1922) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2510 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af10d672)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2652 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5713733)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2679 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2731c20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2087 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62758ba0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2828 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bcfb1fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3111 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70561433)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1554 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d4d2b99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_598 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8114b651)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2213 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f2d3a71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2916 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fea14db1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2009 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3588da78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_865 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f12b78a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2784 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f87bb2ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3330 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2056aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1784 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df404b9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1899 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eaf1c74a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3706 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b56c554b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1029 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd5d8b00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3627 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d845803)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3488 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d674e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_767 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7452378)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1810 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(583a6801)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2208 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a12270a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b5791e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1067 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f208d494)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_664 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28c54599)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1836 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29ac365b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1267 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78448c7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1499 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(641e2e8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_718 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20ea176e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_478 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57416448)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2594 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8256c6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3749 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a15d29cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1912 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a66b93da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1690 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61b95763)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1519 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(749a30f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1158 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b4cb6c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_416 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12be629)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1158 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ff85bdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1262 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1546a46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2940 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de0bdd4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3364 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cae4884e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2443 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98414d20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2357 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7a76aa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2065 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23bdac07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2172 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f5e7ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3075 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(198471c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2415 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7492cbca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2865 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(687b19a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1382 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d982bb72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1952 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97fd667)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2141 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d032709d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2914 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ba125db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_745 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58ccbd63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_889 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3b3002a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1458 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6036560)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dc19442)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_805 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45c55845)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3099 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(731c72e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1801 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f7d3c8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_938 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fc49cb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2892 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36882aa7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_379 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56fb17e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1589 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7091ff69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_782 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b184525f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2845 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ee22394)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3497 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b402ea4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1777 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84d1a44b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3412 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd8ae2d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2833 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a7ca9cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2967 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be3ba659)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2940 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c918729)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3340 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1bba605)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2645 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3147422)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3636 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae80979a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_528 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9faf227)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_871 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e9e57e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1236 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f6a0cfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_631 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(201eb9c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1024 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab4de2e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_501 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51eb4331)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2828 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61b65516)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_830 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99a728c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2752 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2bfc24b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1085 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f317ebb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2714 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(561cc668)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_520 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ec39a6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1996 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac2ce1e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_731 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(271bb41c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1080 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5003a959)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1183 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0d4286f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2574 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a218f9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1253 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb32f9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3505 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17d9cbdc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2129 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a2bc6c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_536 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0ce92a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3785 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(482353d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2726 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86ccb83f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1640 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d081a00d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2391 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be10fb32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_896 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e0710df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1909 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b1ed758)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2830 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dabb2bab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1704 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fa7f1c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2150 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7390040)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3058 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fe53a4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2561 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24bc65a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2053 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3708 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(777e55f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2288 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b99e3c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3057 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5ddbe8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2129 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1da69454)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3121 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44a49c42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2132 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffade156)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3451 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ae4ac83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3354 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5e97459)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_796 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6190f3e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1260 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1e56a80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3107 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(243bab96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2228 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e8ae3ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1802 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dad17268)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2943 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1c99f35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ff91fbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_983 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc24c446)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3107 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7509d952)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3611 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e040d937)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3615 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9409d90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1927 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c39f0e7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54aeae74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_791 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b48b9fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2747 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8278034)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2889 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(226d1123)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3716 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be9114cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1826 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(433d62b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1563 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a06795ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_755 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92120e49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3491 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b154382c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2767 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de43cac8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_874 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aea98d23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3655 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba8a936)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(420672bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3781 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0bdc33b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_899 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26572811)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2603 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89e91bdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1904 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc327d09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1463 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e33dd50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2574 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45e83603)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2230 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c24ced)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_865 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd6f4b77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3282 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b773ab4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1792 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afdfdf8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_944 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a713efa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3460 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a029f5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1446 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b245092)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2505 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(628afed0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38612a75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1515 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81efe7dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2483 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d2c819b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2413 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1480bb32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1162 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f20fe494)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9c6f12a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe4b61c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3301 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8730b40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_574 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28b6aac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(109144d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3304 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70d63efe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1652 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de815b2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1729 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac0443ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3392 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(999df00f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2542 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d7a39b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3274 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35a469af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2510 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f38daac6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2397 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6901fe95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1320 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19448d76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1412 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22a32d46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2142 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(691e9be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1640 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9dbbc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3455 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(affaa1cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(262bf3a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_687 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f21a277c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2133 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29ccd497)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1103 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a06345bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb1aec04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1624 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f56245bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3618 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb8d6149)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3415 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ab760b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3181 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(622be81e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3014 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68583246)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2297 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f04d1be6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_974 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57aab49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_827 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(472ac472)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3297 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a76ac413)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1280 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(935b20ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3378 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a439780e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_387 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c773b613)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3081 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53de1d8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecd506e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3732 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e16e35a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_627 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f76ee99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_810 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8d62bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1809 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0c6fa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1156 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4357a86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3765 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6d83c40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_640 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e93701e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2531 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a2a41d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2626 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe09d9f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_843 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c554c79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_945 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92743836)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3462 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba1bd67c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1236 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d03b6fa1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_525 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(902fb581)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_474 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54cadac3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2473 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c785105c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2891 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(615bd422)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1707 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7769e534)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_901 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c02e116c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2085 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f29c4851)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2502 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52b08852)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3156 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5cfb3a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3656 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(866929d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1829 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c7b6546)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5099fad4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2876 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d2eebaf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1120 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22b46dfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1406 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdd4f858)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_586 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(153e04eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_937 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9478850)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1029 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97e77a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1814 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d80e8b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_460 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c20a2aed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2252 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8787cb34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3300 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(feda58d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2473 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3d69964)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_388 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a9e6b0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2562 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99bfd0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3117 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(490c65ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2323 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afa3dc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3467 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fdc0b6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_741 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12f095b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3407 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ec82f31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1885 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7887d23f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1909 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6ca2d13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_520 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c5e8d02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3720 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ccc8331)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_588 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83de0a98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1107 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a8c1eb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_570 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4be9146a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2617 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a511d5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3563 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68ba608f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3222 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13638104)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1912 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbf3e580)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3384 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ae79d81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2153 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81b2b523)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2670 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecccfca3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8da67a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3028 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1f6da2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2141 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30ab569c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3701 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6910db98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1113 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b64e8174)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d068af1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73e6aa9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1854 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4edd3149)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1173 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89766c55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2916 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27e1b1fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1647 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1788f82f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1501 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2354e9f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1649 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68bd219f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2521 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(376d0587)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2386 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(947c2ea7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2999ecb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11a43526)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1178 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1752e2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_782 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dab363b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3188 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a62dc0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2250 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65a5b88a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3131 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8e94717)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_428 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ce5ef86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2857 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfc11939)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3086 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(866f280f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_898 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3e3ee6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2620 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be773e85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2973 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e403c23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3374 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcbca3e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3692 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e6b421d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1645 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faf29278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2567 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4398d651)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_380 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e75e2d99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2620 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2242756)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_954 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6515c8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3578 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20334ada)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_629 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52209348)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_537 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b7e5a97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2680 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4350e550)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1756 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39fea934)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_978 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58faf6b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1028 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8eb490c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1610 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(157c9ef4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1906 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3f45038)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2221 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bca2a0fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2461 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0889e22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1431 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f85a41b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2860 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a30bf0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3108 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cce302fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3192 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdf38c10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1820 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23f33dcb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1668 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1b58b84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3749 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55b0125e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2152 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78ba4bed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3463 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2dde3c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1712 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98328e09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3362 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae1fc7c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2773 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(552d72c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2640 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15654495)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_531 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2436b8d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be09f90f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2436 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cba072b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3615 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dc8b086)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3818 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4a14f9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1565 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7259ed78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3441 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bae761fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3514 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5348c652)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_811 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73dbcba3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1952 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d904c5ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_926 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d88d81b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d23f011d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1171 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(808814e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3208 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cc12708)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2778 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(946ce571)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3199960)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa345cb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_938 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(384bf0cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_422 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9478285)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1453 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59760e58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_901 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e10aff9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_829 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a584346)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_631 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d484cae3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3243 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56d1d908)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1668 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23eaca43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3646 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99a1e0db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1369 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62a03c17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1248 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee6a5dce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2528 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cab1211a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1265 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa8facc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1605 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8077631)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_593 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(495881c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77a690b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1651 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(181dbce0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3575 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73eeae4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1310 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73e2b1d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1555 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79a2d7e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2391 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d337a4dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2626 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f1bf115)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_729 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1859bda4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1063 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b38a51c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3253 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b98ce50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2867 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4ced0b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_939 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e30f6233)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1415 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(510fd8dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2612 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3369fd49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1848 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(499a5a4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1199 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f001fa7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1092 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31c53a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1259 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(230a37a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3434 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33ffd897)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1554 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f59e45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3792 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b0c7566)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3692 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19f513e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1359 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7925203)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3311 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e0c2e2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_945 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b9703e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_989 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dea0e9c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1248 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b3d44ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1871 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c51c64c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1670 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(243bea88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2049 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11842a8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41bd5ace)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2579 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75f39e36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe09de9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a663fbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2806 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a000ace)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2875 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2cb9be7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2577 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8e361c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1600 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d02e8327)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1704 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(533f582d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_853 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9516b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2779 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3dfcfadc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2783 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8254daae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1816 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b690e96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_594 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd80513e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_811 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49459e4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2630 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4217ee2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1988 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8750597e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2658 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(739b3828)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_816 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c76007b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3616 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(293a3bb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1376 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32f80d74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1918 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0d183a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_756 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(543de5b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_408 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cab60510)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2242 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7af3b9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a60fed7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_523 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11dfd0e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1817 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17b00b2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2242 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ac8c4a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1739 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da35a1b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3565 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72dfadbc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b160230b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2172 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85f4572)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6948abfd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1537 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c483bec0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2394 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6072eced)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3624 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92c350ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1826 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f2b7bc7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1519 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b73abf91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2375 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faf2e20c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3181 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db700be7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3627 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6e53086)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2313 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fee2754)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_664 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f55de14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1775 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8f5cc7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1753 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(770d948e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_940 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c76108e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_422 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2c5aa1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1247 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a24c7f46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_733 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b139d021)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3296 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8aa6d1c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2988 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4ce3766)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_483 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(703622fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3300 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3f7dea6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1558 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3ddce7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_804 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea84777f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2776 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f73cfb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2753 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32d8e4ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2044 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fef622e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2678 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11a8856b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_796 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(668f2817)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3737 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b3611)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1338 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bd700c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3563 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d5bb0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1792 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(440f6dcc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2443 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e68ddb44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2617 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(673b1927)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_515 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58a6c333)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1202 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b85412aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2067 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(148e4bcc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_856 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be6ad680)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1776 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58d7fc67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1830 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bda7d86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a15072)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1134 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b739910)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_805 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7b91c4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2625 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f68a8d1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3092 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dec3ce9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3324 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(847c2b4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_952 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2375ee4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1344 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab8194aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1651 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22d15731)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2942 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdff80e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3077 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1963451)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7225a23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3166 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92805d40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1698 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e8a3e77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3756 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(500d6bbf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2868 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ee22b0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2914 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8c432a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7baa962a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b103ec43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_903 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef964612)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3110 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b0060db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2221 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3821e66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2065 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b0920f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1253 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7605eeed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2036 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f12c89d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1828 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f05504e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_597 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(147b0fb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_380 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79cd031f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_588 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7106071)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2530 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3ec0433)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2751 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c9b821d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2596 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50f62748)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_743 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7465454)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1239 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(312fa7b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2681 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3883f66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1f0838c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1709 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d46b5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1382 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e9630f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_701 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50c937cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2773 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90ab3354)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_838 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(860e09dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3445 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d79f75e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_935 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95dda68b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1254 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f205ce8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee2ba7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3313 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87886d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3082 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47c59f15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_880 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47217df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1841 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e48b409)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_625 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5abd6281)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2416 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(727e688b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_838 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(560df173)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3507 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a01d4e32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1279 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64a0e864)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_666 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2da6fbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1417 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1eba6fba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2800 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8594a34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3572 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a66afd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3063 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8bb0ef5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2009 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62001e8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_525 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b154e66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1828 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9c6f467)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3336 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdbe0390)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84808e25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e0aa833)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2335 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb489339)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2903 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc270869)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3440 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(303542c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3747 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(492e6137)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1857 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcbf451f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2782 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb4ee3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2469 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6abec1b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1446 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d28b0511)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2764 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1dff7678)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1070 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3e66acf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2621 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b97b4562)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3125 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60780f1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1346 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd21744f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3375 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d96d4bb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3074 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33d7d4bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2287 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db2881b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1707 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b10a09f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1431 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc3a0266)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_335 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2467c02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1336 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53e601f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1800 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f779022)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1239 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(143b1fad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_903 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a257a9d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_465 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9024630)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1906 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54d047fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3528 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba7bb8d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_927 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82baef6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2529 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e886c86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_729 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(340a0251)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca027ea7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1901 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(945213dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3378 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7196f20e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2454 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(680b5ddc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3547 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26c9d7da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2152 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a46fd9c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1757 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b8cb2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2902 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85cf3180)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_742 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8031af91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3578 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e420c35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_986 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ffb3db1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3296 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee1546c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2036 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecfc032c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2060 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76926804)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1191 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c957d51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1523 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2defe946)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3256 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19c6fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_905 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c2084fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2715 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31a58cad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_853 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a529e0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1190 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71e904ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_472 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(784a76c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5887efa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3153 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4149f647)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_894 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e0dcaf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1263 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af93b28a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1310 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ff67fdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1005 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ef6bb77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3580 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a183dcff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1916 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10e06b55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38ba80a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1103 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6bb3241)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b75f240c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1308 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bc6cd1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1473 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4164b08a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2638 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78b5207d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3273 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b15a15f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3585 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c7bb004)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1580 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee5d5862)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_437 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26a8bf3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3263 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7eba4e11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2098 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ec5ed2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_887 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87068765)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2072 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b388c564)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_462 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ae7c68a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b4d1f93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3282 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24935eb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3680 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(334fbc4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3294 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be1873a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1473 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e001d5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1249 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cc58a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3699 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cd22de1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1438 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc0488d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_694 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7b9964e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1621 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d503a556)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_410 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1301430)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2577 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12879dfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1946bf99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfee2886)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3192 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a284144e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1800 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bebe8bdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3585 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4797f61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2563 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35d70f0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1502 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa77b7b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1442 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ba1ec06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3697 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69444d84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3792 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a9fc32f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3543 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(104c9f46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2416 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(652a87c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2907 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c4c7f37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2244 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(938c7ee3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3588 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(410bb0cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1501 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64c36be6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3383 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(803bf739)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3910e249)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3580 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(862aa961)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1361 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c050b72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1146 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17074eb1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_635 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10f02eb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1797 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5223d26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2062 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aef7fd50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3560 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa9d8c01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2192 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31f71cfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3036 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bace7b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_641 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1afdc421)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1753 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2da26920)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_474 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c08690da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2766 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cab32e74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d963ded4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3789 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9415cfab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3225 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8b47bb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1464 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24b04c27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1750 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(923b3205)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3646 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dc3e20d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8526c02f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c3d0edc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3766 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(968298c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_803 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20ba85f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_462 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(967b302d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3584 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c09c2ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2830 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6fd3afa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3208 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7310fdfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2596 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(483c709e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2714 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36885b4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2571 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9fffb12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3084 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4dc6b839)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2599 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4cd7817)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2606 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85e4eb2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3656 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccfe61f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3715 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b679912)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_703 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e57be1b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3098 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62b66486)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3516 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91b318bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1573 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ed5c7fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1281 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de4327f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1852 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(612a6481)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1949 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(134b957e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2170 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(882530ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3307 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c87cbed3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_718 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14870494)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_883 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c94ae42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3400 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fcf69dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1661 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cff57bb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_433 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f95b196c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3441 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(472ad81d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2670 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1844e37c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1521 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e44b604)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1364 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b45f1b2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3725a46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1502 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff4683a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3808 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8020a225)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2535 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb310e54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1033 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18d98054)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2341 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72d6e6c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a90f2f10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3392 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(611b54a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2301 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41970d10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1764 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6a0dd1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1522 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e55e3b10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3660 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cae58633)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1705 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d303a0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3199 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cdab695)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2329 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e193dfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2381 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b2ffa59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3008 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aaf58497)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_364 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0693a19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3072 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cc0005)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22faab85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2679 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0b077cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1602 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60fbd9a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2069 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b304a974)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_666 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7b7af5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_573 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e504243)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2038 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a01243a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5080183f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2397 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(811a5c36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3311 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(694df4ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3546 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d60ee58a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1976 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1e50e70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5867dbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1879 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fd0d92e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_677 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cf24fb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3581 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdc6dcba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3381 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7839bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_733 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10eba8f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_745 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db11ed70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2309 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a55a470)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_501 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31b11b44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1997 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62a07776)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1055 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebf70cf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1943 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa5d8f56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3463 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8372579)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2400 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bae97e84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2567 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5c62ac2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1058 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9458cad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2082 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bb25736)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1001 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99b5fd40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3491 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84a95361)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1904 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d1ebe3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1619 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b35e234)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3559 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86c1de5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1260 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6ac4ee6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1819 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78b31c1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3715 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b492d29a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1296 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c400b606)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1062 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faeb3247)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1535 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c099d58f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_824 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19ca667e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1619 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4990d237)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3363 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c269d72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3294 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abd7ef29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1306 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cbb2a04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2502 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44d36841)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_856 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(989eea69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1573 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69e7bc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_981 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f9ec9be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_893 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c7e8783)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1981 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5a68e86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3330 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f8168c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_776 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ef3555f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3827 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fff0769)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1088 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f86c4292)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3081 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ace7bcb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_898 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc6611a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3255 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b1dc147)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1781 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87b64c12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1156 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d714881c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3439 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed5dc9b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_468 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a15e111d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2100 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b78c261)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_446 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ac2cc7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3483 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3628d3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3355 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eeca2891)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_970 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da63596c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3801 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f44508a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(334d2a0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3352 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ceda0e63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1394 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9b9d6cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2243 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49f1bcf9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1288 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7595a158)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_468 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8f6bab2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_892 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b2e2dfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2266 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17a610b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a3b2ea8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2646 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cad97f3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7c00d68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1129 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(180ce570)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3010 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4eb45a9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1229 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5abece8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1288 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac13a48d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f114ea81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1335 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d4c3b8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_648 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e26f65cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3334 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37fe75db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1926 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d68a64d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1002 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(867393f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3797 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c72dc55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2808 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdd61ed3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2872 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1378fb98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a16ec612)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_609 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ea0872e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b73abc77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_589 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f46a9a5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_457 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c52f3955)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_715 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a69cc705)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1371 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d594efc7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_494 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e52a959b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1946 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cecd49d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2454 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23267608)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2094 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82ffb2ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_824 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c2bb1be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3415 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc3a0007)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3643 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65493db6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3413 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5de4d92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3766 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e61f8f54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2601 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9451721)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_714 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df6cc4ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2549 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a71170a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2868 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b26b5abc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1752 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9db8f36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1926 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ae39b16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3747 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae5f762e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3139 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9afb9dd8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2320 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bbd53ebf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_978 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d808e15c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1289 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5091a394)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_490 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31210fb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2018 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f68041a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3631 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb63bb19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1400 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63e7b45b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1674 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cbd0689)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_373 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97457575)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_975 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f46bee16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2638 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(450aa663)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52726fa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1129 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c3954d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_813 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5bc92af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(582e26f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_800 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6b3c4d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1330 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac9effd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_627 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2577b16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3631 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98bc91e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1459 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2532b587)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2969 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b2d51e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1509 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cafa23d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_756 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d478f1f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82635c23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1761 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cda5b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_318 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c203e00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1202 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e23e31b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1245 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(778c35ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1801 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15584f41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1930 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27137c90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3314 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45acf743)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2516 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e93f05a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13b43ef1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2258 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc7521fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2409 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c35f686c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_381 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d36319d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3683 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dd6013d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1781 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d2e29a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_408 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53fbfb9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1683 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a568c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2105 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb43cc78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d943a9f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_950 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b5fd476)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3044 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fac26edc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3550 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5c6e9c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3582 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbfd2cab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2415 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6580b35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3355 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5731812c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2825 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c2eacc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_974 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfad5dad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2269 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f0ff4f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3756 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8985dcc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3659 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60484e80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2346 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab90ed8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1970 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2b4f648)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_892 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9312f68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2304 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe9d34cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2562 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90cf830c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_424 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c712d921)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1616 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac55230c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_893 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cb35557)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3158 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f6d5ec7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15201c40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2702 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87742526)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_694 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faf54c49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_896 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43f0b71d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2108 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0a47e00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3525 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9d90491)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3548 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(324d7257)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1106 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ab8678a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1870 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a378cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1888 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2d64594)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3336 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e3d531f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2176 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f58336c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1225 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac6e2466)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1376 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9349608)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1117 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fbae3a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_429 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f3cbf89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efddee06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3075 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac392006)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2681 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94d6d02a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2805 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9731d4f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2646 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dee59386)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3049 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad15831a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2327 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e35ce095)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2563 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99f18db5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3139 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ba0e288)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1509abcd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97119a97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3274 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2fd21c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1001 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19f3920f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_358 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e682a6b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2049 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b1ef80f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1733 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dbf14d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1579 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eac933d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1817 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d147ab0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_348 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20ce7f4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1106 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(229f9c2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3029 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36d2fdd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3538 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5d35729)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2460 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e6ba775)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_573 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bebd59c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_515 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0857a57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2513 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3ea7107)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1179 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce505542)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2511 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58fcf79d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2658 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5c8168e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db917cd8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1664 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(626bdc73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2509 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e3645d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2803 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(368749cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1203 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(277dc68b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1709 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6747852)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_364 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f92f31db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3007 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(494506a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1791 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aaa8c250)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1555 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8113d00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2900 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(857b084)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3111 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8528db53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_562 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d36703af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1279 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b3aff74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1670 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46b4a82d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1575 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b70e74c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfe106c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2313 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(141cd003)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2164 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efe2d47a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2209 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b90d73f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1997 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44f1ec48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2572 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b467e359)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3713 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(657aebf3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2844 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ad7fc52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3397 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30b6d2f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_816 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc8f19cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_731 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cab898ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2993 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93a7a5c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_556 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1629c3db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3077 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc92bb68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3759 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15e38c3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3660 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70392c80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1396 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8037ac6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3497 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4c7c0d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2148 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80e78a98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef18a541)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_937 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3521f415)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(678d6cf0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1409 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(281e38db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2292 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b954f72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_884 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e7a7a17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_661 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bc5dc9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2599 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2669166)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1245 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cc84ddd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3588 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edd815c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3353 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(999e70bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_831 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6eec7113)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_827 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d5d81ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2182 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a89d7060)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2150 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79627fad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_971 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(559343bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2444 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ded3707)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1624 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8debcd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59e6b1fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_598 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7a276e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3197 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(182afb9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2723 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e978e135)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3191 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb072615)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3486 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd4184d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2013 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bc73d1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1074 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77bbad88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3460 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdae4aee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3785 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89cbff9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_899 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb516f1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3554 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e0f5dac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2990 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d93c6c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1162 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62a657a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b4b4109)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1336 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98f5d17a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_373 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f0c7d2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50c28c88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1763 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38392a61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2393 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(816c25d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2350 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b53bcf0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2263 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f1db204)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3618 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(637c029e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2170 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40eb6145)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2281 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5423da3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1526 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d013a88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_839 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a06693a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1809 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5adb6cfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_429 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c9aa69f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2131 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e037548)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1761 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c4e3350)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3467 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61474fd2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_709 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(518028e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1389 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a2a643a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2902 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db8d9b4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3582 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31ec9ce6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1042 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5bcc688)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1735 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a6b610b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2601 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(914c693b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2833 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a700b03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2361 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93ee2987)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1923 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bec93b66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2747 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(feb7fb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4247502f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3367 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd6b5dcf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_698 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d139da9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1058 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ecd44cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1072 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a1e6625)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64c48a63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1199 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(529f3b72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d47ff688)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2983 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba98c569)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_701 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f35889c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_456 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95e11b97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_688 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52c4459a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3514 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb575f5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2904 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c3923b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2244 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1949b8f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2625 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8c2c098)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_848 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3b6af17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_693 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b5e51bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3072 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e2594b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_394 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e38e1cda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1344 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45cd8370)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_633 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a92f46b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1858 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cb99ed2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_975 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d5a1441)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3625 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7993ce1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_902 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(779c73b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2446 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cb93956)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3525 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ded8a78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_917 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8820b5eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2462 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(313b36e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2543 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f567a14c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2813 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0039e63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3199 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc092ff9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2213 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(668d46c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1291 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15c2a1e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3559 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(421f5ab5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3462 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae4ac25a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2898 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ace39fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_787 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25b754c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2561 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94ea2aa1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_424 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8431c5f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2784 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f40834c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2461 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4a5f14e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1458 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb0ac790)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3191 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(884b1c0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3180 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b81d729)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1757 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa0f62bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2975 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3684cd36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3446 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(922dd204)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1932 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e57f5d00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_843 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96fd525a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_405 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36621084)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2892 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d980bdef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_830 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b89cf5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2273 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70bb3c81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3478 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b266c81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3335 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1cbbf76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3044 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3adec6f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2337 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(681b2952)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3242 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(469d33a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3732 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c74ccfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2798 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1eebd29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1660 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bbb983f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2900 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4d0c33d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2754 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f9dbe54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3108 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8bd5af2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2151 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16dae96f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1464 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93c43e3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2329 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f194b16a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1192 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8466c4a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1225 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(409ca0e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2266 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89a940b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3340 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66ff8f95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1302 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c7c28b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3601 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64e29c6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2441 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cce31ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c88654e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1605 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0e80ec5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1266 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a595ddb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2808 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fc87c86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2785 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c97e890)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1183 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1837effb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10bc5c63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1316 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4d9a999)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2159 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f51511cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2184 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d17051ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2357 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d76e1a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_532 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c143353c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2147 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(657caef9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2450 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71a86b62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1600 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c1384c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3260 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(878eb0ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3607 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98d73684)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3572 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa1354dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2844 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46fa6c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1636 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab68b6f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1741 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(484abc8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc05f8d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_814 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(216566e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d57c2ff3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3051 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86c774ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1184 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(675fa836)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3184 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fc9c311)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1521 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a83f8f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1137 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12ccfff4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3702 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ef0b9b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1451 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17864147)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_864 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(745e4bfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1907 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1ee946f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3333 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c3ed7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3538 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(606b3a41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7afc0ddb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2171 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9444477)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1481 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dc8ba9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3570 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d1488b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1770 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ece1800f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1663 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ef93ee2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2132 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a036263)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1866 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70c56b53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2042 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(926603)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2814 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4db1a39b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8623269c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2766 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2682864)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1107 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea5d20b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_500 & _EVAL_1730) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4bd5a2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_639 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b959b7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1f5becd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1412 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0772689)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2966 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5c60a02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2587 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4d38b17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1674 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cff4b398)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3131 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(593ff74e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1229 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b051334)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2867 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2c05eaa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2594 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8f7701b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3301 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22537e65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2630 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ba23103)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3397 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(229afbe2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1427 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb4dee75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3552 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18591578)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3092 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9956e3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3697 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc28c95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1858 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3da92e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2467 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7145b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1943 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18d8a01d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_786 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(226f505b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1092 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a199112)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c7ac584)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1315 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42f72480)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1515 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf99cf1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_342 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(258929b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3664 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cdad874)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_928 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3015fc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2293 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6232689b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3028 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39366c59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2181 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(906c1e7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2434 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1ebf760)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1080 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d26e24ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3078 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e737419)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2976 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0808006)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76b2dae6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3716 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea3e733a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3010 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a205ab3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3197 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c90696b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2088 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13dfd71f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_562 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9014bbe2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2153 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95389fd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1130 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afda2fb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_775 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d87aada1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2872 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16d28d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1608 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9712a4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1286 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f2bfe4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_591 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c22e0af3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_926 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e3c2607)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1281 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e748c3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1025 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4435aad1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1369 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(630056c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1617 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7a8aeee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2030 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d7fc53e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1749 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5681c0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1901 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da3234a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1929 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6d2c782)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2536 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d9b9cd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1671 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(723952ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_369 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5c46be8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1663 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d86a2e7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3126 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dcf9e87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1333 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abf14699)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2583 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be46864b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(feaf6ae4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2239 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44c56458)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_663 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8c07d7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2752 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7e21385)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2232 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9485a23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3501 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19f2ef62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2607 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(393f8e0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3659 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99907baf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1255 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_976 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37127841)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1717 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be4e278b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(979aa45c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3648 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c1cfec1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_597 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(795b7e43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1252 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f62bd8a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2441 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(363dbd8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1323 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9192f3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1223 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f216258c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2331 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f22dbbc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1203 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1393a86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15773e43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3629 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ed60ac3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eca28028)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_935 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fcd802d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_465 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64e14390)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2029 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a258ed9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31d4fe34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2518 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9f67acf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_907 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb3c36bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1575 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(692cc939)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_724 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9e2a275)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1249 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18e1c957)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3605 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddfce2b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3451 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfdd49f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2200 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3413cd2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_529 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e04fdd72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3528 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60aa8fc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3263 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92eb14b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7fa30cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1649 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b38fe11d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3380 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bf12f89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6bdd99e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2346 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd3cd946)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_668 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87da572d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3188 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b446b380)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3833 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcf6cb4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2426) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e3eb251)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_665 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1d2ae0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6826adac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1233 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99df2de8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2243 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(625bfbbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1947 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3df4ca34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2805 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(781d35d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3215 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae9d7a0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1492 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d19840)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3264 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ee616c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1522 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2072b56b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1652 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea0dd17d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1083 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1dc03845)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2356 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6aa39f7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3053 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b55691a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2917 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c4c070a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3414 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7f4fc1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3819 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40303ca4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1067 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a133f9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2800 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ffdc986)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_776 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58fad2bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1744 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1219f5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3752 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5e6d395)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2680 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35019389)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2191 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f68a5c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2070 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cf66b12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2070 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(509d0499)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2408 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e6636dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2469 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(872c187)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_644 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d7ab9ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_775 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5603ef21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3680 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(409b5a68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1259 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8bd7438)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1802 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2ab61e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_786 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(292998ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1293 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(459d85c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3767 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c2f58eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_714 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc0bc527)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2564 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5afdcfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3828 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63614f8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2988 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ceb836b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1923 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d72dad6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1024 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab3cfcb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2783 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c33961b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1726 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f4b1452)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1932 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38d4d89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3117 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26ece127)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1929 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6112d66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3519 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(145ae8f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_435 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(875545)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1330 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5520e55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1306 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a913078c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14aebbb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b1015fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2409 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b8aa5a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3713 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ded1e8a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2209 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91a19ca0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3268 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7e000e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1877 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65567545)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3635 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36dfed16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2923 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56853e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_852 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db8b75a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1144 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcc9128f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7762bdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_976 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd27aed0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2288 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9769cd7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1834 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af55ceb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1427 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8a824fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2107 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b217b633)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3407 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(655996eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3125 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c56f849)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1267 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0ed17e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3705 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8de751b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2000 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83e20d98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2112 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18a4c095)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_490 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d479d020)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14f44682)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3277 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2acc251)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ace57377)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1918 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb319d6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3056 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35d99639)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2835 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c31558e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9892eb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_767 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(250bea59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1505 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7998ba94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10a220d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_381 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1db18417)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31be34aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_423 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afdfaa2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_394 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47040aa6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b34db3a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1117 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86a93d6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3256 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7299f588)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1535 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(387146a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2545 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(311a39c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_927 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bcd9e4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2362 & _EVAL_1730) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8ee57e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2582 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81a41873)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2726 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(910d00c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1142 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d0cc8b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1171 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d09e4c56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1852 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(963e4882)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2967 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af51e8b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1625 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62a2649c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2814 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1882046)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2147 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8d7ef8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_456 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f86d46d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8043f47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1385 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89fec70b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3210 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e842776)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3702 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(622a1cc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_803 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5a7d110)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1054 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d010fb1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1492 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b48e4122)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2690 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c881ac4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1745 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aff1e475)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1688 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fe6770e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_609 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57b224fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c3252ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3291 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45498e52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1796 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35210c29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_435 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d634ef2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1510 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d5f5b14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2386 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6227c2ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_874 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(534ff1af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3565 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f4b7fe2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3492 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86e7f76f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3471 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d76c69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3752 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c3a4f2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1988 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64e34c5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2155 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f86b5dd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2085 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9fa204)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2018 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47386e8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2133 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfdfac55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3353 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edf755f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_466 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3166213)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3401 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f661118c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_359 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bf95876)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3625 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a319c968)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2529 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b5b7198)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3163 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54400db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1608 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f57d66ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2071 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7869443)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1990 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7707627)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3658 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0eb84db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2776 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8b2e337)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_658 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5fcbfcd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2897 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e60b6e3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2226 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6ad1674)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_437 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5e2a831)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3286 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(719a0eba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_743 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a218ee65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3381 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70ec09e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2434 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(decfc35b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1588 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7ff044e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3552 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e9f142c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2239 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(273571b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2228 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a0378c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f8b0be6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1179 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e63291d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2943 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9c8d89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1079 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e53eed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_883 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbca5b81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1387 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad01c88e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_800 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(358a9f57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2672 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(caba51cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e35c7f1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2708 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea33e0f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_940 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3262bd45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_989 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc236e28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2044 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95e2d106)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1612 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3999c026)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_928 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(475fda88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_536 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b492e19b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1287 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(835e2d43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_640 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(577fd45a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3304 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de094b25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_952 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56d00af1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1927 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dce8c916)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_787 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78e6f278)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2269 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e650509b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3215 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(521b177d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1033 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0c34aab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2192 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b37fe7f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2875 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(326fe536)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3570 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25d223c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1fcfba6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2516 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(449e561c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5ae2d36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2094 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92518c3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2350 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ca0d8b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2963 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b373753c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_603 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3e27bba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2973 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93d1955b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_663 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e61a9a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3507 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c2791ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3401 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0b6ec3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1705 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a8680bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2341 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f2f5bc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2884 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18d3db35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3242 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bbb3fbc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_715 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4578269)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3486 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28471ecd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2470 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(439873da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2151 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d2f7150)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2863 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba4f998a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2087 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16445682)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2376 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d84ddd3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3277 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a6eb67c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_804 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5cca852)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3434 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87ea4c78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3211 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d87cc71a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1737 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_405 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8cb8d99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1537 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92164e26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b1253c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_862 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76c7571)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3624 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ab4e09b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2462 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b9b00fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1636 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e1456d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1610 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(540b02e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2685 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b31b911)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1690 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5aa77553)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2413 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a72b76ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_738 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3bc4965)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1489 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71463160)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1398 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24f01336)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3121 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(967d91b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2377 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d096dea6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a0fcce7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1284 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39f3d622)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3445 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8fd53a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2013 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(418e8007)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1178 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5f38bd2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3156 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8779ed7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3130 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aaa2e7c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2803 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(387ed6a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1443 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fd161f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1889 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f328640c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2587 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85716c3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2323 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78663546)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1632 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7ab264)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3240 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7fb5907)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3056 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ed39a0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3720 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b97e95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1526 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d879f1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2483 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23f4a47f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1632 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41877cbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3014 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(345a85a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2011 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5080f941)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3602 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27769747)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1749 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bc7da1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_773 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ece0df9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1814 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97bc7208)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1871 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f107a2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3479 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3bfc9ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2321 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fed948c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2702 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a072a66b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3543 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4152dbdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3334 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e57194c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3163 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6df09a90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2869 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a42784c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_923 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6f1d58e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_764 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(917c3b45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2923 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4fb5419)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2572 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60b7c481)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2947 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a009a68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3413 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(738fb6cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1616 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5c4a7ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4607652d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2528 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79481c8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1283 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98b2a2ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c602b5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_644 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bc6b96a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2983 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1519266)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1076 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d02a595)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3278 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef8a1f90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3412 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa359124)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3211 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7dd9d5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5edadd4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_672 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c25ebc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1661 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a79a1d27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1144 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87f8c664)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3616 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27361248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1735 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d42ccc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8034232b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1262 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3bdc177)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2159 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39439aba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1265 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38f114e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2369 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd2819e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_528 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(525d1f86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3414 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc8234e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1417 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e79a1060)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2444 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e07424c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_1922) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ecc7916)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
