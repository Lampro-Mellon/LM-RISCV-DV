//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_6(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  output        _EVAL_3,
  output        _EVAL_4,
  input         _EVAL_5,
  output [31:0] _EVAL_6,
  output        _EVAL_7,
  output        _EVAL_8,
  output        _EVAL_9,
  input  [31:0] _EVAL_10,
  output        _EVAL_11,
  input         _EVAL_12,
  input  [31:0] _EVAL_13,
  output        _EVAL_14,
  output        _EVAL_15,
  input         _EVAL_16,
  input  [1:0]  _EVAL_17,
  input         _EVAL_18,
  output        _EVAL_19,
  output [31:0] _EVAL_20,
  output        _EVAL_21,
  output        _EVAL_22,
  output        _EVAL_23,
  output [3:0]  _EVAL_24,
  input         _EVAL_25,
  output [31:0] _EVAL_26,
  output [3:0]  _EVAL_27,
  output        _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  output [1:0]  _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_34,
  output [3:0]  _EVAL_35,
  output [2:0]  _EVAL_36,
  input  [3:0]  _EVAL_37,
  input         _EVAL_38,
  output [3:0]  _EVAL_39,
  input         _EVAL_40,
  input         _EVAL_41,
  input         _EVAL_42,
  input  [3:0]  _EVAL_43,
  input         _EVAL_44,
  output [2:0]  _EVAL_45,
  output        _EVAL_46,
  output        _EVAL_47,
  output [1:0]  _EVAL_48,
  input         _EVAL_49,
  output        _EVAL_50,
  input         _EVAL_51,
  output [3:0]  _EVAL_52,
  input  [31:0] _EVAL_53,
  input  [2:0]  _EVAL_54,
  output        _EVAL_55,
  input  [2:0]  _EVAL_56,
  output        _EVAL_57,
  input         _EVAL_58,
  output        _EVAL_59,
  output        _EVAL_60,
  input  [2:0]  _EVAL_61,
  output        _EVAL_62,
  input         _EVAL_63,
  output        _EVAL_64,
  input         _EVAL_65,
  input  [31:0] _EVAL_66,
  input  [3:0]  _EVAL_67,
  output [2:0]  _EVAL_68,
  input         _EVAL_69,
  output        _EVAL_70,
  output        _EVAL_71,
  output [2:0]  _EVAL_72,
  input  [2:0]  _EVAL_73,
  input         _EVAL_74,
  input  [31:0] _EVAL_75,
  input         _EVAL_76,
  output        _EVAL_77,
  input         _EVAL_78,
  input         _EVAL_79,
  output        _EVAL_80,
  input  [1:0]  _EVAL_81,
  input         _EVAL_82,
  output        _EVAL_83,
  output [31:0] _EVAL_84,
  input         _EVAL_85,
  input  [3:0]  _EVAL_86,
  output [2:0]  _EVAL_87,
  output        _EVAL_88,
  input         _EVAL_89,
  input  [3:0]  _EVAL_90,
  input         _EVAL_91,
  input         _EVAL_92,
  output [2:0]  _EVAL_93,
  output        _EVAL_94,
  output        _EVAL_95,
  input  [31:0] _EVAL_96,
  input         _EVAL_97,
  output [31:0] _EVAL_98,
  output        _EVAL_99,
  input  [3:0]  _EVAL_100,
  output        _EVAL_101,
  output [3:0]  _EVAL_102,
  input         _EVAL_103,
  output        _EVAL_104,
  input         _EVAL_105,
  output [31:0] _EVAL_106,
  output        _EVAL_107,
  input         _EVAL_108
);
  assign _EVAL_101 = _EVAL_91;
  assign _EVAL_106 = _EVAL_66;
  assign _EVAL_8 = _EVAL_63;
  assign _EVAL_59 = _EVAL_42;
  assign _EVAL_104 = _EVAL_38;
  assign _EVAL_11 = _EVAL_51;
  assign _EVAL_26 = _EVAL_13;
  assign _EVAL_20 = _EVAL_10;
  assign _EVAL_107 = _EVAL_2;
  assign _EVAL_45 = _EVAL_61;
  assign _EVAL_46 = _EVAL_44;
  assign _EVAL_72 = _EVAL_54;
  assign _EVAL_87 = _EVAL_73;
  assign _EVAL_50 = _EVAL_92;
  assign _EVAL_24 = _EVAL_100;
  assign _EVAL_57 = _EVAL_58;
  assign _EVAL_15 = _EVAL_78;
  assign _EVAL_99 = _EVAL_25;
  assign _EVAL_4 = _EVAL_97;
  assign _EVAL_102 = _EVAL_67;
  assign _EVAL_68 = _EVAL_0;
  assign _EVAL_3 = _EVAL;
  assign _EVAL_7 = _EVAL_30;
  assign _EVAL_84 = _EVAL_53;
  assign _EVAL_64 = _EVAL_31;
  assign _EVAL_9 = _EVAL_18;
  assign _EVAL_70 = _EVAL_74;
  assign _EVAL_32 = _EVAL_81;
  assign _EVAL_22 = _EVAL_69;
  assign _EVAL_19 = _EVAL_103;
  assign _EVAL_14 = _EVAL_108;
  assign _EVAL_35 = _EVAL_90;
  assign _EVAL_21 = _EVAL_105;
  assign _EVAL_28 = _EVAL_16;
  assign _EVAL_95 = _EVAL_82;
  assign _EVAL_98 = _EVAL_96;
  assign _EVAL_62 = _EVAL_5;
  assign _EVAL_77 = _EVAL_89;
  assign _EVAL_48 = _EVAL_17;
  assign _EVAL_47 = _EVAL_49;
  assign _EVAL_88 = _EVAL_65;
  assign _EVAL_27 = _EVAL_37;
  assign _EVAL_80 = _EVAL_29;
  assign _EVAL_39 = _EVAL_86;
  assign _EVAL_6 = _EVAL_75;
  assign _EVAL_60 = _EVAL_76;
  assign _EVAL_36 = _EVAL_1;
  assign _EVAL_93 = _EVAL_56;
  assign _EVAL_23 = _EVAL_79;
  assign _EVAL_83 = _EVAL_34;
  assign _EVAL_55 = _EVAL_41;
  assign _EVAL_52 = _EVAL_43;
  assign _EVAL_71 = _EVAL_85;
  assign _EVAL_94 = _EVAL_12;
endmodule
