//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_164(
  input  [2:0]  _EVAL,
  input  [3:0]  _EVAL_0,
  input         _EVAL_1,
  output        _EVAL_2,
  output        _EVAL_3,
  output [3:0]  _EVAL_4,
  output [3:0]  _EVAL_5,
  input  [31:0] _EVAL_6,
  output [31:0] _EVAL_7,
  output        _EVAL_8,
  output [31:0] _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  output        _EVAL_12,
  output        _EVAL_13,
  input         _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16,
  output        _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19,
  input         _EVAL_20,
  input         _EVAL_21,
  output        _EVAL_22,
  output        _EVAL_23,
  input         _EVAL_24,
  input  [3:0]  _EVAL_25,
  input  [3:0]  _EVAL_26,
  input  [31:0] _EVAL_27,
  input         _EVAL_28,
  output        _EVAL_29,
  output [2:0]  _EVAL_30,
  input         _EVAL_31,
  output        _EVAL_32,
  output        _EVAL_33,
  input         _EVAL_34,
  input  [31:0] _EVAL_35,
  output [31:0] _EVAL_36,
  output [31:0] _EVAL_37,
  input         _EVAL_38,
  input  [1:0]  _EVAL_39,
  input         _EVAL_40,
  input         _EVAL_41,
  output        _EVAL_42,
  input  [31:0] _EVAL_43,
  input         _EVAL_44,
  input         _EVAL_45,
  output [2:0]  _EVAL_46,
  output [3:0]  _EVAL_47,
  input  [2:0]  _EVAL_48,
  output        _EVAL_49,
  output        _EVAL_50,
  output        _EVAL_51,
  input         _EVAL_52,
  input         _EVAL_53,
  output [1:0]  _EVAL_54,
  output        _EVAL_55,
  output [2:0]  _EVAL_56,
  output [31:0] _EVAL_57,
  input         _EVAL_58,
  input         _EVAL_59,
  output        _EVAL_60,
  input  [3:0]  _EVAL_61,
  input         _EVAL_62,
  output [31:0] _EVAL_63,
  output [3:0]  _EVAL_64,
  input         _EVAL_65,
  input         _EVAL_66,
  input         _EVAL_67,
  output        _EVAL_68,
  output        _EVAL_69,
  output        _EVAL_70,
  input         _EVAL_71,
  input  [2:0]  _EVAL_72,
  output [2:0]  _EVAL_73,
  input         _EVAL_74,
  input         _EVAL_75,
  output        _EVAL_76,
  output [3:0]  _EVAL_77,
  output        _EVAL_78,
  output        _EVAL_79,
  output        _EVAL_80,
  output        _EVAL_81,
  input  [1:0]  _EVAL_82,
  output        _EVAL_83,
  input  [3:0]  _EVAL_84,
  input         _EVAL_85,
  output        _EVAL_86,
  output [2:0]  _EVAL_87,
  output        _EVAL_88,
  output        _EVAL_89,
  input         _EVAL_90,
  input         _EVAL_91,
  input  [31:0] _EVAL_92,
  output [3:0]  _EVAL_93,
  input  [2:0]  _EVAL_94,
  output [1:0]  _EVAL_95,
  input         _EVAL_96,
  output        _EVAL_97,
  input         _EVAL_98,
  output        _EVAL_99,
  input  [3:0]  _EVAL_100,
  output [2:0]  _EVAL_101,
  input  [31:0] _EVAL_102,
  input         _EVAL_103,
  input         _EVAL_104,
  input         _EVAL_105,
  input         _EVAL_106,
  output        _EVAL_107,
  output        _EVAL_108
);
  assign _EVAL_8 = _EVAL_24;
  assign _EVAL_86 = _EVAL_28;
  assign _EVAL_108 = _EVAL_65;
  assign _EVAL_50 = _EVAL_11;
  assign _EVAL_55 = _EVAL_66;
  assign _EVAL_64 = _EVAL_84;
  assign _EVAL_12 = _EVAL_71;
  assign _EVAL_63 = _EVAL_6;
  assign _EVAL_30 = _EVAL_10;
  assign _EVAL_46 = _EVAL;
  assign _EVAL_77 = _EVAL_61;
  assign _EVAL_23 = _EVAL_58;
  assign _EVAL_7 = _EVAL_35;
  assign _EVAL_17 = _EVAL_62;
  assign _EVAL_81 = _EVAL_103;
  assign _EVAL_57 = _EVAL_102;
  assign _EVAL_29 = _EVAL_104;
  assign _EVAL_4 = _EVAL_0;
  assign _EVAL_37 = _EVAL_43;
  assign _EVAL_83 = _EVAL_74;
  assign _EVAL_22 = _EVAL_41;
  assign _EVAL_80 = _EVAL_98;
  assign _EVAL_93 = _EVAL_100;
  assign _EVAL_60 = _EVAL_45;
  assign _EVAL_68 = _EVAL_75;
  assign _EVAL_88 = _EVAL_31;
  assign _EVAL_33 = _EVAL_38;
  assign _EVAL_9 = _EVAL_92;
  assign _EVAL_3 = _EVAL_59;
  assign _EVAL_42 = _EVAL_91;
  assign _EVAL_69 = _EVAL_67;
  assign _EVAL_70 = _EVAL_14;
  assign _EVAL_54 = _EVAL_39;
  assign _EVAL_36 = _EVAL_27;
  assign _EVAL_101 = _EVAL_94;
  assign _EVAL_76 = _EVAL_44;
  assign _EVAL_107 = _EVAL_1;
  assign _EVAL_49 = _EVAL_96;
  assign _EVAL_32 = _EVAL_20;
  assign _EVAL_97 = _EVAL_53;
  assign _EVAL_78 = _EVAL_34;
  assign _EVAL_5 = _EVAL_25;
  assign _EVAL_2 = _EVAL_21;
  assign _EVAL_99 = _EVAL_106;
  assign _EVAL_47 = _EVAL_26;
  assign _EVAL_95 = _EVAL_82;
  assign _EVAL_13 = _EVAL_19;
  assign _EVAL_18 = _EVAL_16;
  assign _EVAL_56 = _EVAL_15;
  assign _EVAL_87 = _EVAL_48;
  assign _EVAL_73 = _EVAL_72;
  assign _EVAL_79 = _EVAL_52;
  assign _EVAL_89 = _EVAL_40;
  assign _EVAL_51 = _EVAL_90;
endmodule
