//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_35(
  input  [1:0]  _EVAL,
  output        _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  output [3:0]  _EVAL_3,
  input         _EVAL_4,
  output        _EVAL_5,
  output        _EVAL_6,
  input  [31:0] _EVAL_7,
  input         _EVAL_8,
  output        _EVAL_9,
  output        _EVAL_10,
  input         _EVAL_11,
  output        _EVAL_12,
  input  [2:0]  _EVAL_13,
  output [31:0] _EVAL_14,
  input         _EVAL_15,
  output        _EVAL_16,
  input         _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19,
  input  [31:0] _EVAL_20,
  output        _EVAL_21,
  input         _EVAL_22,
  output [3:0]  _EVAL_23,
  input         _EVAL_24,
  output        _EVAL_25,
  output [2:0]  _EVAL_26,
  output [31:0] _EVAL_27,
  input  [3:0]  _EVAL_28,
  output        _EVAL_29,
  output [1:0]  _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  output        _EVAL_33,
  input         _EVAL_34,
  output [2:0]  _EVAL_35,
  input  [3:0]  _EVAL_36,
  input         _EVAL_37,
  input  [3:0]  _EVAL_38,
  input  [31:0] _EVAL_39,
  input         _EVAL_40,
  input         _EVAL_41,
  input  [2:0]  _EVAL_42,
  output        _EVAL_43,
  output [2:0]  _EVAL_44,
  output        _EVAL_45,
  output        _EVAL_46,
  output        _EVAL_47,
  input         _EVAL_48,
  output [3:0]  _EVAL_49,
  input         _EVAL_50,
  input         _EVAL_51,
  output [31:0] _EVAL_52
);
  assign _EVAL_0 = _EVAL_34;
  assign _EVAL_5 = _EVAL_50;
  assign _EVAL_30 = _EVAL;
  assign _EVAL_10 = _EVAL_37;
  assign _EVAL_52 = _EVAL_20;
  assign _EVAL_18 = _EVAL_48;
  assign _EVAL_45 = _EVAL_41;
  assign _EVAL_14 = _EVAL_7;
  assign _EVAL_6 = _EVAL_4;
  assign _EVAL_21 = _EVAL_24;
  assign _EVAL_49 = _EVAL_28;
  assign _EVAL_23 = _EVAL_38;
  assign _EVAL_12 = _EVAL_17;
  assign _EVAL_29 = _EVAL_51;
  assign _EVAL_46 = _EVAL_11;
  assign _EVAL_35 = _EVAL_1;
  assign _EVAL_33 = _EVAL_8;
  assign _EVAL_47 = _EVAL_40;
  assign _EVAL_44 = _EVAL_42;
  assign _EVAL_16 = _EVAL_22;
  assign _EVAL_26 = _EVAL_13;
  assign _EVAL_43 = _EVAL_15;
  assign _EVAL_27 = _EVAL_39;
  assign _EVAL_25 = _EVAL_31;
  assign _EVAL_9 = _EVAL_2;
  assign _EVAL_3 = _EVAL_36;
endmodule
