//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_27_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input  [3:0]  _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input  [1:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [30:0] _EVAL_13,
  input         _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16,
  input  [2:0]  _EVAL_17,
  input         _EVAL_18
);
  wire [4:0] _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire [5:0] _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire [31:0] _EVAL_30;
  wire [4:0] _EVAL_31;
  reg [2:0] _EVAL_32;
  reg [31:0] _RAND_0;
  wire  _EVAL_33;
  reg [1:0] _EVAL_34;
  reg [31:0] _RAND_1;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire [3:0] _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire [3:0] _EVAL_49;
  wire  _EVAL_50;
  reg [3:0] _EVAL_51;
  reg [31:0] _RAND_2;
  wire  _EVAL_52;
  wire [31:0] _EVAL_53;
  wire [7:0] _EVAL_54;
  wire  _EVAL_55;
  wire [1:0] _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire [32:0] _EVAL_61;
  reg  _EVAL_62;
  reg [31:0] _RAND_3;
  wire [12:0] _EVAL_63;
  wire [4:0] _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  reg  _EVAL_67;
  reg [31:0] _RAND_4;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire [3:0] _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire [4:0] _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire [3:0] _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire [30:0] _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_95;
  wire [5:0] _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire [1:0] _EVAL_101;
  wire  _EVAL_102;
  reg [2:0] _EVAL_103;
  reg [31:0] _RAND_5;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire [7:0] _EVAL_108;
  reg [30:0] _EVAL_109;
  reg [31:0] _RAND_6;
  wire  _EVAL_110;
  wire [4:0] _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire [4:0] _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  reg [2:0] _EVAL_121;
  reg [31:0] _RAND_7;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire [3:0] _EVAL_124;
  wire [5:0] _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire [31:0] _EVAL_130;
  wire [12:0] _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  reg [2:0] _EVAL_137;
  reg [31:0] _RAND_8;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [7:0] _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  reg [2:0] _EVAL_149;
  reg [31:0] _RAND_9;
  wire  _EVAL_150;
  wire [3:0] _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire [30:0] _EVAL_154;
  wire  _EVAL_155;
  wire [4:0] _EVAL_156;
  reg [4:0] _EVAL_157;
  reg [31:0] _RAND_10;
  wire [7:0] _EVAL_158;
  wire [3:0] _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire [4:0] _EVAL_169;
  wire  _EVAL_170;
  wire [30:0] _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire [5:0] _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire [4:0] _EVAL_192;
  wire  _EVAL_194;
  reg [2:0] _EVAL_195;
  reg [31:0] _RAND_11;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire [31:0] _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire [3:0] _EVAL_207;
  reg [31:0] _EVAL_208;
  reg [31:0] _RAND_12;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire [1:0] _EVAL_218;
  wire [1:0] _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire [4:0] _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_236;
  wire [4:0] _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  reg [3:0] _EVAL_245;
  reg [31:0] _RAND_13;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_250;
  reg [2:0] _EVAL_251;
  reg [31:0] _RAND_14;
  wire  _EVAL_252;
  wire [4:0] _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  reg [3:0] _EVAL_267;
  reg [31:0] _RAND_15;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire [3:0] _EVAL_287;
  wire [3:0] _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  reg [3:0] _EVAL_293;
  reg [31:0] _RAND_16;
  wire  _EVAL_294;
  wire  _EVAL_295;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_105 = _EVAL_0 == 3'h1;
  assign _EVAL_269 = ~_EVAL_176;
  assign _EVAL_36 = _EVAL_56 == 2'h1;
  assign _EVAL_86 = _EVAL_203 | _EVAL_11;
  assign _EVAL_96 = _EVAL_131[5:0];
  assign _EVAL_54 = 8'h1 << _EVAL_10;
  assign _EVAL_63 = 13'h3f << _EVAL_9;
  assign _EVAL_218 = _EVAL_219 | 2'h1;
  assign _EVAL_187 = _EVAL_98 & _EVAL_75;
  assign _EVAL_76 = _EVAL_148 | _EVAL_11;
  assign _EVAL_28 = _EVAL_140 | _EVAL_11;
  assign _EVAL_23 = _EVAL_201 & _EVAL_126;
  assign _EVAL_176 = _EVAL_172 | _EVAL_11;
  assign _EVAL_37 = _EVAL_13 == _EVAL_109;
  assign _EVAL_213 = _EVAL_263 | _EVAL_11;
  assign _EVAL_61 = _EVAL_208 + 32'h1;
  assign _EVAL_98 = _EVAL_218[0];
  assign _EVAL_74 = _EVAL_0[0];
  assign _EVAL_85 = _EVAL_194 | _EVAL_16;
  assign _EVAL_87 = _EVAL_17 == 3'h7;
  assign _EVAL_153 = _EVAL_29 | _EVAL_11;
  assign _EVAL_152 = _EVAL_201 & _EVAL_27;
  assign _EVAL_128 = _EVAL_72 & _EVAL_38;
  assign _EVAL_275 = _EVAL_17[2];
  assign _EVAL_225 = _EVAL_118 | _EVAL_11;
  assign _EVAL_203 = _EVAL_4 == _EVAL_32;
  assign _EVAL_21 = _EVAL_5 & _EVAL_268;
  assign _EVAL_189 = ~_EVAL_285;
  assign _EVAL_219 = 2'h1 << _EVAL_290;
  assign _EVAL_119 = _EVAL_55 & _EVAL_173;
  assign _EVAL_53 = {1'b0,$signed(_EVAL_171)};
  assign _EVAL_46 = _EVAL_253 != _EVAL_229;
  assign _EVAL_148 = _EVAL_4 <= 3'h3;
  assign _EVAL_201 = _EVAL_18 & _EVAL_1;
  assign _EVAL_252 = _EVAL_13[1];
  assign _EVAL_106 = ~_EVAL_146;
  assign _EVAL_262 = ~_EVAL_277;
  assign _EVAL_171 = _EVAL_13 ^ 31'h40000000;
  assign _EVAL_29 = _EVAL_6 == _EVAL_103;
  assign _EVAL_35 = _EVAL_97 | _EVAL_11;
  assign _EVAL_174 = ~_EVAL_27;
  assign _EVAL_194 = ~_EVAL_7;
  assign _EVAL_209 = ~_EVAL_231;
  assign _EVAL_124 = _EVAL_156[3:0];
  assign _EVAL_100 = ~_EVAL_196;
  assign _EVAL_281 = _EVAL_52 | _EVAL_11;
  assign _EVAL_57 = _EVAL_147 | _EVAL_184;
  assign _EVAL_116 = _EVAL_293 - 4'h1;
  assign _EVAL_265 = _EVAL_253 != 5'h0;
  assign _EVAL_31 = _EVAL_19 & _EVAL_237;
  assign _EVAL_81 = _EVAL_5 & _EVAL_295;
  assign _EVAL_192 = _EVAL_157 >> _EVAL_10;
  assign _EVAL_228 = ~_EVAL_265;
  assign _EVAL_141 = _EVAL_284 | _EVAL_11;
  assign _EVAL_284 = _EVAL_8 == 2'h0;
  assign _EVAL_294 = _EVAL_17 == _EVAL_149;
  assign _EVAL_144 = _EVAL_10 == _EVAL_251;
  assign _EVAL_283 = _EVAL_170 | _EVAL_11;
  assign _EVAL_156 = _EVAL_267 - 4'h1;
  assign _EVAL_160 = _EVAL_17 == 3'h5;
  assign _EVAL_40 = _EVAL_119 | _EVAL_11;
  assign _EVAL_38 = _EVAL_267 == 4'h0;
  assign _EVAL_111 = _EVAL_169 >> _EVAL_6;
  assign _EVAL_285 = _EVAL_192[0];
  assign _EVAL_68 = _EVAL_198 | _EVAL_11;
  assign _EVAL_264 = _EVAL_236 | _EVAL_11;
  assign _EVAL_184 = _EVAL_98 & _EVAL_79;
  assign _EVAL_282 = _EVAL_24 | _EVAL_255;
  assign _EVAL_291 = _EVAL_201 | _EVAL_72;
  assign _EVAL_224 = ~_EVAL_206;
  assign _EVAL_185 = ~_EVAL_153;
  assign _EVAL_78 = _EVAL_51 - 4'h1;
  assign _EVAL_134 = ~_EVAL_210;
  assign _EVAL_48 = _EVAL_0 == 3'h0;
  assign _EVAL_173 = $signed(_EVAL_130) == 32'sh0;
  assign _EVAL_142 = ~_EVAL_141;
  assign _EVAL_227 = _EVAL_39 == 4'h0;
  assign _EVAL_49 = ~_EVAL_3;
  assign _EVAL_289 = _EVAL_102 | _EVAL_11;
  assign _EVAL_199 = _EVAL_61[31:0];
  assign _EVAL_220 = ~_EVAL_271;
  assign _EVAL_210 = _EVAL_37 | _EVAL_11;
  assign _EVAL_47 = _EVAL_4 <= 3'h2;
  assign _EVAL_135 = _EVAL_98 & _EVAL_292;
  assign _EVAL_45 = _EVAL_8 != 2'h2;
  assign _EVAL_64 = _EVAL_245 - 4'h1;
  assign _EVAL_260 = _EVAL_157 != 5'h0;
  assign _EVAL_151 = ~_EVAL_70;
  assign _EVAL_177 = ~_EVAL_200;
  assign _EVAL_178 = _EVAL_5 & _EVAL_240;
  assign _EVAL_39 = _EVAL_3 & _EVAL_151;
  assign _EVAL_212 = _EVAL_8 == _EVAL_34;
  assign _EVAL_138 = ~_EVAL_182;
  assign _EVAL_287 = _EVAL_116[3:0];
  assign _EVAL_136 = _EVAL_5 & _EVAL_105;
  assign _EVAL_232 = _EVAL_111[0];
  assign _EVAL_19 = _EVAL_157 | _EVAL_253;
  assign _EVAL_169 = _EVAL_253 | _EVAL_157;
  assign _EVAL_41 = _EVAL_194 | _EVAL_11;
  assign _EVAL_167 = ~_EVAL_264;
  assign _EVAL_290 = _EVAL_9[0];
  assign _EVAL_211 = ~_EVAL_295;
  assign _EVAL_58 = _EVAL_17 == 3'h0;
  assign _EVAL_107 = _EVAL_45 | _EVAL_11;
  assign _EVAL_114 = ~_EVAL_270;
  assign _EVAL_243 = _EVAL_9 >= 3'h2;
  assign _EVAL_259 = _EVAL_5 & _EVAL_215;
  assign _EVAL_271 = _EVAL_47 | _EVAL_11;
  assign _EVAL_233 = _EVAL_17 == 3'h4;
  assign _EVAL_129 = _EVAL_133 | _EVAL_187;
  assign _EVAL_254 = _EVAL_43 & _EVAL_252;
  assign _EVAL_263 = _EVAL_3 == _EVAL_70;
  assign _EVAL_240 = _EVAL_0 == 3'h2;
  assign _EVAL_188 = ~_EVAL_69;
  assign _EVAL_255 = _EVAL_10 == 3'h4;
  assign _EVAL_75 = _EVAL_252 & _EVAL_277;
  assign _EVAL_143 = _EVAL_23 ? _EVAL_54 : 8'h0;
  assign _EVAL_159 = _EVAL_78[3:0];
  assign _EVAL_92 = _EVAL_13 & _EVAL_154;
  assign _EVAL_113 = ~_EVAL_16;
  assign _EVAL_33 = ~_EVAL_155;
  assign _EVAL_93 = _EVAL_145 & _EVAL_211;
  assign _EVAL_97 = _EVAL_15 >= 3'h2;
  assign _EVAL_24 = _EVAL_36 | _EVAL_127;
  assign _EVAL_27 = _EVAL_293 == 4'h0;
  assign _EVAL_237 = ~_EVAL_229;
  assign _EVAL_277 = _EVAL_13[0];
  assign _EVAL_89 = _EVAL_64[3:0];
  assign _EVAL_288 = _EVAL_125[5:2];
  assign _EVAL_268 = ~_EVAL_38;
  assign _EVAL_145 = _EVAL_72 & _EVAL_22;
  assign _EVAL_241 = _EVAL_208 < plusarg_reader_out;
  assign _EVAL_236 = _EVAL_0 == _EVAL_195;
  assign _EVAL_166 = _EVAL_101 == 2'h1;
  assign _EVAL_276 = _EVAL_101 == 2'h0;
  assign _EVAL_170 = _EVAL_279 | _EVAL_241;
  assign _EVAL_207 = _EVAL_186[5:2];
  assign _EVAL_26 = _EVAL_63[5:0];
  assign _EVAL_215 = _EVAL_0 == 3'h4;
  assign _EVAL_158 = 8'h1 << _EVAL_6;
  assign _EVAL_112 = ~_EVAL_76;
  assign _EVAL_126 = _EVAL_245 == 4'h0;
  assign _EVAL_80 = _EVAL_17 == 3'h3;
  assign _EVAL_216 = _EVAL_1 & _EVAL_87;
  assign _EVAL_72 = _EVAL_14 & _EVAL_5;
  assign _EVAL_154 = {{25'd0}, _EVAL_186};
  assign _EVAL_190 = _EVAL_133 | _EVAL_246;
  assign _EVAL_146 = _EVAL_189 | _EVAL_11;
  assign _EVAL_205 = ~_EVAL_132;
  assign _EVAL_183 = ~_EVAL_281;
  assign _EVAL_246 = _EVAL_98 & _EVAL_123;
  assign _EVAL_186 = ~_EVAL_26;
  assign _EVAL_278 = ~_EVAL_86;
  assign _EVAL_102 = ~_EVAL_2;
  assign _EVAL_110 = ~_EVAL_20;
  assign _EVAL_198 = _EVAL_7 == _EVAL_62;
  assign _EVAL_161 = ~_EVAL_40;
  assign _EVAL_65 = _EVAL_166 | _EVAL_276;
  assign _EVAL_175 = _EVAL_5 & _EVAL_84;
  assign _EVAL_147 = _EVAL_243 | _EVAL_73;
  assign _EVAL_66 = _EVAL_6 == 3'h4;
  assign _EVAL_56 = _EVAL_10[2:1];
  assign _EVAL_82 = _EVAL_46 | _EVAL_228;
  assign _EVAL_130 = _EVAL_30;
  assign _EVAL_292 = _EVAL_242 & _EVAL_262;
  assign _EVAL_261 = _EVAL_0 <= 3'h6;
  assign _EVAL_117 = ~_EVAL_164;
  assign _EVAL_242 = ~_EVAL_252;
  assign _EVAL_95 = ~_EVAL_99;
  assign _EVAL_204 = _EVAL_1 & _EVAL_80;
  assign _EVAL_139 = ~_EVAL_275;
  assign _EVAL_206 = _EVAL_232 | _EVAL_11;
  assign _EVAL_60 = _EVAL_4 != 3'h0;
  assign _EVAL_239 = _EVAL_4 == 3'h0;
  assign _EVAL_238 = _EVAL_4 <= 3'h4;
  assign _EVAL_270 = _EVAL_85 | _EVAL_11;
  assign _EVAL_182 = _EVAL_282 | _EVAL_11;
  assign _EVAL_168 = _EVAL_17 == 3'h2;
  assign _EVAL_191 = _EVAL_49 == 4'h0;
  assign _EVAL_253 = _EVAL_143[4:0];
  assign _EVAL_77 = ~_EVAL_260;
  assign _EVAL_279 = _EVAL_77 | _EVAL_25;
  assign _EVAL_123 = _EVAL_252 & _EVAL_262;
  assign _EVAL_280 = _EVAL_5 & _EVAL_48;
  assign _EVAL_122 = ~_EVAL_197;
  assign _EVAL_250 = _EVAL_71 | _EVAL_11;
  assign _EVAL_88 = _EVAL_144 | _EVAL_11;
  assign _EVAL_202 = ~_EVAL_289;
  assign _EVAL_221 = _EVAL_1 & _EVAL_233;
  assign _EVAL_230 = _EVAL_147 | _EVAL_135;
  assign _EVAL_42 = ~_EVAL_283;
  assign _EVAL_44 = ~_EVAL_104;
  assign _EVAL_131 = 13'h3f << _EVAL_15;
  assign _EVAL_155 = _EVAL_191 | _EVAL_11;
  assign _EVAL_59 = _EVAL_294 | _EVAL_11;
  assign _EVAL_197 = _EVAL_115 | _EVAL_11;
  assign _EVAL_273 = _EVAL_65 | _EVAL_66;
  assign _EVAL_226 = ~_EVAL_225;
  assign _EVAL_52 = _EVAL_12 == _EVAL_67;
  assign _EVAL_71 = _EVAL_9 == _EVAL_121;
  assign _EVAL_274 = ~_EVAL_50;
  assign _EVAL_181 = ~_EVAL_250;
  assign _EVAL_118 = _EVAL_4 <= 3'h1;
  assign _EVAL_73 = _EVAL_43 & _EVAL_242;
  assign _EVAL_196 = _EVAL_212 | _EVAL_11;
  assign _EVAL_172 = _EVAL_15 == _EVAL_137;
  assign _EVAL_257 = _EVAL_1 & _EVAL_174;
  assign _EVAL_234 = _EVAL_1 & _EVAL_160;
  assign _EVAL_84 = _EVAL_0 == 3'h5;
  assign _EVAL_108 = _EVAL_93 ? _EVAL_158 : 8'h0;
  assign _EVAL_115 = _EVAL_92 == 31'h0;
  assign _EVAL_20 = _EVAL_82 | _EVAL_11;
  assign _EVAL_256 = _EVAL_1 & _EVAL_168;
  assign _EVAL_79 = _EVAL_242 & _EVAL_277;
  assign _EVAL_180 = ~_EVAL_213;
  assign _EVAL_55 = _EVAL_9 <= 3'h6;
  assign _EVAL_83 = ~_EVAL_35;
  assign _EVAL_132 = _EVAL_60 | _EVAL_11;
  assign _EVAL_179 = ~_EVAL_11;
  assign _EVAL_164 = _EVAL_243 | _EVAL_11;
  assign _EVAL_231 = _EVAL_273 | _EVAL_11;
  assign _EVAL_140 = _EVAL_8 <= 2'h2;
  assign _EVAL_248 = ~_EVAL_41;
  assign _EVAL_295 = _EVAL_0 == 3'h6;
  assign _EVAL_150 = _EVAL_17 == 3'h6;
  assign _EVAL_99 = _EVAL_261 | _EVAL_11;
  assign _EVAL_165 = _EVAL_1 & _EVAL_58;
  assign _EVAL_30 = $signed(_EVAL_53) & -32'sh2000;
  assign _EVAL_50 = _EVAL_239 | _EVAL_11;
  assign _EVAL_120 = _EVAL_17 == 3'h1;
  assign _EVAL_25 = plusarg_reader_out == 32'h0;
  assign _EVAL_69 = _EVAL_238 | _EVAL_11;
  assign _EVAL_286 = ~_EVAL_88;
  assign _EVAL_222 = _EVAL_1 & _EVAL_120;
  assign _EVAL_244 = _EVAL_1 & _EVAL_150;
  assign _EVAL_70 = {_EVAL_129,_EVAL_190,_EVAL_57,_EVAL_230};
  assign _EVAL_200 = _EVAL_113 | _EVAL_11;
  assign _EVAL_272 = ~_EVAL_107;
  assign _EVAL_101 = _EVAL_6[2:1];
  assign _EVAL_247 = ~_EVAL_28;
  assign _EVAL_127 = _EVAL_56 == 2'h0;
  assign _EVAL_133 = _EVAL_243 | _EVAL_254;
  assign _EVAL_125 = ~_EVAL_96;
  assign _EVAL_104 = _EVAL_227 | _EVAL_11;
  assign _EVAL_22 = _EVAL_51 == 4'h0;
  assign _EVAL_229 = _EVAL_108[4:0];
  assign _EVAL_90 = ~_EVAL_59;
  assign _EVAL_91 = ~_EVAL_68;
  assign _EVAL_43 = _EVAL_218[1];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_32 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_34 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_51 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_62 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_67 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_103 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_109 = _RAND_6[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_121 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_137 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_149 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_157 = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_195 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_208 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_245 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_251 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_267 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_293 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL) begin
    if (_EVAL_152) begin
      _EVAL_32 <= _EVAL_4;
    end
    if (_EVAL_128) begin
      _EVAL_34 <= _EVAL_8;
    end
    if (_EVAL_11) begin
      _EVAL_51 <= 4'h0;
    end else if (_EVAL_72) begin
      if (_EVAL_22) begin
        if (_EVAL_74) begin
          _EVAL_51 <= _EVAL_288;
        end else begin
          _EVAL_51 <= 4'h0;
        end
      end else begin
        _EVAL_51 <= _EVAL_159;
      end
    end
    if (_EVAL_128) begin
      _EVAL_62 <= _EVAL_7;
    end
    if (_EVAL_128) begin
      _EVAL_67 <= _EVAL_12;
    end
    if (_EVAL_128) begin
      _EVAL_103 <= _EVAL_6;
    end
    if (_EVAL_152) begin
      _EVAL_109 <= _EVAL_13;
    end
    if (_EVAL_152) begin
      _EVAL_121 <= _EVAL_9;
    end
    if (_EVAL_128) begin
      _EVAL_137 <= _EVAL_15;
    end
    if (_EVAL_152) begin
      _EVAL_149 <= _EVAL_17;
    end
    if (_EVAL_11) begin
      _EVAL_157 <= 5'h0;
    end else begin
      _EVAL_157 <= _EVAL_31;
    end
    if (_EVAL_128) begin
      _EVAL_195 <= _EVAL_0;
    end
    if (_EVAL_11) begin
      _EVAL_208 <= 32'h0;
    end else if (_EVAL_291) begin
      _EVAL_208 <= 32'h0;
    end else begin
      _EVAL_208 <= _EVAL_199;
    end
    if (_EVAL_11) begin
      _EVAL_245 <= 4'h0;
    end else if (_EVAL_201) begin
      if (_EVAL_126) begin
        if (_EVAL_139) begin
          _EVAL_245 <= _EVAL_207;
        end else begin
          _EVAL_245 <= 4'h0;
        end
      end else begin
        _EVAL_245 <= _EVAL_89;
      end
    end
    if (_EVAL_152) begin
      _EVAL_251 <= _EVAL_10;
    end
    if (_EVAL_11) begin
      _EVAL_267 <= 4'h0;
    end else if (_EVAL_72) begin
      if (_EVAL_38) begin
        if (_EVAL_74) begin
          _EVAL_267 <= _EVAL_288;
        end else begin
          _EVAL_267 <= 4'h0;
        end
      end else begin
        _EVAL_267 <= _EVAL_124;
      end
    end
    if (_EVAL_11) begin
      _EVAL_293 <= 4'h0;
    end else if (_EVAL_201) begin
      if (_EVAL_27) begin
        if (_EVAL_139) begin
          _EVAL_293 <= _EVAL_207;
        end else begin
          _EVAL_293 <= 4'h0;
        end
      end else begin
        _EVAL_293 <= _EVAL_287;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(590bb7d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfd182b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c381a7ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7dc98393)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(150a644a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b678d6cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9f85e8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1f9d6d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5aae083d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3da1149)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a219997d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a5edf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ec0dfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_274) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(496c40de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(838057cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2403d296)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bfb7ba4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4d2bb3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5244e582)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acc598bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d614e5d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(728d8a14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ae2289c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af548851)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45e0894)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abba8d6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9407c91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18934298)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6f5b029)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68a92bf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4367091a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49152e2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64d4e109)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39b5627b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dad53424)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e392ce7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5946042)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d86af58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1356846a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_274) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9699482e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5438e4c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68c4cb41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4636123)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5dd58177)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ed2fe4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b779dd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11c42c7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dec3c92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(718f49b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9ff4cc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89ebfc64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f84e455d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bb9c118)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(496acfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5f76373)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85dd8d47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(659c7995)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bec8c2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38025dae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed3a95ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_274) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(843195cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f1e19cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1d26a0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c92c8c4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e90a2d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(affd3034)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10f8eb3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50ae2cbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(888f78f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(258b1158)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6603b2fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3490b4cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5da18dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a1c53ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a2f2223)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19821de5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69acf6a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(affc04c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe37cd3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d7381ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15185c62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b587bf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5efab74c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d99851b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1d5f1a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(914787fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fafae22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b9b066e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7383f7fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89967b03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_256 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bffcb25d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56696367)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da660764)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
