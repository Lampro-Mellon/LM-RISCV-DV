//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_37(
  output        _EVAL,
  input         _EVAL_0,
  output [30:0] _EVAL_1,
  output [31:0] _EVAL_2,
  output [3:0]  _EVAL_3,
  input  [3:0]  _EVAL_4,
  output [1:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  output        _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [1:0]  _EVAL_10,
  input  [3:0]  _EVAL_11,
  output [2:0]  _EVAL_12,
  output [1:0]  _EVAL_13,
  output        _EVAL_14,
  output [31:0] _EVAL_15,
  output        _EVAL_16,
  output        _EVAL_17,
  output        _EVAL_18,
  output        _EVAL_19,
  output        _EVAL_20,
  output [2:0]  _EVAL_21,
  output        _EVAL_23,
  output        _EVAL_24,
  input  [2:0]  _EVAL_25,
  output [1:0]  _EVAL_26,
  output [3:0]  _EVAL_27,
  output        _EVAL_28,
  output        _EVAL_29,
  output [31:0] _EVAL_30,
  input         _EVAL_31,
  input  [3:0]  _EVAL_32,
  input  [2:0]  _EVAL_33,
  output        _EVAL_34,
  input         _EVAL_36,
  output        _EVAL_37,
  input  [2:0]  _EVAL_38,
  input         _EVAL_39,
  input  [1:0]  _EVAL_41,
  input  [31:0] _EVAL_42,
  input         _EVAL_43,
  input  [2:0]  _EVAL_44,
  input         _EVAL_45,
  input         _EVAL_46,
  output [2:0]  _EVAL_47,
  input         _EVAL_48,
  output        _EVAL_50,
  input         _EVAL_51,
  output [2:0]  _EVAL_52,
  input         _EVAL_53,
  output        _EVAL_54,
  input         _EVAL_55,
  input  [31:0] _EVAL_56,
  output [3:0]  _EVAL_57,
  output [2:0]  _EVAL_58,
  input         _EVAL_59,
  output        _EVAL_60,
  output        _EVAL_61,
  output        _EVAL_62,
  input         _EVAL_63,
  input  [2:0]  _EVAL_64,
  input  [3:0]  _EVAL_65,
  output [2:0]  _EVAL_66,
  output [3:0]  _EVAL_67,
  input         _EVAL_68,
  output        _EVAL_69,
  output [2:0]  _EVAL_70,
  input         _EVAL_71,
  input         _EVAL_72,
  input  [31:0] _EVAL_73,
  input         _EVAL_74,
  output        _EVAL_76,
  input         _EVAL_77,
  input         _EVAL_78,
  output [31:0] _EVAL_79,
  output [3:0]  _EVAL_80,
  output        _EVAL_81,
  input         _EVAL_82,
  output        _EVAL_83,
  input         _EVAL_84,
  input         _EVAL_85,
  output [3:0]  _EVAL_86,
  input  [31:0] _EVAL_87,
  output [1:0]  _EVAL_89,
  output [2:0]  _EVAL_90,
  input         _EVAL_91,
  input         _EVAL_92,
  input         _EVAL_93,
  input  [2:0]  _EVAL_94,
  input         _EVAL_95,
  output        _EVAL_96,
  input         _EVAL_97,
  input  [3:0]  _EVAL_98,
  output [29:0] _EVAL_99,
  output        _EVAL_100,
  input         _EVAL_101,
  input  [3:0]  _EVAL_102,
  input         _EVAL_103,
  input  [31:0] _EVAL_104,
  output        _EVAL_105,
  input  [31:0] _EVAL_106,
  input         _EVAL_107,
  input  [31:0] _EVAL_108,
  input  [1:0]  _EVAL_109,
  input         _EVAL_110,
  input  [31:0] _EVAL_111,
  input  [2:0]  _EVAL_112,
  input         _EVAL_113,
  input         _EVAL_114,
  input  [31:0] _EVAL_115,
  output [2:0]  _EVAL_116,
  input         _EVAL_117,
  output [2:0]  _EVAL_118,
  output [2:0]  _EVAL_119,
  output        _EVAL_120,
  input         _EVAL_121,
  output        _EVAL_122,
  output [2:0]  _EVAL_123,
  output [3:0]  _EVAL_124,
  input  [2:0]  _EVAL_125,
  input  [2:0]  _EVAL_126,
  output [1:0]  _EVAL_128,
  input         _EVAL_129,
  output        _EVAL_130,
  output        _EVAL_131,
  output [3:0]  _EVAL_132,
  input         _EVAL_133,
  input         _EVAL_134,
  output        _EVAL_135,
  output        _EVAL_136,
  input         _EVAL_137,
  output        _EVAL_138,
  input         _EVAL_139,
  output        _EVAL_140,
  input         _EVAL_141,
  output        _EVAL_142,
  input         _EVAL_143,
  output        _EVAL_144,
  input  [2:0]  _EVAL_146,
  output [31:0] _EVAL_147,
  output [31:0] _EVAL_148,
  output [31:0] _EVAL_150,
  input  [3:0]  _EVAL_151,
  input  [2:0]  _EVAL_152,
  input         _EVAL_153,
  output [31:0] _EVAL_154,
  output        _EVAL_156,
  output        _EVAL_157,
  input         _EVAL_158,
  input         _EVAL_159,
  output        _EVAL_160,
  input  [31:0] _EVAL_161,
  output [1:0]  _EVAL_162,
  output [31:0] _EVAL_164,
  output        _EVAL_165,
  output [2:0]  _EVAL_167,
  output [2:0]  _EVAL_168,
  input         _EVAL_169,
  input         _EVAL_170,
  input         _EVAL_171
);
  wire  system_bus_xbar__EVAL;
  wire  system_bus_xbar__EVAL_0;
  wire  system_bus_xbar__EVAL_1;
  wire [2:0] system_bus_xbar__EVAL_2;
  wire [29:0] system_bus_xbar__EVAL_3;
  wire  system_bus_xbar__EVAL_4;
  wire  system_bus_xbar__EVAL_5;
  wire [3:0] system_bus_xbar__EVAL_6;
  wire [3:0] system_bus_xbar__EVAL_7;
  wire [1:0] system_bus_xbar__EVAL_8;
  wire  system_bus_xbar__EVAL_9;
  wire [2:0] system_bus_xbar__EVAL_10;
  wire [3:0] system_bus_xbar__EVAL_11;
  wire  system_bus_xbar__EVAL_12;
  wire  system_bus_xbar__EVAL_13;
  wire  system_bus_xbar__EVAL_14;
  wire [2:0] system_bus_xbar__EVAL_15;
  wire [31:0] system_bus_xbar__EVAL_16;
  wire [1:0] system_bus_xbar__EVAL_17;
  wire  system_bus_xbar__EVAL_18;
  wire [1:0] system_bus_xbar__EVAL_19;
  wire  system_bus_xbar__EVAL_20;
  wire  system_bus_xbar__EVAL_21;
  wire [2:0] system_bus_xbar__EVAL_22;
  wire  system_bus_xbar__EVAL_23;
  wire  system_bus_xbar__EVAL_24;
  wire [2:0] system_bus_xbar__EVAL_25;
  wire  system_bus_xbar__EVAL_26;
  wire [2:0] system_bus_xbar__EVAL_27;
  wire  system_bus_xbar__EVAL_28;
  wire [1:0] system_bus_xbar__EVAL_29;
  wire [2:0] system_bus_xbar__EVAL_30;
  wire  system_bus_xbar__EVAL_31;
  wire  system_bus_xbar__EVAL_32;
  wire  system_bus_xbar__EVAL_33;
  wire [2:0] system_bus_xbar__EVAL_34;
  wire [2:0] system_bus_xbar__EVAL_35;
  wire  system_bus_xbar__EVAL_36;
  wire  system_bus_xbar__EVAL_37;
  wire [1:0] system_bus_xbar__EVAL_38;
  wire [31:0] system_bus_xbar__EVAL_39;
  wire  system_bus_xbar__EVAL_40;
  wire [3:0] system_bus_xbar__EVAL_41;
  wire  system_bus_xbar__EVAL_42;
  wire [2:0] system_bus_xbar__EVAL_43;
  wire  system_bus_xbar__EVAL_44;
  wire  system_bus_xbar__EVAL_45;
  wire  system_bus_xbar__EVAL_46;
  wire  system_bus_xbar__EVAL_47;
  wire  system_bus_xbar__EVAL_48;
  wire  system_bus_xbar__EVAL_49;
  wire [31:0] system_bus_xbar__EVAL_50;
  wire [2:0] system_bus_xbar__EVAL_51;
  wire [3:0] system_bus_xbar__EVAL_52;
  wire [2:0] system_bus_xbar__EVAL_53;
  wire  system_bus_xbar__EVAL_54;
  wire  system_bus_xbar__EVAL_55;
  wire  system_bus_xbar__EVAL_56;
  wire [31:0] system_bus_xbar__EVAL_57;
  wire [31:0] system_bus_xbar__EVAL_58;
  wire [1:0] system_bus_xbar__EVAL_59;
  wire [31:0] system_bus_xbar__EVAL_60;
  wire [3:0] system_bus_xbar__EVAL_61;
  wire  system_bus_xbar__EVAL_62;
  wire  system_bus_xbar__EVAL_63;
  wire  system_bus_xbar__EVAL_64;
  wire [3:0] system_bus_xbar__EVAL_65;
  wire  system_bus_xbar__EVAL_66;
  wire  system_bus_xbar__EVAL_67;
  wire [30:0] system_bus_xbar__EVAL_68;
  wire  system_bus_xbar__EVAL_69;
  wire [2:0] system_bus_xbar__EVAL_70;
  wire  system_bus_xbar__EVAL_71;
  wire [31:0] system_bus_xbar__EVAL_72;
  wire  system_bus_xbar__EVAL_73;
  wire  system_bus_xbar__EVAL_74;
  wire  system_bus_xbar__EVAL_75;
  wire  system_bus_xbar__EVAL_76;
  wire [31:0] system_bus_xbar__EVAL_77;
  wire [2:0] system_bus_xbar__EVAL_78;
  wire [2:0] system_bus_xbar__EVAL_79;
  wire  system_bus_xbar__EVAL_80;
  wire  system_bus_xbar__EVAL_81;
  wire [1:0] system_bus_xbar__EVAL_82;
  wire [31:0] system_bus_xbar__EVAL_83;
  wire  system_bus_xbar__EVAL_84;
  wire [31:0] system_bus_xbar__EVAL_85;
  wire [2:0] system_bus_xbar__EVAL_86;
  wire [2:0] system_bus_xbar__EVAL_87;
  wire  system_bus_xbar__EVAL_88;
  wire [2:0] system_bus_xbar__EVAL_89;
  wire  system_bus_xbar__EVAL_90;
  wire  system_bus_xbar__EVAL_91;
  wire [3:0] system_bus_xbar__EVAL_92;
  wire [2:0] system_bus_xbar__EVAL_93;
  wire  system_bus_xbar__EVAL_94;
  wire [1:0] system_bus_xbar__EVAL_95;
  wire  system_bus_xbar__EVAL_96;
  wire  system_bus_xbar__EVAL_97;
  wire  system_bus_xbar__EVAL_98;
  wire [31:0] system_bus_xbar__EVAL_99;
  wire [31:0] system_bus_xbar__EVAL_100;
  wire [2:0] system_bus_xbar__EVAL_101;
  wire [31:0] system_bus_xbar__EVAL_102;
  wire  system_bus_xbar__EVAL_103;
  wire  system_bus_xbar__EVAL_104;
  wire [3:0] system_bus_xbar__EVAL_105;
  wire [2:0] system_bus_xbar__EVAL_106;
  wire  system_bus_xbar__EVAL_107;
  wire  system_bus_xbar__EVAL_108;
  wire  system_bus_xbar__EVAL_109;
  wire [31:0] system_bus_xbar__EVAL_110;
  wire  system_bus_xbar__EVAL_111;
  wire [2:0] system_bus_xbar__EVAL_112;
  wire  system_bus_xbar__EVAL_113;
  wire [2:0] system_bus_xbar__EVAL_114;
  wire [3:0] system_bus_xbar__EVAL_115;
  wire  system_bus_xbar__EVAL_116;
  wire [31:0] system_bus_xbar__EVAL_117;
  wire [2:0] system_bus_xbar__EVAL_118;
  wire  system_bus_xbar__EVAL_119;
  wire [3:0] system_bus_xbar__EVAL_120;
  wire [2:0] system_bus_xbar__EVAL_121;
  wire  system_bus_xbar__EVAL_122;
  wire [31:0] system_bus_xbar__EVAL_123;
  wire  system_bus_xbar__EVAL_124;
  wire  system_bus_xbar__EVAL_125;
  wire  system_bus_xbar__EVAL_126;
  wire  system_bus_xbar__EVAL_127;
  wire [2:0] system_bus_xbar__EVAL_128;
  wire [2:0] system_bus_xbar__EVAL_129;
  wire [3:0] system_bus_xbar__EVAL_130;
  wire [3:0] system_bus_xbar__EVAL_131;
  wire [31:0] system_bus_xbar__EVAL_132;
  wire  system_bus_xbar__EVAL_133;
  wire [31:0] system_bus_xbar__EVAL_134;
  wire [2:0] system_bus_xbar__EVAL_135;
  wire [31:0] system_bus_xbar__EVAL_136;
  wire [2:0] system_bus_xbar__EVAL_137;
  wire  system_bus_xbar__EVAL_138;
  wire  system_bus_xbar__EVAL_139;
  wire [2:0] system_bus_xbar__EVAL_140;
  wire [3:0] system_bus_xbar__EVAL_141;
  wire [3:0] system_bus_xbar__EVAL_142;
  wire [1:0] system_bus_xbar__EVAL_143;
  wire  system_bus_xbar__EVAL_144;
  wire  system_bus_xbar__EVAL_145;
  wire  system_bus_xbar__EVAL_146;
  wire  system_bus_xbar__EVAL_147;
  wire  system_bus_xbar__EVAL_148;
  wire  system_bus_xbar__EVAL_149;
  wire  system_bus_xbar__EVAL_150;
  wire  system_bus_xbar__EVAL_151;
  wire  system_bus_xbar__EVAL_152;
  wire [2:0] system_bus_xbar__EVAL_153;
  wire  system_bus_xbar__EVAL_154;
  wire  system_bus_xbar__EVAL_155;
  wire  system_bus_xbar__EVAL_156;
  wire  system_bus_xbar__EVAL_157;
  wire  system_bus_xbar__EVAL_158;
  wire  system_bus_xbar__EVAL_159;
  wire  system_bus_xbar__EVAL_160;
  wire  system_bus_xbar__EVAL_161;
  wire  system_bus_xbar__EVAL_162;
  wire  system_bus_xbar__EVAL_163;
  wire  fixedClockNode__EVAL;
  wire  fixedClockNode__EVAL_0;
  wire  fixedClockNode__EVAL_1;
  wire  fixedClockNode__EVAL_2;
  wire  coupler_to_bus_named_cbus__EVAL;
  wire [1:0] coupler_to_bus_named_cbus__EVAL_0;
  wire [3:0] coupler_to_bus_named_cbus__EVAL_1;
  wire  coupler_to_bus_named_cbus__EVAL_2;
  wire [31:0] coupler_to_bus_named_cbus__EVAL_3;
  wire  coupler_to_bus_named_cbus__EVAL_4;
  wire [2:0] coupler_to_bus_named_cbus__EVAL_5;
  wire  coupler_to_bus_named_cbus__EVAL_6;
  wire [31:0] coupler_to_bus_named_cbus__EVAL_7;
  wire [3:0] coupler_to_bus_named_cbus__EVAL_8;
  wire [2:0] coupler_to_bus_named_cbus__EVAL_9;
  wire  coupler_to_bus_named_cbus__EVAL_10;
  wire  coupler_to_bus_named_cbus__EVAL_11;
  wire [3:0] coupler_to_bus_named_cbus__EVAL_12;
  wire  coupler_to_bus_named_cbus__EVAL_13;
  wire [2:0] coupler_to_bus_named_cbus__EVAL_14;
  wire  coupler_to_bus_named_cbus__EVAL_15;
  wire [2:0] coupler_to_bus_named_cbus__EVAL_16;
  wire  coupler_to_bus_named_cbus__EVAL_17;
  wire  coupler_to_bus_named_cbus__EVAL_18;
  wire [2:0] coupler_to_bus_named_cbus__EVAL_19;
  wire  coupler_to_bus_named_cbus__EVAL_20;
  wire [31:0] coupler_to_bus_named_cbus__EVAL_21;
  wire [29:0] coupler_to_bus_named_cbus__EVAL_22;
  wire  coupler_to_bus_named_cbus__EVAL_23;
  wire  coupler_to_bus_named_cbus__EVAL_24;
  wire  coupler_to_bus_named_cbus__EVAL_25;
  wire  coupler_to_bus_named_cbus__EVAL_26;
  wire  coupler_to_bus_named_cbus__EVAL_27;
  wire  coupler_to_bus_named_cbus__EVAL_28;
  wire  coupler_to_bus_named_cbus__EVAL_29;
  wire  coupler_to_bus_named_cbus__EVAL_30;
  wire  coupler_to_bus_named_cbus__EVAL_31;
  wire  coupler_to_bus_named_cbus__EVAL_32;
  wire  coupler_to_bus_named_cbus__EVAL_33;
  wire  coupler_to_bus_named_cbus__EVAL_34;
  wire [2:0] coupler_to_bus_named_cbus__EVAL_35;
  wire  coupler_to_bus_named_cbus__EVAL_36;
  wire [3:0] coupler_to_bus_named_cbus__EVAL_37;
  wire [2:0] coupler_to_bus_named_cbus__EVAL_38;
  wire [2:0] coupler_to_bus_named_cbus__EVAL_39;
  wire [2:0] coupler_to_bus_named_cbus__EVAL_40;
  wire  coupler_to_bus_named_cbus__EVAL_41;
  wire [3:0] coupler_to_bus_named_cbus__EVAL_42;
  wire  coupler_to_bus_named_cbus__EVAL_43;
  wire  coupler_to_bus_named_cbus__EVAL_44;
  wire  coupler_to_bus_named_cbus__EVAL_45;
  wire  coupler_to_bus_named_cbus__EVAL_46;
  wire  coupler_to_bus_named_cbus__EVAL_47;
  wire [29:0] coupler_to_bus_named_cbus__EVAL_48;
  wire [3:0] coupler_to_bus_named_cbus__EVAL_49;
  wire [2:0] coupler_to_bus_named_cbus__EVAL_50;
  wire [31:0] coupler_to_bus_named_cbus__EVAL_51;
  wire  coupler_to_bus_named_cbus__EVAL_52;
  wire  coupler_to_bus_named_cbus__EVAL_53;
  wire [1:0] coupler_to_bus_named_cbus__EVAL_54;
  wire  coupler_from_bus_named_front_bus__EVAL;
  wire [1:0] coupler_from_bus_named_front_bus__EVAL_0;
  wire  coupler_from_bus_named_front_bus__EVAL_1;
  wire [31:0] coupler_from_bus_named_front_bus__EVAL_2;
  wire  coupler_from_bus_named_front_bus__EVAL_3;
  wire [2:0] coupler_from_bus_named_front_bus__EVAL_4;
  wire  coupler_from_bus_named_front_bus__EVAL_5;
  wire  coupler_from_bus_named_front_bus__EVAL_6;
  wire [3:0] coupler_from_bus_named_front_bus__EVAL_7;
  wire [31:0] coupler_from_bus_named_front_bus__EVAL_8;
  wire  coupler_from_bus_named_front_bus__EVAL_9;
  wire [31:0] coupler_from_bus_named_front_bus__EVAL_10;
  wire  coupler_from_bus_named_front_bus__EVAL_11;
  wire  coupler_from_bus_named_front_bus__EVAL_12;
  wire  coupler_from_bus_named_front_bus__EVAL_13;
  wire  coupler_from_bus_named_front_bus__EVAL_14;
  wire  coupler_from_bus_named_front_bus__EVAL_15;
  wire [3:0] coupler_from_bus_named_front_bus__EVAL_16;
  wire  coupler_from_bus_named_front_bus__EVAL_17;
  wire  coupler_from_bus_named_front_bus__EVAL_18;
  wire [2:0] coupler_from_bus_named_front_bus__EVAL_19;
  wire  coupler_from_bus_named_front_bus__EVAL_20;
  wire [3:0] coupler_from_bus_named_front_bus__EVAL_21;
  wire [2:0] coupler_from_bus_named_front_bus__EVAL_22;
  wire  coupler_from_bus_named_front_bus__EVAL_23;
  wire  coupler_from_bus_named_front_bus__EVAL_24;
  wire  coupler_from_bus_named_front_bus__EVAL_25;
  wire [2:0] coupler_from_bus_named_front_bus__EVAL_26;
  wire [31:0] coupler_from_bus_named_front_bus__EVAL_27;
  wire  coupler_from_bus_named_front_bus__EVAL_28;
  wire  coupler_from_bus_named_front_bus__EVAL_29;
  wire  coupler_from_bus_named_front_bus__EVAL_30;
  wire  coupler_from_bus_named_front_bus__EVAL_31;
  wire  coupler_from_bus_named_front_bus__EVAL_32;
  wire [31:0] coupler_from_bus_named_front_bus__EVAL_33;
  wire  coupler_from_bus_named_front_bus__EVAL_34;
  wire  coupler_from_bus_named_front_bus__EVAL_35;
  wire [2:0] coupler_from_bus_named_front_bus__EVAL_36;
  wire  coupler_from_bus_named_front_bus__EVAL_37;
  wire  coupler_from_bus_named_front_bus__EVAL_38;
  wire  coupler_from_bus_named_front_bus__EVAL_39;
  wire [3:0] coupler_from_bus_named_front_bus__EVAL_40;
  wire [3:0] coupler_from_bus_named_front_bus__EVAL_41;
  wire  coupler_from_bus_named_front_bus__EVAL_42;
  wire  coupler_from_bus_named_front_bus__EVAL_43;
  wire [3:0] coupler_from_bus_named_front_bus__EVAL_44;
  wire  coupler_from_bus_named_front_bus__EVAL_45;
  wire [1:0] coupler_from_bus_named_front_bus__EVAL_46;
  wire  coupler_from_bus_named_front_bus__EVAL_47;
  wire  coupler_from_bus_named_front_bus__EVAL_48;
  wire  coupler_from_bus_named_front_bus__EVAL_49;
  wire [31:0] coupler_from_bus_named_front_bus__EVAL_50;
  wire  coupler_from_bus_named_front_bus__EVAL_51;
  wire [2:0] coupler_from_bus_named_front_bus__EVAL_52;
  wire  coupler_from_tile_with_no_name__EVAL;
  wire  coupler_from_tile_with_no_name__EVAL_0;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_1;
  wire  coupler_from_tile_with_no_name__EVAL_2;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_3;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_4;
  wire  coupler_from_tile_with_no_name__EVAL_5;
  wire  coupler_from_tile_with_no_name__EVAL_6;
  wire  coupler_from_tile_with_no_name__EVAL_7;
  wire  coupler_from_tile_with_no_name__EVAL_8;
  wire  coupler_from_tile_with_no_name__EVAL_9;
  wire  coupler_from_tile_with_no_name__EVAL_10;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_11;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_12;
  wire  coupler_from_tile_with_no_name__EVAL_13;
  wire  coupler_from_tile_with_no_name__EVAL_14;
  wire  coupler_from_tile_with_no_name__EVAL_15;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_16;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_17;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_18;
  wire  coupler_from_tile_with_no_name__EVAL_19;
  wire  coupler_from_tile_with_no_name__EVAL_20;
  wire  coupler_from_tile_with_no_name__EVAL_21;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_22;
  wire  coupler_from_tile_with_no_name__EVAL_23;
  wire  coupler_from_tile_with_no_name__EVAL_24;
  wire  coupler_from_tile_with_no_name__EVAL_25;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_26;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_27;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_28;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_29;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_30;
  wire  coupler_from_tile_with_no_name__EVAL_31;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_32;
  wire  coupler_from_tile_with_no_name__EVAL_33;
  wire  coupler_from_tile_with_no_name__EVAL_34;
  wire  coupler_from_tile_with_no_name__EVAL_35;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_36;
  wire  coupler_from_tile_with_no_name__EVAL_37;
  wire  coupler_from_tile_with_no_name__EVAL_38;
  wire  coupler_from_tile_with_no_name__EVAL_39;
  wire  coupler_from_tile_with_no_name__EVAL_40;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_41;
  wire  coupler_from_tile_with_no_name__EVAL_42;
  wire  coupler_from_tile_with_no_name__EVAL_43;
  wire  coupler_from_tile_with_no_name__EVAL_44;
  wire  coupler_from_tile_with_no_name__EVAL_45;
  wire  coupler_from_tile_with_no_name__EVAL_46;
  wire  coupler_from_tile_with_no_name__EVAL_47;
  wire  coupler_from_tile_with_no_name__EVAL_48;
  wire  coupler_from_tile_with_no_name__EVAL_49;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_50;
  wire  coupler_from_tile_with_no_name__EVAL_51;
  wire  coupler_from_tile_with_no_name__EVAL_52;
  wire  coupler_from_tile_with_no_name__EVAL_53;
  wire  coupler_from_tile_with_no_name__EVAL_54;
  wire  coupler_from_tile_with_no_name__EVAL_55;
  wire  coupler_from_tile_with_no_name__EVAL_56;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_57;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_58;
  wire  coupler_from_tile_with_no_name__EVAL_59;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_60;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_61;
  wire  coupler_from_tile_with_no_name__EVAL_62;
  wire  coupler_from_tile_with_no_name__EVAL_63;
  wire  coupler_from_tile_with_no_name__EVAL_64;
  wire  coupler_from_tile_with_no_name__EVAL_65;
  wire  coupler_from_tile_with_no_name__EVAL_66;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_67;
  wire  coupler_from_tile_with_no_name__EVAL_68;
  wire  coupler_from_tile_with_no_name__EVAL_69;
  wire  coupler_from_tile_with_no_name__EVAL_70;
  wire [1:0] coupler_from_tile_with_no_name__EVAL_71;
  wire  coupler_from_tile_with_no_name__EVAL_72;
  wire  coupler_from_tile_with_no_name__EVAL_73;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_74;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_75;
  wire  coupler_from_tile_with_no_name__EVAL_76;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_77;
  wire  coupler_from_tile_with_no_name__EVAL_78;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_79;
  wire  coupler_from_tile_with_no_name__EVAL_80;
  wire  coupler_from_tile_with_no_name__EVAL_81;
  wire  coupler_from_tile_with_no_name__EVAL_82;
  wire  coupler_from_tile_with_no_name__EVAL_83;
  wire  coupler_from_tile_with_no_name__EVAL_84;
  wire  coupler_from_tile_with_no_name__EVAL_85;
  wire  coupler_from_tile_with_no_name__EVAL_86;
  wire  coupler_from_tile_with_no_name__EVAL_87;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_88;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_89;
  wire  coupler_from_tile_with_no_name__EVAL_90;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_91;
  wire  coupler_from_tile_with_no_name__EVAL_92;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_93;
  wire  coupler_from_tile_with_no_name__EVAL_94;
  wire  coupler_from_tile_with_no_name__EVAL_95;
  wire  coupler_from_tile_with_no_name__EVAL_96;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_97;
  wire  coupler_from_tile_with_no_name__EVAL_98;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_99;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_100;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_101;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_102;
  wire  coupler_from_tile_with_no_name__EVAL_103;
  wire [31:0] coupler_from_tile_with_no_name__EVAL_104;
  wire  coupler_from_tile_with_no_name__EVAL_105;
  wire  coupler_from_tile_with_no_name__EVAL_106;
  wire [3:0] coupler_from_tile_with_no_name__EVAL_107;
  wire [2:0] coupler_from_tile_with_no_name__EVAL_108;
  wire [3:0] coupler_to_sys_sram_1__EVAL;
  wire [2:0] coupler_to_sys_sram_1__EVAL_0;
  wire  coupler_to_sys_sram_1__EVAL_1;
  wire [31:0] coupler_to_sys_sram_1__EVAL_2;
  wire  coupler_to_sys_sram_1__EVAL_3;
  wire  coupler_to_sys_sram_1__EVAL_4;
  wire [31:0] coupler_to_sys_sram_1__EVAL_5;
  wire [1:0] coupler_to_sys_sram_1__EVAL_6;
  wire [31:0] coupler_to_sys_sram_1__EVAL_7;
  wire [31:0] coupler_to_sys_sram_1__EVAL_8;
  wire [2:0] coupler_to_sys_sram_1__EVAL_9;
  wire  coupler_to_sys_sram_1__EVAL_10;
  wire [2:0] coupler_to_sys_sram_1__EVAL_11;
  wire  coupler_to_sys_sram_1__EVAL_12;
  wire [2:0] coupler_to_sys_sram_1__EVAL_13;
  wire [2:0] coupler_to_sys_sram_1__EVAL_14;
  wire [1:0] coupler_to_sys_sram_1__EVAL_15;
  wire [2:0] coupler_to_sys_sram_1__EVAL_16;
  wire [3:0] coupler_to_sys_sram_1__EVAL_17;
  wire [31:0] coupler_to_sys_sram_1__EVAL_18;
  wire [2:0] coupler_to_sys_sram_1__EVAL_19;
  wire  coupler_to_sys_sram_1__EVAL_20;
  wire  coupler_to_sys_sram_1__EVAL_21;
  wire  coupler_to_sys_sram_1__EVAL_22;
  wire  coupler_to_sys_sram_1__EVAL_23;
  wire  coupler_to_sys_sram_1__EVAL_24;
  wire [1:0] coupler_to_sys_sram_1__EVAL_25;
  wire  coupler_to_sys_sram_1__EVAL_26;
  wire  coupler_to_sys_sram_1__EVAL_27;
  wire [2:0] coupler_to_sys_sram_1__EVAL_28;
  wire [31:0] coupler_to_sys_sram_1__EVAL_29;
  wire [2:0] coupler_to_sys_sram_1__EVAL_30;
  wire [1:0] coupler_to_sys_sram_1__EVAL_31;
  wire [2:0] coupler_to_sys_sram_1__EVAL_32;
  wire  system_bus_clock_groups__EVAL_1;
  wire  system_bus_clock_groups__EVAL_2;
  wire  system_bus_clock_groups__EVAL_3;
  wire  system_bus_clock_groups__EVAL_4;
  wire  system_bus_clock_groups__EVAL_7;
  wire  system_bus_clock_groups__EVAL_10;
  wire  system_bus_clock_groups__EVAL_11;
  wire  system_bus_clock_groups__EVAL_12;
  wire  system_bus_clock_groups__EVAL_15;
  wire  system_bus_clock_groups__EVAL_17;
  wire  system_bus_clock_groups__EVAL_19;
  wire  system_bus_clock_groups__EVAL_22;
  wire  coupler_to_port_named_ahb_sys_port__EVAL;
  wire [31:0] coupler_to_port_named_ahb_sys_port__EVAL_0;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_1;
  wire [2:0] coupler_to_port_named_ahb_sys_port__EVAL_2;
  wire [2:0] coupler_to_port_named_ahb_sys_port__EVAL_3;
  wire [1:0] coupler_to_port_named_ahb_sys_port__EVAL_4;
  wire [2:0] coupler_to_port_named_ahb_sys_port__EVAL_5;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_6;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_7;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_8;
  wire [2:0] coupler_to_port_named_ahb_sys_port__EVAL_9;
  wire [31:0] coupler_to_port_named_ahb_sys_port__EVAL_10;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_11;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_12;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_13;
  wire [1:0] coupler_to_port_named_ahb_sys_port__EVAL_14;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_15;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_16;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_17;
  wire [31:0] coupler_to_port_named_ahb_sys_port__EVAL_18;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_19;
  wire [30:0] coupler_to_port_named_ahb_sys_port__EVAL_20;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_21;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_22;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_23;
  wire [31:0] coupler_to_port_named_ahb_sys_port__EVAL_24;
  wire [2:0] coupler_to_port_named_ahb_sys_port__EVAL_25;
  wire [3:0] coupler_to_port_named_ahb_sys_port__EVAL_26;
  wire [2:0] coupler_to_port_named_ahb_sys_port__EVAL_27;
  wire [30:0] coupler_to_port_named_ahb_sys_port__EVAL_28;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_29;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_30;
  wire [2:0] coupler_to_port_named_ahb_sys_port__EVAL_31;
  wire [2:0] coupler_to_port_named_ahb_sys_port__EVAL_32;
  wire [2:0] coupler_to_port_named_ahb_sys_port__EVAL_33;
  wire [3:0] coupler_to_port_named_ahb_sys_port__EVAL_34;
  wire [31:0] coupler_to_sys_sram_0__EVAL;
  wire  coupler_to_sys_sram_0__EVAL_0;
  wire [31:0] coupler_to_sys_sram_0__EVAL_1;
  wire [1:0] coupler_to_sys_sram_0__EVAL_2;
  wire [31:0] coupler_to_sys_sram_0__EVAL_3;
  wire  coupler_to_sys_sram_0__EVAL_4;
  wire  coupler_to_sys_sram_0__EVAL_5;
  wire [31:0] coupler_to_sys_sram_0__EVAL_6;
  wire [2:0] coupler_to_sys_sram_0__EVAL_7;
  wire [2:0] coupler_to_sys_sram_0__EVAL_8;
  wire  coupler_to_sys_sram_0__EVAL_9;
  wire  coupler_to_sys_sram_0__EVAL_10;
  wire [2:0] coupler_to_sys_sram_0__EVAL_11;
  wire [3:0] coupler_to_sys_sram_0__EVAL_12;
  wire  coupler_to_sys_sram_0__EVAL_13;
  wire [1:0] coupler_to_sys_sram_0__EVAL_14;
  wire  coupler_to_sys_sram_0__EVAL_15;
  wire [2:0] coupler_to_sys_sram_0__EVAL_16;
  wire [2:0] coupler_to_sys_sram_0__EVAL_17;
  wire [2:0] coupler_to_sys_sram_0__EVAL_18;
  wire [3:0] coupler_to_sys_sram_0__EVAL_19;
  wire  coupler_to_sys_sram_0__EVAL_20;
  wire  coupler_to_sys_sram_0__EVAL_21;
  wire [1:0] coupler_to_sys_sram_0__EVAL_22;
  wire [2:0] coupler_to_sys_sram_0__EVAL_23;
  wire  coupler_to_sys_sram_0__EVAL_24;
  wire [1:0] coupler_to_sys_sram_0__EVAL_25;
  wire  coupler_to_sys_sram_0__EVAL_26;
  wire  coupler_to_sys_sram_0__EVAL_27;
  wire [2:0] coupler_to_sys_sram_0__EVAL_28;
  wire [2:0] coupler_to_sys_sram_0__EVAL_29;
  wire [2:0] coupler_to_sys_sram_0__EVAL_30;
  wire [31:0] coupler_to_sys_sram_0__EVAL_31;
  wire [31:0] coupler_to_sys_sram_0__EVAL_32;
  wire  clockGroup__EVAL;
  wire  clockGroup__EVAL_0;
  wire  clockGroup__EVAL_1;
  wire  clockGroup__EVAL_2;
  _EVAL_4 system_bus_xbar (
    ._EVAL(system_bus_xbar__EVAL),
    ._EVAL_0(system_bus_xbar__EVAL_0),
    ._EVAL_1(system_bus_xbar__EVAL_1),
    ._EVAL_2(system_bus_xbar__EVAL_2),
    ._EVAL_3(system_bus_xbar__EVAL_3),
    ._EVAL_4(system_bus_xbar__EVAL_4),
    ._EVAL_5(system_bus_xbar__EVAL_5),
    ._EVAL_6(system_bus_xbar__EVAL_6),
    ._EVAL_7(system_bus_xbar__EVAL_7),
    ._EVAL_8(system_bus_xbar__EVAL_8),
    ._EVAL_9(system_bus_xbar__EVAL_9),
    ._EVAL_10(system_bus_xbar__EVAL_10),
    ._EVAL_11(system_bus_xbar__EVAL_11),
    ._EVAL_12(system_bus_xbar__EVAL_12),
    ._EVAL_13(system_bus_xbar__EVAL_13),
    ._EVAL_14(system_bus_xbar__EVAL_14),
    ._EVAL_15(system_bus_xbar__EVAL_15),
    ._EVAL_16(system_bus_xbar__EVAL_16),
    ._EVAL_17(system_bus_xbar__EVAL_17),
    ._EVAL_18(system_bus_xbar__EVAL_18),
    ._EVAL_19(system_bus_xbar__EVAL_19),
    ._EVAL_20(system_bus_xbar__EVAL_20),
    ._EVAL_21(system_bus_xbar__EVAL_21),
    ._EVAL_22(system_bus_xbar__EVAL_22),
    ._EVAL_23(system_bus_xbar__EVAL_23),
    ._EVAL_24(system_bus_xbar__EVAL_24),
    ._EVAL_25(system_bus_xbar__EVAL_25),
    ._EVAL_26(system_bus_xbar__EVAL_26),
    ._EVAL_27(system_bus_xbar__EVAL_27),
    ._EVAL_28(system_bus_xbar__EVAL_28),
    ._EVAL_29(system_bus_xbar__EVAL_29),
    ._EVAL_30(system_bus_xbar__EVAL_30),
    ._EVAL_31(system_bus_xbar__EVAL_31),
    ._EVAL_32(system_bus_xbar__EVAL_32),
    ._EVAL_33(system_bus_xbar__EVAL_33),
    ._EVAL_34(system_bus_xbar__EVAL_34),
    ._EVAL_35(system_bus_xbar__EVAL_35),
    ._EVAL_36(system_bus_xbar__EVAL_36),
    ._EVAL_37(system_bus_xbar__EVAL_37),
    ._EVAL_38(system_bus_xbar__EVAL_38),
    ._EVAL_39(system_bus_xbar__EVAL_39),
    ._EVAL_40(system_bus_xbar__EVAL_40),
    ._EVAL_41(system_bus_xbar__EVAL_41),
    ._EVAL_42(system_bus_xbar__EVAL_42),
    ._EVAL_43(system_bus_xbar__EVAL_43),
    ._EVAL_44(system_bus_xbar__EVAL_44),
    ._EVAL_45(system_bus_xbar__EVAL_45),
    ._EVAL_46(system_bus_xbar__EVAL_46),
    ._EVAL_47(system_bus_xbar__EVAL_47),
    ._EVAL_48(system_bus_xbar__EVAL_48),
    ._EVAL_49(system_bus_xbar__EVAL_49),
    ._EVAL_50(system_bus_xbar__EVAL_50),
    ._EVAL_51(system_bus_xbar__EVAL_51),
    ._EVAL_52(system_bus_xbar__EVAL_52),
    ._EVAL_53(system_bus_xbar__EVAL_53),
    ._EVAL_54(system_bus_xbar__EVAL_54),
    ._EVAL_55(system_bus_xbar__EVAL_55),
    ._EVAL_56(system_bus_xbar__EVAL_56),
    ._EVAL_57(system_bus_xbar__EVAL_57),
    ._EVAL_58(system_bus_xbar__EVAL_58),
    ._EVAL_59(system_bus_xbar__EVAL_59),
    ._EVAL_60(system_bus_xbar__EVAL_60),
    ._EVAL_61(system_bus_xbar__EVAL_61),
    ._EVAL_62(system_bus_xbar__EVAL_62),
    ._EVAL_63(system_bus_xbar__EVAL_63),
    ._EVAL_64(system_bus_xbar__EVAL_64),
    ._EVAL_65(system_bus_xbar__EVAL_65),
    ._EVAL_66(system_bus_xbar__EVAL_66),
    ._EVAL_67(system_bus_xbar__EVAL_67),
    ._EVAL_68(system_bus_xbar__EVAL_68),
    ._EVAL_69(system_bus_xbar__EVAL_69),
    ._EVAL_70(system_bus_xbar__EVAL_70),
    ._EVAL_71(system_bus_xbar__EVAL_71),
    ._EVAL_72(system_bus_xbar__EVAL_72),
    ._EVAL_73(system_bus_xbar__EVAL_73),
    ._EVAL_74(system_bus_xbar__EVAL_74),
    ._EVAL_75(system_bus_xbar__EVAL_75),
    ._EVAL_76(system_bus_xbar__EVAL_76),
    ._EVAL_77(system_bus_xbar__EVAL_77),
    ._EVAL_78(system_bus_xbar__EVAL_78),
    ._EVAL_79(system_bus_xbar__EVAL_79),
    ._EVAL_80(system_bus_xbar__EVAL_80),
    ._EVAL_81(system_bus_xbar__EVAL_81),
    ._EVAL_82(system_bus_xbar__EVAL_82),
    ._EVAL_83(system_bus_xbar__EVAL_83),
    ._EVAL_84(system_bus_xbar__EVAL_84),
    ._EVAL_85(system_bus_xbar__EVAL_85),
    ._EVAL_86(system_bus_xbar__EVAL_86),
    ._EVAL_87(system_bus_xbar__EVAL_87),
    ._EVAL_88(system_bus_xbar__EVAL_88),
    ._EVAL_89(system_bus_xbar__EVAL_89),
    ._EVAL_90(system_bus_xbar__EVAL_90),
    ._EVAL_91(system_bus_xbar__EVAL_91),
    ._EVAL_92(system_bus_xbar__EVAL_92),
    ._EVAL_93(system_bus_xbar__EVAL_93),
    ._EVAL_94(system_bus_xbar__EVAL_94),
    ._EVAL_95(system_bus_xbar__EVAL_95),
    ._EVAL_96(system_bus_xbar__EVAL_96),
    ._EVAL_97(system_bus_xbar__EVAL_97),
    ._EVAL_98(system_bus_xbar__EVAL_98),
    ._EVAL_99(system_bus_xbar__EVAL_99),
    ._EVAL_100(system_bus_xbar__EVAL_100),
    ._EVAL_101(system_bus_xbar__EVAL_101),
    ._EVAL_102(system_bus_xbar__EVAL_102),
    ._EVAL_103(system_bus_xbar__EVAL_103),
    ._EVAL_104(system_bus_xbar__EVAL_104),
    ._EVAL_105(system_bus_xbar__EVAL_105),
    ._EVAL_106(system_bus_xbar__EVAL_106),
    ._EVAL_107(system_bus_xbar__EVAL_107),
    ._EVAL_108(system_bus_xbar__EVAL_108),
    ._EVAL_109(system_bus_xbar__EVAL_109),
    ._EVAL_110(system_bus_xbar__EVAL_110),
    ._EVAL_111(system_bus_xbar__EVAL_111),
    ._EVAL_112(system_bus_xbar__EVAL_112),
    ._EVAL_113(system_bus_xbar__EVAL_113),
    ._EVAL_114(system_bus_xbar__EVAL_114),
    ._EVAL_115(system_bus_xbar__EVAL_115),
    ._EVAL_116(system_bus_xbar__EVAL_116),
    ._EVAL_117(system_bus_xbar__EVAL_117),
    ._EVAL_118(system_bus_xbar__EVAL_118),
    ._EVAL_119(system_bus_xbar__EVAL_119),
    ._EVAL_120(system_bus_xbar__EVAL_120),
    ._EVAL_121(system_bus_xbar__EVAL_121),
    ._EVAL_122(system_bus_xbar__EVAL_122),
    ._EVAL_123(system_bus_xbar__EVAL_123),
    ._EVAL_124(system_bus_xbar__EVAL_124),
    ._EVAL_125(system_bus_xbar__EVAL_125),
    ._EVAL_126(system_bus_xbar__EVAL_126),
    ._EVAL_127(system_bus_xbar__EVAL_127),
    ._EVAL_128(system_bus_xbar__EVAL_128),
    ._EVAL_129(system_bus_xbar__EVAL_129),
    ._EVAL_130(system_bus_xbar__EVAL_130),
    ._EVAL_131(system_bus_xbar__EVAL_131),
    ._EVAL_132(system_bus_xbar__EVAL_132),
    ._EVAL_133(system_bus_xbar__EVAL_133),
    ._EVAL_134(system_bus_xbar__EVAL_134),
    ._EVAL_135(system_bus_xbar__EVAL_135),
    ._EVAL_136(system_bus_xbar__EVAL_136),
    ._EVAL_137(system_bus_xbar__EVAL_137),
    ._EVAL_138(system_bus_xbar__EVAL_138),
    ._EVAL_139(system_bus_xbar__EVAL_139),
    ._EVAL_140(system_bus_xbar__EVAL_140),
    ._EVAL_141(system_bus_xbar__EVAL_141),
    ._EVAL_142(system_bus_xbar__EVAL_142),
    ._EVAL_143(system_bus_xbar__EVAL_143),
    ._EVAL_144(system_bus_xbar__EVAL_144),
    ._EVAL_145(system_bus_xbar__EVAL_145),
    ._EVAL_146(system_bus_xbar__EVAL_146),
    ._EVAL_147(system_bus_xbar__EVAL_147),
    ._EVAL_148(system_bus_xbar__EVAL_148),
    ._EVAL_149(system_bus_xbar__EVAL_149),
    ._EVAL_150(system_bus_xbar__EVAL_150),
    ._EVAL_151(system_bus_xbar__EVAL_151),
    ._EVAL_152(system_bus_xbar__EVAL_152),
    ._EVAL_153(system_bus_xbar__EVAL_153),
    ._EVAL_154(system_bus_xbar__EVAL_154),
    ._EVAL_155(system_bus_xbar__EVAL_155),
    ._EVAL_156(system_bus_xbar__EVAL_156),
    ._EVAL_157(system_bus_xbar__EVAL_157),
    ._EVAL_158(system_bus_xbar__EVAL_158),
    ._EVAL_159(system_bus_xbar__EVAL_159),
    ._EVAL_160(system_bus_xbar__EVAL_160),
    ._EVAL_161(system_bus_xbar__EVAL_161),
    ._EVAL_162(system_bus_xbar__EVAL_162),
    ._EVAL_163(system_bus_xbar__EVAL_163)
  );
  _EVAL_1 fixedClockNode (
    ._EVAL(fixedClockNode__EVAL),
    ._EVAL_0(fixedClockNode__EVAL_0),
    ._EVAL_1(fixedClockNode__EVAL_1),
    ._EVAL_2(fixedClockNode__EVAL_2)
  );
  _EVAL_33 coupler_to_bus_named_cbus (
    ._EVAL(coupler_to_bus_named_cbus__EVAL),
    ._EVAL_0(coupler_to_bus_named_cbus__EVAL_0),
    ._EVAL_1(coupler_to_bus_named_cbus__EVAL_1),
    ._EVAL_2(coupler_to_bus_named_cbus__EVAL_2),
    ._EVAL_3(coupler_to_bus_named_cbus__EVAL_3),
    ._EVAL_4(coupler_to_bus_named_cbus__EVAL_4),
    ._EVAL_5(coupler_to_bus_named_cbus__EVAL_5),
    ._EVAL_6(coupler_to_bus_named_cbus__EVAL_6),
    ._EVAL_7(coupler_to_bus_named_cbus__EVAL_7),
    ._EVAL_8(coupler_to_bus_named_cbus__EVAL_8),
    ._EVAL_9(coupler_to_bus_named_cbus__EVAL_9),
    ._EVAL_10(coupler_to_bus_named_cbus__EVAL_10),
    ._EVAL_11(coupler_to_bus_named_cbus__EVAL_11),
    ._EVAL_12(coupler_to_bus_named_cbus__EVAL_12),
    ._EVAL_13(coupler_to_bus_named_cbus__EVAL_13),
    ._EVAL_14(coupler_to_bus_named_cbus__EVAL_14),
    ._EVAL_15(coupler_to_bus_named_cbus__EVAL_15),
    ._EVAL_16(coupler_to_bus_named_cbus__EVAL_16),
    ._EVAL_17(coupler_to_bus_named_cbus__EVAL_17),
    ._EVAL_18(coupler_to_bus_named_cbus__EVAL_18),
    ._EVAL_19(coupler_to_bus_named_cbus__EVAL_19),
    ._EVAL_20(coupler_to_bus_named_cbus__EVAL_20),
    ._EVAL_21(coupler_to_bus_named_cbus__EVAL_21),
    ._EVAL_22(coupler_to_bus_named_cbus__EVAL_22),
    ._EVAL_23(coupler_to_bus_named_cbus__EVAL_23),
    ._EVAL_24(coupler_to_bus_named_cbus__EVAL_24),
    ._EVAL_25(coupler_to_bus_named_cbus__EVAL_25),
    ._EVAL_26(coupler_to_bus_named_cbus__EVAL_26),
    ._EVAL_27(coupler_to_bus_named_cbus__EVAL_27),
    ._EVAL_28(coupler_to_bus_named_cbus__EVAL_28),
    ._EVAL_29(coupler_to_bus_named_cbus__EVAL_29),
    ._EVAL_30(coupler_to_bus_named_cbus__EVAL_30),
    ._EVAL_31(coupler_to_bus_named_cbus__EVAL_31),
    ._EVAL_32(coupler_to_bus_named_cbus__EVAL_32),
    ._EVAL_33(coupler_to_bus_named_cbus__EVAL_33),
    ._EVAL_34(coupler_to_bus_named_cbus__EVAL_34),
    ._EVAL_35(coupler_to_bus_named_cbus__EVAL_35),
    ._EVAL_36(coupler_to_bus_named_cbus__EVAL_36),
    ._EVAL_37(coupler_to_bus_named_cbus__EVAL_37),
    ._EVAL_38(coupler_to_bus_named_cbus__EVAL_38),
    ._EVAL_39(coupler_to_bus_named_cbus__EVAL_39),
    ._EVAL_40(coupler_to_bus_named_cbus__EVAL_40),
    ._EVAL_41(coupler_to_bus_named_cbus__EVAL_41),
    ._EVAL_42(coupler_to_bus_named_cbus__EVAL_42),
    ._EVAL_43(coupler_to_bus_named_cbus__EVAL_43),
    ._EVAL_44(coupler_to_bus_named_cbus__EVAL_44),
    ._EVAL_45(coupler_to_bus_named_cbus__EVAL_45),
    ._EVAL_46(coupler_to_bus_named_cbus__EVAL_46),
    ._EVAL_47(coupler_to_bus_named_cbus__EVAL_47),
    ._EVAL_48(coupler_to_bus_named_cbus__EVAL_48),
    ._EVAL_49(coupler_to_bus_named_cbus__EVAL_49),
    ._EVAL_50(coupler_to_bus_named_cbus__EVAL_50),
    ._EVAL_51(coupler_to_bus_named_cbus__EVAL_51),
    ._EVAL_52(coupler_to_bus_named_cbus__EVAL_52),
    ._EVAL_53(coupler_to_bus_named_cbus__EVAL_53),
    ._EVAL_54(coupler_to_bus_named_cbus__EVAL_54)
  );
  _EVAL_36 coupler_from_bus_named_front_bus (
    ._EVAL(coupler_from_bus_named_front_bus__EVAL),
    ._EVAL_0(coupler_from_bus_named_front_bus__EVAL_0),
    ._EVAL_1(coupler_from_bus_named_front_bus__EVAL_1),
    ._EVAL_2(coupler_from_bus_named_front_bus__EVAL_2),
    ._EVAL_3(coupler_from_bus_named_front_bus__EVAL_3),
    ._EVAL_4(coupler_from_bus_named_front_bus__EVAL_4),
    ._EVAL_5(coupler_from_bus_named_front_bus__EVAL_5),
    ._EVAL_6(coupler_from_bus_named_front_bus__EVAL_6),
    ._EVAL_7(coupler_from_bus_named_front_bus__EVAL_7),
    ._EVAL_8(coupler_from_bus_named_front_bus__EVAL_8),
    ._EVAL_9(coupler_from_bus_named_front_bus__EVAL_9),
    ._EVAL_10(coupler_from_bus_named_front_bus__EVAL_10),
    ._EVAL_11(coupler_from_bus_named_front_bus__EVAL_11),
    ._EVAL_12(coupler_from_bus_named_front_bus__EVAL_12),
    ._EVAL_13(coupler_from_bus_named_front_bus__EVAL_13),
    ._EVAL_14(coupler_from_bus_named_front_bus__EVAL_14),
    ._EVAL_15(coupler_from_bus_named_front_bus__EVAL_15),
    ._EVAL_16(coupler_from_bus_named_front_bus__EVAL_16),
    ._EVAL_17(coupler_from_bus_named_front_bus__EVAL_17),
    ._EVAL_18(coupler_from_bus_named_front_bus__EVAL_18),
    ._EVAL_19(coupler_from_bus_named_front_bus__EVAL_19),
    ._EVAL_20(coupler_from_bus_named_front_bus__EVAL_20),
    ._EVAL_21(coupler_from_bus_named_front_bus__EVAL_21),
    ._EVAL_22(coupler_from_bus_named_front_bus__EVAL_22),
    ._EVAL_23(coupler_from_bus_named_front_bus__EVAL_23),
    ._EVAL_24(coupler_from_bus_named_front_bus__EVAL_24),
    ._EVAL_25(coupler_from_bus_named_front_bus__EVAL_25),
    ._EVAL_26(coupler_from_bus_named_front_bus__EVAL_26),
    ._EVAL_27(coupler_from_bus_named_front_bus__EVAL_27),
    ._EVAL_28(coupler_from_bus_named_front_bus__EVAL_28),
    ._EVAL_29(coupler_from_bus_named_front_bus__EVAL_29),
    ._EVAL_30(coupler_from_bus_named_front_bus__EVAL_30),
    ._EVAL_31(coupler_from_bus_named_front_bus__EVAL_31),
    ._EVAL_32(coupler_from_bus_named_front_bus__EVAL_32),
    ._EVAL_33(coupler_from_bus_named_front_bus__EVAL_33),
    ._EVAL_34(coupler_from_bus_named_front_bus__EVAL_34),
    ._EVAL_35(coupler_from_bus_named_front_bus__EVAL_35),
    ._EVAL_36(coupler_from_bus_named_front_bus__EVAL_36),
    ._EVAL_37(coupler_from_bus_named_front_bus__EVAL_37),
    ._EVAL_38(coupler_from_bus_named_front_bus__EVAL_38),
    ._EVAL_39(coupler_from_bus_named_front_bus__EVAL_39),
    ._EVAL_40(coupler_from_bus_named_front_bus__EVAL_40),
    ._EVAL_41(coupler_from_bus_named_front_bus__EVAL_41),
    ._EVAL_42(coupler_from_bus_named_front_bus__EVAL_42),
    ._EVAL_43(coupler_from_bus_named_front_bus__EVAL_43),
    ._EVAL_44(coupler_from_bus_named_front_bus__EVAL_44),
    ._EVAL_45(coupler_from_bus_named_front_bus__EVAL_45),
    ._EVAL_46(coupler_from_bus_named_front_bus__EVAL_46),
    ._EVAL_47(coupler_from_bus_named_front_bus__EVAL_47),
    ._EVAL_48(coupler_from_bus_named_front_bus__EVAL_48),
    ._EVAL_49(coupler_from_bus_named_front_bus__EVAL_49),
    ._EVAL_50(coupler_from_bus_named_front_bus__EVAL_50),
    ._EVAL_51(coupler_from_bus_named_front_bus__EVAL_51),
    ._EVAL_52(coupler_from_bus_named_front_bus__EVAL_52)
  );
  _EVAL_9 coupler_from_tile_with_no_name (
    ._EVAL(coupler_from_tile_with_no_name__EVAL),
    ._EVAL_0(coupler_from_tile_with_no_name__EVAL_0),
    ._EVAL_1(coupler_from_tile_with_no_name__EVAL_1),
    ._EVAL_2(coupler_from_tile_with_no_name__EVAL_2),
    ._EVAL_3(coupler_from_tile_with_no_name__EVAL_3),
    ._EVAL_4(coupler_from_tile_with_no_name__EVAL_4),
    ._EVAL_5(coupler_from_tile_with_no_name__EVAL_5),
    ._EVAL_6(coupler_from_tile_with_no_name__EVAL_6),
    ._EVAL_7(coupler_from_tile_with_no_name__EVAL_7),
    ._EVAL_8(coupler_from_tile_with_no_name__EVAL_8),
    ._EVAL_9(coupler_from_tile_with_no_name__EVAL_9),
    ._EVAL_10(coupler_from_tile_with_no_name__EVAL_10),
    ._EVAL_11(coupler_from_tile_with_no_name__EVAL_11),
    ._EVAL_12(coupler_from_tile_with_no_name__EVAL_12),
    ._EVAL_13(coupler_from_tile_with_no_name__EVAL_13),
    ._EVAL_14(coupler_from_tile_with_no_name__EVAL_14),
    ._EVAL_15(coupler_from_tile_with_no_name__EVAL_15),
    ._EVAL_16(coupler_from_tile_with_no_name__EVAL_16),
    ._EVAL_17(coupler_from_tile_with_no_name__EVAL_17),
    ._EVAL_18(coupler_from_tile_with_no_name__EVAL_18),
    ._EVAL_19(coupler_from_tile_with_no_name__EVAL_19),
    ._EVAL_20(coupler_from_tile_with_no_name__EVAL_20),
    ._EVAL_21(coupler_from_tile_with_no_name__EVAL_21),
    ._EVAL_22(coupler_from_tile_with_no_name__EVAL_22),
    ._EVAL_23(coupler_from_tile_with_no_name__EVAL_23),
    ._EVAL_24(coupler_from_tile_with_no_name__EVAL_24),
    ._EVAL_25(coupler_from_tile_with_no_name__EVAL_25),
    ._EVAL_26(coupler_from_tile_with_no_name__EVAL_26),
    ._EVAL_27(coupler_from_tile_with_no_name__EVAL_27),
    ._EVAL_28(coupler_from_tile_with_no_name__EVAL_28),
    ._EVAL_29(coupler_from_tile_with_no_name__EVAL_29),
    ._EVAL_30(coupler_from_tile_with_no_name__EVAL_30),
    ._EVAL_31(coupler_from_tile_with_no_name__EVAL_31),
    ._EVAL_32(coupler_from_tile_with_no_name__EVAL_32),
    ._EVAL_33(coupler_from_tile_with_no_name__EVAL_33),
    ._EVAL_34(coupler_from_tile_with_no_name__EVAL_34),
    ._EVAL_35(coupler_from_tile_with_no_name__EVAL_35),
    ._EVAL_36(coupler_from_tile_with_no_name__EVAL_36),
    ._EVAL_37(coupler_from_tile_with_no_name__EVAL_37),
    ._EVAL_38(coupler_from_tile_with_no_name__EVAL_38),
    ._EVAL_39(coupler_from_tile_with_no_name__EVAL_39),
    ._EVAL_40(coupler_from_tile_with_no_name__EVAL_40),
    ._EVAL_41(coupler_from_tile_with_no_name__EVAL_41),
    ._EVAL_42(coupler_from_tile_with_no_name__EVAL_42),
    ._EVAL_43(coupler_from_tile_with_no_name__EVAL_43),
    ._EVAL_44(coupler_from_tile_with_no_name__EVAL_44),
    ._EVAL_45(coupler_from_tile_with_no_name__EVAL_45),
    ._EVAL_46(coupler_from_tile_with_no_name__EVAL_46),
    ._EVAL_47(coupler_from_tile_with_no_name__EVAL_47),
    ._EVAL_48(coupler_from_tile_with_no_name__EVAL_48),
    ._EVAL_49(coupler_from_tile_with_no_name__EVAL_49),
    ._EVAL_50(coupler_from_tile_with_no_name__EVAL_50),
    ._EVAL_51(coupler_from_tile_with_no_name__EVAL_51),
    ._EVAL_52(coupler_from_tile_with_no_name__EVAL_52),
    ._EVAL_53(coupler_from_tile_with_no_name__EVAL_53),
    ._EVAL_54(coupler_from_tile_with_no_name__EVAL_54),
    ._EVAL_55(coupler_from_tile_with_no_name__EVAL_55),
    ._EVAL_56(coupler_from_tile_with_no_name__EVAL_56),
    ._EVAL_57(coupler_from_tile_with_no_name__EVAL_57),
    ._EVAL_58(coupler_from_tile_with_no_name__EVAL_58),
    ._EVAL_59(coupler_from_tile_with_no_name__EVAL_59),
    ._EVAL_60(coupler_from_tile_with_no_name__EVAL_60),
    ._EVAL_61(coupler_from_tile_with_no_name__EVAL_61),
    ._EVAL_62(coupler_from_tile_with_no_name__EVAL_62),
    ._EVAL_63(coupler_from_tile_with_no_name__EVAL_63),
    ._EVAL_64(coupler_from_tile_with_no_name__EVAL_64),
    ._EVAL_65(coupler_from_tile_with_no_name__EVAL_65),
    ._EVAL_66(coupler_from_tile_with_no_name__EVAL_66),
    ._EVAL_67(coupler_from_tile_with_no_name__EVAL_67),
    ._EVAL_68(coupler_from_tile_with_no_name__EVAL_68),
    ._EVAL_69(coupler_from_tile_with_no_name__EVAL_69),
    ._EVAL_70(coupler_from_tile_with_no_name__EVAL_70),
    ._EVAL_71(coupler_from_tile_with_no_name__EVAL_71),
    ._EVAL_72(coupler_from_tile_with_no_name__EVAL_72),
    ._EVAL_73(coupler_from_tile_with_no_name__EVAL_73),
    ._EVAL_74(coupler_from_tile_with_no_name__EVAL_74),
    ._EVAL_75(coupler_from_tile_with_no_name__EVAL_75),
    ._EVAL_76(coupler_from_tile_with_no_name__EVAL_76),
    ._EVAL_77(coupler_from_tile_with_no_name__EVAL_77),
    ._EVAL_78(coupler_from_tile_with_no_name__EVAL_78),
    ._EVAL_79(coupler_from_tile_with_no_name__EVAL_79),
    ._EVAL_80(coupler_from_tile_with_no_name__EVAL_80),
    ._EVAL_81(coupler_from_tile_with_no_name__EVAL_81),
    ._EVAL_82(coupler_from_tile_with_no_name__EVAL_82),
    ._EVAL_83(coupler_from_tile_with_no_name__EVAL_83),
    ._EVAL_84(coupler_from_tile_with_no_name__EVAL_84),
    ._EVAL_85(coupler_from_tile_with_no_name__EVAL_85),
    ._EVAL_86(coupler_from_tile_with_no_name__EVAL_86),
    ._EVAL_87(coupler_from_tile_with_no_name__EVAL_87),
    ._EVAL_88(coupler_from_tile_with_no_name__EVAL_88),
    ._EVAL_89(coupler_from_tile_with_no_name__EVAL_89),
    ._EVAL_90(coupler_from_tile_with_no_name__EVAL_90),
    ._EVAL_91(coupler_from_tile_with_no_name__EVAL_91),
    ._EVAL_92(coupler_from_tile_with_no_name__EVAL_92),
    ._EVAL_93(coupler_from_tile_with_no_name__EVAL_93),
    ._EVAL_94(coupler_from_tile_with_no_name__EVAL_94),
    ._EVAL_95(coupler_from_tile_with_no_name__EVAL_95),
    ._EVAL_96(coupler_from_tile_with_no_name__EVAL_96),
    ._EVAL_97(coupler_from_tile_with_no_name__EVAL_97),
    ._EVAL_98(coupler_from_tile_with_no_name__EVAL_98),
    ._EVAL_99(coupler_from_tile_with_no_name__EVAL_99),
    ._EVAL_100(coupler_from_tile_with_no_name__EVAL_100),
    ._EVAL_101(coupler_from_tile_with_no_name__EVAL_101),
    ._EVAL_102(coupler_from_tile_with_no_name__EVAL_102),
    ._EVAL_103(coupler_from_tile_with_no_name__EVAL_103),
    ._EVAL_104(coupler_from_tile_with_no_name__EVAL_104),
    ._EVAL_105(coupler_from_tile_with_no_name__EVAL_105),
    ._EVAL_106(coupler_from_tile_with_no_name__EVAL_106),
    ._EVAL_107(coupler_from_tile_with_no_name__EVAL_107),
    ._EVAL_108(coupler_from_tile_with_no_name__EVAL_108)
  );
  _EVAL_19 coupler_to_sys_sram_1 (
    ._EVAL(coupler_to_sys_sram_1__EVAL),
    ._EVAL_0(coupler_to_sys_sram_1__EVAL_0),
    ._EVAL_1(coupler_to_sys_sram_1__EVAL_1),
    ._EVAL_2(coupler_to_sys_sram_1__EVAL_2),
    ._EVAL_3(coupler_to_sys_sram_1__EVAL_3),
    ._EVAL_4(coupler_to_sys_sram_1__EVAL_4),
    ._EVAL_5(coupler_to_sys_sram_1__EVAL_5),
    ._EVAL_6(coupler_to_sys_sram_1__EVAL_6),
    ._EVAL_7(coupler_to_sys_sram_1__EVAL_7),
    ._EVAL_8(coupler_to_sys_sram_1__EVAL_8),
    ._EVAL_9(coupler_to_sys_sram_1__EVAL_9),
    ._EVAL_10(coupler_to_sys_sram_1__EVAL_10),
    ._EVAL_11(coupler_to_sys_sram_1__EVAL_11),
    ._EVAL_12(coupler_to_sys_sram_1__EVAL_12),
    ._EVAL_13(coupler_to_sys_sram_1__EVAL_13),
    ._EVAL_14(coupler_to_sys_sram_1__EVAL_14),
    ._EVAL_15(coupler_to_sys_sram_1__EVAL_15),
    ._EVAL_16(coupler_to_sys_sram_1__EVAL_16),
    ._EVAL_17(coupler_to_sys_sram_1__EVAL_17),
    ._EVAL_18(coupler_to_sys_sram_1__EVAL_18),
    ._EVAL_19(coupler_to_sys_sram_1__EVAL_19),
    ._EVAL_20(coupler_to_sys_sram_1__EVAL_20),
    ._EVAL_21(coupler_to_sys_sram_1__EVAL_21),
    ._EVAL_22(coupler_to_sys_sram_1__EVAL_22),
    ._EVAL_23(coupler_to_sys_sram_1__EVAL_23),
    ._EVAL_24(coupler_to_sys_sram_1__EVAL_24),
    ._EVAL_25(coupler_to_sys_sram_1__EVAL_25),
    ._EVAL_26(coupler_to_sys_sram_1__EVAL_26),
    ._EVAL_27(coupler_to_sys_sram_1__EVAL_27),
    ._EVAL_28(coupler_to_sys_sram_1__EVAL_28),
    ._EVAL_29(coupler_to_sys_sram_1__EVAL_29),
    ._EVAL_30(coupler_to_sys_sram_1__EVAL_30),
    ._EVAL_31(coupler_to_sys_sram_1__EVAL_31),
    ._EVAL_32(coupler_to_sys_sram_1__EVAL_32)
  );
  _EVAL system_bus_clock_groups (
    ._EVAL_1(system_bus_clock_groups__EVAL_1),
    ._EVAL_2(system_bus_clock_groups__EVAL_2),
    ._EVAL_3(system_bus_clock_groups__EVAL_3),
    ._EVAL_4(system_bus_clock_groups__EVAL_4),
    ._EVAL_7(system_bus_clock_groups__EVAL_7),
    ._EVAL_10(system_bus_clock_groups__EVAL_10),
    ._EVAL_11(system_bus_clock_groups__EVAL_11),
    ._EVAL_12(system_bus_clock_groups__EVAL_12),
    ._EVAL_15(system_bus_clock_groups__EVAL_15),
    ._EVAL_17(system_bus_clock_groups__EVAL_17),
    ._EVAL_19(system_bus_clock_groups__EVAL_19),
    ._EVAL_22(system_bus_clock_groups__EVAL_22)
  );
  _EVAL_30 coupler_to_port_named_ahb_sys_port (
    ._EVAL(coupler_to_port_named_ahb_sys_port__EVAL),
    ._EVAL_0(coupler_to_port_named_ahb_sys_port__EVAL_0),
    ._EVAL_1(coupler_to_port_named_ahb_sys_port__EVAL_1),
    ._EVAL_2(coupler_to_port_named_ahb_sys_port__EVAL_2),
    ._EVAL_3(coupler_to_port_named_ahb_sys_port__EVAL_3),
    ._EVAL_4(coupler_to_port_named_ahb_sys_port__EVAL_4),
    ._EVAL_5(coupler_to_port_named_ahb_sys_port__EVAL_5),
    ._EVAL_6(coupler_to_port_named_ahb_sys_port__EVAL_6),
    ._EVAL_7(coupler_to_port_named_ahb_sys_port__EVAL_7),
    ._EVAL_8(coupler_to_port_named_ahb_sys_port__EVAL_8),
    ._EVAL_9(coupler_to_port_named_ahb_sys_port__EVAL_9),
    ._EVAL_10(coupler_to_port_named_ahb_sys_port__EVAL_10),
    ._EVAL_11(coupler_to_port_named_ahb_sys_port__EVAL_11),
    ._EVAL_12(coupler_to_port_named_ahb_sys_port__EVAL_12),
    ._EVAL_13(coupler_to_port_named_ahb_sys_port__EVAL_13),
    ._EVAL_14(coupler_to_port_named_ahb_sys_port__EVAL_14),
    ._EVAL_15(coupler_to_port_named_ahb_sys_port__EVAL_15),
    ._EVAL_16(coupler_to_port_named_ahb_sys_port__EVAL_16),
    ._EVAL_17(coupler_to_port_named_ahb_sys_port__EVAL_17),
    ._EVAL_18(coupler_to_port_named_ahb_sys_port__EVAL_18),
    ._EVAL_19(coupler_to_port_named_ahb_sys_port__EVAL_19),
    ._EVAL_20(coupler_to_port_named_ahb_sys_port__EVAL_20),
    ._EVAL_21(coupler_to_port_named_ahb_sys_port__EVAL_21),
    ._EVAL_22(coupler_to_port_named_ahb_sys_port__EVAL_22),
    ._EVAL_23(coupler_to_port_named_ahb_sys_port__EVAL_23),
    ._EVAL_24(coupler_to_port_named_ahb_sys_port__EVAL_24),
    ._EVAL_25(coupler_to_port_named_ahb_sys_port__EVAL_25),
    ._EVAL_26(coupler_to_port_named_ahb_sys_port__EVAL_26),
    ._EVAL_27(coupler_to_port_named_ahb_sys_port__EVAL_27),
    ._EVAL_28(coupler_to_port_named_ahb_sys_port__EVAL_28),
    ._EVAL_29(coupler_to_port_named_ahb_sys_port__EVAL_29),
    ._EVAL_30(coupler_to_port_named_ahb_sys_port__EVAL_30),
    ._EVAL_31(coupler_to_port_named_ahb_sys_port__EVAL_31),
    ._EVAL_32(coupler_to_port_named_ahb_sys_port__EVAL_32),
    ._EVAL_33(coupler_to_port_named_ahb_sys_port__EVAL_33),
    ._EVAL_34(coupler_to_port_named_ahb_sys_port__EVAL_34)
  );
  _EVAL_14 coupler_to_sys_sram_0 (
    ._EVAL(coupler_to_sys_sram_0__EVAL),
    ._EVAL_0(coupler_to_sys_sram_0__EVAL_0),
    ._EVAL_1(coupler_to_sys_sram_0__EVAL_1),
    ._EVAL_2(coupler_to_sys_sram_0__EVAL_2),
    ._EVAL_3(coupler_to_sys_sram_0__EVAL_3),
    ._EVAL_4(coupler_to_sys_sram_0__EVAL_4),
    ._EVAL_5(coupler_to_sys_sram_0__EVAL_5),
    ._EVAL_6(coupler_to_sys_sram_0__EVAL_6),
    ._EVAL_7(coupler_to_sys_sram_0__EVAL_7),
    ._EVAL_8(coupler_to_sys_sram_0__EVAL_8),
    ._EVAL_9(coupler_to_sys_sram_0__EVAL_9),
    ._EVAL_10(coupler_to_sys_sram_0__EVAL_10),
    ._EVAL_11(coupler_to_sys_sram_0__EVAL_11),
    ._EVAL_12(coupler_to_sys_sram_0__EVAL_12),
    ._EVAL_13(coupler_to_sys_sram_0__EVAL_13),
    ._EVAL_14(coupler_to_sys_sram_0__EVAL_14),
    ._EVAL_15(coupler_to_sys_sram_0__EVAL_15),
    ._EVAL_16(coupler_to_sys_sram_0__EVAL_16),
    ._EVAL_17(coupler_to_sys_sram_0__EVAL_17),
    ._EVAL_18(coupler_to_sys_sram_0__EVAL_18),
    ._EVAL_19(coupler_to_sys_sram_0__EVAL_19),
    ._EVAL_20(coupler_to_sys_sram_0__EVAL_20),
    ._EVAL_21(coupler_to_sys_sram_0__EVAL_21),
    ._EVAL_22(coupler_to_sys_sram_0__EVAL_22),
    ._EVAL_23(coupler_to_sys_sram_0__EVAL_23),
    ._EVAL_24(coupler_to_sys_sram_0__EVAL_24),
    ._EVAL_25(coupler_to_sys_sram_0__EVAL_25),
    ._EVAL_26(coupler_to_sys_sram_0__EVAL_26),
    ._EVAL_27(coupler_to_sys_sram_0__EVAL_27),
    ._EVAL_28(coupler_to_sys_sram_0__EVAL_28),
    ._EVAL_29(coupler_to_sys_sram_0__EVAL_29),
    ._EVAL_30(coupler_to_sys_sram_0__EVAL_30),
    ._EVAL_31(coupler_to_sys_sram_0__EVAL_31),
    ._EVAL_32(coupler_to_sys_sram_0__EVAL_32)
  );
  _EVAL_0 clockGroup (
    ._EVAL(clockGroup__EVAL),
    ._EVAL_0(clockGroup__EVAL_0),
    ._EVAL_1(clockGroup__EVAL_1),
    ._EVAL_2(clockGroup__EVAL_2)
  );
  assign _EVAL_13 = coupler_to_sys_sram_1__EVAL_6;
  assign coupler_to_port_named_ahb_sys_port__EVAL_0 = _EVAL_161;
  assign system_bus_xbar__EVAL_154 = fixedClockNode__EVAL_0;
  assign coupler_to_bus_named_cbus__EVAL_42 = system_bus_xbar__EVAL_130;
  assign fixedClockNode__EVAL = clockGroup__EVAL_1;
  assign _EVAL_167 = coupler_from_tile_with_no_name__EVAL_26;
  assign coupler_to_sys_sram_0__EVAL_7 = _EVAL_94;
  assign _EVAL_70 = coupler_to_sys_sram_0__EVAL_18;
  assign coupler_from_bus_named_front_bus__EVAL_14 = _EVAL_91;
  assign coupler_to_sys_sram_0__EVAL_32 = system_bus_xbar__EVAL_77;
  assign coupler_to_sys_sram_0__EVAL_9 = system_bus_xbar__EVAL_32;
  assign coupler_from_tile_with_no_name__EVAL_84 = _EVAL_117;
  assign _EVAL_81 = coupler_to_bus_named_cbus__EVAL_24;
  assign system_bus_xbar__EVAL_71 = coupler_from_tile_with_no_name__EVAL_24;
  assign _EVAL_26 = coupler_from_tile_with_no_name__EVAL_1;
  assign coupler_to_bus_named_cbus__EVAL_38 = system_bus_xbar__EVAL_43;
  assign coupler_from_tile_with_no_name__EVAL_52 = system_bus_xbar__EVAL_63;
  assign coupler_to_sys_sram_0__EVAL_28 = system_bus_xbar__EVAL_118;
  assign coupler_to_bus_named_cbus__EVAL_53 = system_bus_xbar__EVAL_26;
  assign _EVAL_1 = coupler_to_port_named_ahb_sys_port__EVAL_20;
  assign coupler_from_tile_with_no_name__EVAL_46 = _EVAL_59;
  assign _EVAL_164 = coupler_to_bus_named_cbus__EVAL_51;
  assign system_bus_xbar__EVAL_143 = coupler_to_bus_named_cbus__EVAL_0;
  assign _EVAL_119 = coupler_to_sys_sram_1__EVAL_16;
  assign system_bus_xbar__EVAL_58 = coupler_from_tile_with_no_name__EVAL_89;
  assign system_bus_xbar__EVAL_119 = coupler_from_bus_named_front_bus__EVAL_47;
  assign coupler_from_tile_with_no_name__EVAL_3 = system_bus_xbar__EVAL_105;
  assign coupler_to_bus_named_cbus__EVAL_16 = system_bus_xbar__EVAL_137;
  assign system_bus_xbar__EVAL_83 = coupler_from_tile_with_no_name__EVAL_88;
  assign _EVAL_60 = coupler_to_sys_sram_0__EVAL_0;
  assign coupler_from_tile_with_no_name__EVAL_87 = _EVAL_46;
  assign system_bus_xbar__EVAL_150 = coupler_from_tile_with_no_name__EVAL_69;
  assign _EVAL_160 = coupler_to_bus_named_cbus__EVAL_52;
  assign _EVAL_140 = coupler_from_bus_named_front_bus__EVAL_34;
  assign coupler_from_bus_named_front_bus__EVAL_42 = system_bus_xbar__EVAL_126;
  assign coupler_to_port_named_ahb_sys_port__EVAL_16 = system_bus_xbar__EVAL_88;
  assign _EVAL_58 = coupler_from_bus_named_front_bus__EVAL_4;
  assign coupler_from_tile_with_no_name__EVAL_96 = _EVAL_92;
  assign _EVAL_105 = coupler_to_bus_named_cbus__EVAL_4;
  assign coupler_from_tile_with_no_name__EVAL_25 = _EVAL_82;
  assign coupler_from_tile_with_no_name__EVAL_103 = _EVAL_170;
  assign coupler_to_port_named_ahb_sys_port__EVAL_12 = system_bus_xbar__EVAL_54;
  assign _EVAL_23 = coupler_to_sys_sram_1__EVAL_26;
  assign coupler_from_tile_with_no_name__EVAL_56 = system_bus_xbar__EVAL_24;
  assign _EVAL_154 = coupler_to_sys_sram_0__EVAL_3;
  assign coupler_to_port_named_ahb_sys_port__EVAL_15 = _EVAL_97;
  assign system_bus_xbar__EVAL_101 = coupler_to_port_named_ahb_sys_port__EVAL_33;
  assign coupler_from_tile_with_no_name__EVAL_70 = system_bus_xbar__EVAL_4;
  assign _EVAL_76 = coupler_to_port_named_ahb_sys_port__EVAL_8;
  assign _EVAL_130 = coupler_to_bus_named_cbus__EVAL_11;
  assign system_bus_xbar__EVAL_86 = coupler_from_tile_with_no_name__EVAL_100;
  assign coupler_to_port_named_ahb_sys_port__EVAL_34 = system_bus_xbar__EVAL_65;
  assign _EVAL_80 = coupler_to_bus_named_cbus__EVAL_8;
  assign coupler_from_tile_with_no_name__EVAL_83 = _EVAL_171;
  assign coupler_from_tile_with_no_name__EVAL_104 = system_bus_xbar__EVAL_39;
  assign coupler_from_bus_named_front_bus__EVAL_39 = _EVAL_85;
  assign coupler_from_tile_with_no_name__EVAL_105 = system_bus_xbar__EVAL_159;
  assign coupler_to_sys_sram_0__EVAL_14 = _EVAL_10;
  assign coupler_from_bus_named_front_bus__EVAL_6 = system_bus_xbar__EVAL_158;
  assign system_bus_xbar__EVAL_104 = coupler_from_tile_with_no_name__EVAL_39;
  assign coupler_to_sys_sram_1__EVAL_15 = system_bus_xbar__EVAL_29;
  assign coupler_from_tile_with_no_name__EVAL_13 = _EVAL_93;
  assign coupler_from_tile_with_no_name__EVAL_8 = _EVAL_169;
  assign coupler_to_bus_named_cbus__EVAL_2 = _EVAL_78;
  assign system_bus_xbar__EVAL_85 = coupler_from_bus_named_front_bus__EVAL_10;
  assign coupler_to_bus_named_cbus__EVAL_47 = system_bus_xbar__EVAL_31;
  assign _EVAL_20 = coupler_to_bus_named_cbus__EVAL_31;
  assign _EVAL_90 = coupler_to_sys_sram_0__EVAL_17;
  assign system_bus_xbar__EVAL_135 = coupler_from_tile_with_no_name__EVAL_99;
  assign system_bus_xbar__EVAL_28 = coupler_from_tile_with_no_name__EVAL_35;
  assign system_bus_xbar__EVAL_7 = coupler_from_tile_with_no_name__EVAL_58;
  assign system_bus_xbar__EVAL_37 = coupler_to_sys_sram_1__EVAL_4;
  assign coupler_to_port_named_ahb_sys_port__EVAL_18 = system_bus_xbar__EVAL_57;
  assign _EVAL_148 = coupler_from_tile_with_no_name__EVAL_41;
  assign coupler_from_bus_named_front_bus__EVAL_28 = _EVAL_101;
  assign coupler_to_sys_sram_1__EVAL = system_bus_xbar__EVAL_142;
  assign coupler_to_bus_named_cbus__EVAL_43 = _EVAL_68;
  assign system_bus_xbar__EVAL_14 = coupler_from_tile_with_no_name__EVAL_31;
  assign coupler_to_bus_named_cbus__EVAL_19 = _EVAL_44;
  assign _EVAL_34 = fixedClockNode__EVAL_2;
  assign system_bus_xbar__EVAL_133 = coupler_from_tile_with_no_name__EVAL_73;
  assign _EVAL_168 = coupler_to_bus_named_cbus__EVAL_50;
  assign coupler_to_sys_sram_1__EVAL_8 = system_bus_xbar__EVAL_100;
  assign coupler_to_bus_named_cbus__EVAL_15 = system_bus_xbar__EVAL_49;
  assign system_bus_xbar__EVAL_162 = fixedClockNode__EVAL_2;
  assign _EVAL_123 = coupler_to_port_named_ahb_sys_port__EVAL_27;
  assign system_bus_xbar__EVAL_121 = coupler_to_port_named_ahb_sys_port__EVAL_5;
  assign _EVAL_136 = coupler_from_tile_with_no_name__EVAL_2;
  assign _EVAL_54 = coupler_from_tile_with_no_name__EVAL_63;
  assign coupler_from_tile_with_no_name__EVAL_86 = _EVAL_77;
  assign system_bus_xbar__EVAL_138 = coupler_from_bus_named_front_bus__EVAL_45;
  assign _EVAL_62 = system_bus_clock_groups__EVAL_4;
  assign coupler_from_bus_named_front_bus__EVAL_32 = system_bus_xbar__EVAL_147;
  assign coupler_to_sys_sram_0__EVAL_16 = system_bus_xbar__EVAL_2;
  assign system_bus_xbar__EVAL_108 = coupler_from_bus_named_front_bus__EVAL_49;
  assign system_bus_xbar__EVAL_34 = coupler_to_port_named_ahb_sys_port__EVAL_32;
  assign _EVAL_99 = coupler_to_bus_named_cbus__EVAL_22;
  assign coupler_from_tile_with_no_name__EVAL_38 = _EVAL_134;
  assign coupler_from_tile_with_no_name__EVAL_75 = _EVAL_125;
  assign coupler_from_tile_with_no_name__EVAL_67 = system_bus_xbar__EVAL_106;
  assign system_bus_xbar__EVAL_61 = coupler_from_bus_named_front_bus__EVAL_44;
  assign coupler_to_sys_sram_1__EVAL_21 = _EVAL_45;
  assign _EVAL_29 = coupler_to_sys_sram_0__EVAL_24;
  assign coupler_to_bus_named_cbus__EVAL_41 = fixedClockNode__EVAL_2;
  assign coupler_from_tile_with_no_name__EVAL_108 = _EVAL_152;
  assign coupler_from_bus_named_front_bus__EVAL_13 = _EVAL_129;
  assign system_bus_xbar__EVAL_91 = coupler_from_bus_named_front_bus__EVAL_48;
  assign _EVAL_52 = coupler_to_bus_named_cbus__EVAL_9;
  assign _EVAL_14 = coupler_from_tile_with_no_name__EVAL_20;
  assign coupler_from_tile_with_no_name__EVAL_71 = system_bus_xbar__EVAL_38;
  assign system_bus_xbar__EVAL_112 = coupler_to_bus_named_cbus__EVAL_39;
  assign _EVAL_67 = coupler_from_tile_with_no_name__EVAL_61;
  assign coupler_to_sys_sram_1__EVAL_3 = system_bus_xbar__EVAL_146;
  assign coupler_to_sys_sram_1__EVAL_32 = system_bus_xbar__EVAL_27;
  assign coupler_to_sys_sram_0__EVAL_12 = system_bus_xbar__EVAL_41;
  assign coupler_to_port_named_ahb_sys_port__EVAL = system_bus_xbar__EVAL_84;
  assign _EVAL_17 = fixedClockNode__EVAL_0;
  assign coupler_to_bus_named_cbus__EVAL_48 = system_bus_xbar__EVAL_3;
  assign system_bus_clock_groups__EVAL_17 = _EVAL_63;
  assign coupler_from_tile_with_no_name__EVAL_29 = system_bus_xbar__EVAL_17;
  assign _EVAL_7 = coupler_from_tile_with_no_name__EVAL_19;
  assign coupler_to_sys_sram_1__EVAL_24 = fixedClockNode__EVAL_2;
  assign system_bus_xbar__EVAL_117 = coupler_to_bus_named_cbus__EVAL_7;
  assign coupler_to_bus_named_cbus__EVAL_54 = _EVAL_41;
  assign system_bus_xbar__EVAL_120 = coupler_from_tile_with_no_name__EVAL_36;
  assign system_bus_xbar__EVAL_93 = coupler_to_bus_named_cbus__EVAL_40;
  assign system_bus_xbar__EVAL_141 = coupler_from_bus_named_front_bus__EVAL_21;
  assign coupler_from_bus_named_front_bus__EVAL = system_bus_xbar__EVAL_157;
  assign coupler_from_tile_with_no_name__EVAL_50 = system_bus_xbar__EVAL_60;
  assign system_bus_xbar__EVAL_125 = coupler_from_bus_named_front_bus__EVAL_38;
  assign clockGroup__EVAL = system_bus_clock_groups__EVAL_7;
  assign coupler_to_sys_sram_0__EVAL_1 = _EVAL_56;
  assign system_bus_xbar__EVAL_52 = coupler_from_tile_with_no_name__EVAL_101;
  assign _EVAL_120 = system_bus_clock_groups__EVAL_22;
  assign coupler_to_sys_sram_0__EVAL_21 = _EVAL_74;
  assign system_bus_xbar__EVAL_94 = coupler_from_tile_with_no_name__EVAL_6;
  assign _EVAL_21 = coupler_to_bus_named_cbus__EVAL_14;
  assign system_bus_xbar__EVAL_149 = coupler_from_tile_with_no_name__EVAL_55;
  assign coupler_from_tile_with_no_name__EVAL_33 = _EVAL_139;
  assign system_bus_xbar__EVAL_132 = coupler_to_sys_sram_0__EVAL_6;
  assign system_bus_xbar__EVAL_160 = coupler_to_port_named_ahb_sys_port__EVAL_23;
  assign coupler_to_sys_sram_1__EVAL_20 = _EVAL_141;
  assign coupler_from_tile_with_no_name__EVAL_81 = system_bus_xbar__EVAL_18;
  assign system_bus_xbar__EVAL_96 = coupler_to_sys_sram_1__EVAL_1;
  assign coupler_from_tile_with_no_name__EVAL_95 = _EVAL_114;
  assign coupler_to_bus_named_cbus__EVAL_5 = system_bus_xbar__EVAL_51;
  assign coupler_to_bus_named_cbus__EVAL_30 = system_bus_xbar__EVAL_5;
  assign coupler_to_sys_sram_0__EVAL_10 = system_bus_xbar__EVAL_80;
  assign _EVAL_30 = coupler_to_sys_sram_1__EVAL_2;
  assign _EVAL_132 = coupler_from_bus_named_front_bus__EVAL_41;
  assign coupler_from_bus_named_front_bus__EVAL_18 = _EVAL_95;
  assign coupler_from_tile_with_no_name__EVAL_62 = fixedClockNode__EVAL_0;
  assign system_bus_xbar__EVAL_139 = coupler_from_bus_named_front_bus__EVAL_51;
  assign system_bus_xbar__EVAL_87 = coupler_from_bus_named_front_bus__EVAL_52;
  assign coupler_to_sys_sram_0__EVAL_29 = system_bus_xbar__EVAL_70;
  assign coupler_to_port_named_ahb_sys_port__EVAL_25 = system_bus_xbar__EVAL_78;
  assign coupler_from_bus_named_front_bus__EVAL_26 = system_bus_xbar__EVAL_129;
  assign system_bus_xbar__EVAL_97 = coupler_from_bus_named_front_bus__EVAL_12;
  assign _EVAL_2 = coupler_from_bus_named_front_bus__EVAL_8;
  assign system_bus_xbar__EVAL_89 = coupler_from_bus_named_front_bus__EVAL_19;
  assign _EVAL_142 = coupler_to_bus_named_cbus__EVAL_32;
  assign coupler_from_tile_with_no_name__EVAL_76 = system_bus_xbar__EVAL_67;
  assign coupler_to_sys_sram_0__EVAL_31 = system_bus_xbar__EVAL_102;
  assign _EVAL_37 = coupler_from_tile_with_no_name__EVAL_5;
  assign system_bus_xbar__EVAL_72 = coupler_to_sys_sram_1__EVAL_7;
  assign _EVAL_124 = coupler_to_port_named_ahb_sys_port__EVAL_26;
  assign coupler_from_tile_with_no_name__EVAL_65 = _EVAL_143;
  assign _EVAL = coupler_from_tile_with_no_name__EVAL_37;
  assign coupler_to_port_named_ahb_sys_port__EVAL_13 = system_bus_xbar__EVAL_144;
  assign coupler_from_bus_named_front_bus__EVAL_24 = _EVAL_9;
  assign coupler_from_tile_with_no_name__EVAL_23 = system_bus_xbar__EVAL_151;
  assign _EVAL_116 = coupler_to_sys_sram_1__EVAL_0;
  assign system_bus_xbar__EVAL_148 = coupler_to_sys_sram_0__EVAL_15;
  assign system_bus_xbar__EVAL_73 = coupler_from_tile_with_no_name__EVAL_21;
  assign system_bus_xbar__EVAL_8 = coupler_to_sys_sram_0__EVAL_22;
  assign coupler_to_sys_sram_1__EVAL_27 = system_bus_xbar__EVAL_103;
  assign coupler_from_tile_with_no_name__EVAL_77 = system_bus_xbar__EVAL_140;
  assign coupler_from_bus_named_front_bus__EVAL_2 = system_bus_xbar__EVAL_123;
  assign coupler_to_bus_named_cbus__EVAL_46 = system_bus_xbar__EVAL_107;
  assign coupler_to_sys_sram_1__EVAL_28 = _EVAL_25;
  assign coupler_to_sys_sram_0__EVAL_11 = _EVAL_33;
  assign _EVAL_135 = coupler_to_bus_named_cbus__EVAL_36;
  assign _EVAL_162 = coupler_to_port_named_ahb_sys_port__EVAL_14;
  assign coupler_from_tile_with_no_name__EVAL_98 = fixedClockNode__EVAL_2;
  assign coupler_to_port_named_ahb_sys_port__EVAL_31 = system_bus_xbar__EVAL_53;
  assign coupler_from_tile_with_no_name__EVAL_90 = system_bus_xbar__EVAL_64;
  assign coupler_from_tile_with_no_name__EVAL_53 = _EVAL_43;
  assign coupler_from_bus_named_front_bus__EVAL_15 = fixedClockNode__EVAL_0;
  assign _EVAL_138 = coupler_from_tile_with_no_name__EVAL_48;
  assign coupler_to_bus_named_cbus__EVAL_3 = _EVAL_73;
  assign coupler_to_bus_named_cbus__EVAL_6 = system_bus_xbar__EVAL_66;
  assign coupler_to_port_named_ahb_sys_port__EVAL_6 = system_bus_xbar__EVAL_44;
  assign coupler_to_sys_sram_1__EVAL_12 = fixedClockNode__EVAL_0;
  assign coupler_to_bus_named_cbus__EVAL_49 = system_bus_xbar__EVAL_92;
  assign coupler_from_tile_with_no_name__EVAL_107 = _EVAL_4;
  assign coupler_from_tile_with_no_name__EVAL_64 = _EVAL_71;
  assign _EVAL_61 = coupler_from_tile_with_no_name__EVAL_54;
  assign system_bus_xbar__EVAL_45 = coupler_from_tile_with_no_name__EVAL_10;
  assign coupler_from_tile_with_no_name__EVAL_106 = _EVAL_107;
  assign coupler_from_tile_with_no_name__EVAL_22 = _EVAL_38;
  assign system_bus_xbar__EVAL_113 = coupler_from_bus_named_front_bus__EVAL_11;
  assign coupler_from_tile_with_no_name__EVAL_47 = _EVAL_53;
  assign _EVAL_50 = system_bus_clock_groups__EVAL_11;
  assign _EVAL_150 = coupler_to_sys_sram_1__EVAL_18;
  assign _EVAL_147 = coupler_to_sys_sram_0__EVAL;
  assign coupler_to_sys_sram_1__EVAL_29 = _EVAL_108;
  assign system_bus_xbar__EVAL_12 = coupler_from_tile_with_no_name__EVAL_49;
  assign _EVAL_122 = coupler_from_bus_named_front_bus__EVAL_43;
  assign _EVAL_100 = coupler_from_tile_with_no_name__EVAL_59;
  assign coupler_from_bus_named_front_bus__EVAL_20 = _EVAL_137;
  assign coupler_to_bus_named_cbus__EVAL_18 = _EVAL_72;
  assign system_bus_xbar__EVAL_25 = coupler_to_sys_sram_0__EVAL_23;
  assign coupler_from_tile_with_no_name__EVAL_102 = _EVAL_98;
  assign coupler_from_tile_with_no_name__EVAL_72 = system_bus_xbar__EVAL_145;
  assign coupler_from_tile_with_no_name__EVAL_44 = system_bus_xbar__EVAL_62;
  assign system_bus_xbar__EVAL_74 = coupler_to_bus_named_cbus__EVAL_29;
  assign coupler_to_bus_named_cbus__EVAL = _EVAL_39;
  assign system_bus_xbar__EVAL_110 = coupler_from_tile_with_no_name__EVAL_97;
  assign system_bus_xbar__EVAL_50 = coupler_from_bus_named_front_bus__EVAL_27;
  assign system_bus_xbar__EVAL_20 = coupler_from_tile_with_no_name__EVAL_14;
  assign system_bus_xbar__EVAL_48 = coupler_from_tile_with_no_name__EVAL;
  assign coupler_to_port_named_ahb_sys_port__EVAL_3 = system_bus_xbar__EVAL_153;
  assign system_bus_clock_groups__EVAL_2 = _EVAL_84;
  assign system_bus_xbar__EVAL_75 = coupler_from_bus_named_front_bus__EVAL_29;
  assign system_bus_xbar__EVAL_55 = coupler_from_tile_with_no_name__EVAL_92;
  assign coupler_from_bus_named_front_bus__EVAL_22 = _EVAL_64;
  assign system_bus_xbar__EVAL_59 = coupler_to_port_named_ahb_sys_port__EVAL_4;
  assign _EVAL_144 = coupler_to_sys_sram_0__EVAL_27;
  assign coupler_to_sys_sram_0__EVAL_20 = _EVAL_110;
  assign system_bus_xbar__EVAL_163 = coupler_from_bus_named_front_bus__EVAL_23;
  assign _EVAL_96 = coupler_from_tile_with_no_name__EVAL_78;
  assign coupler_to_bus_named_cbus__EVAL_34 = system_bus_xbar__EVAL_76;
  assign system_bus_xbar__EVAL_136 = coupler_from_tile_with_no_name__EVAL_4;
  assign coupler_from_bus_named_front_bus__EVAL_5 = system_bus_xbar__EVAL_127;
  assign fixedClockNode__EVAL_1 = clockGroup__EVAL_0;
  assign _EVAL_131 = coupler_from_bus_named_front_bus__EVAL_25;
  assign coupler_from_tile_with_no_name__EVAL_66 = system_bus_xbar__EVAL_156;
  assign _EVAL_118 = coupler_to_sys_sram_0__EVAL_8;
  assign coupler_from_tile_with_no_name__EVAL_79 = _EVAL_6;
  assign system_bus_xbar__EVAL = coupler_to_sys_sram_0__EVAL_4;
  assign system_bus_xbar__EVAL_6 = coupler_to_bus_named_cbus__EVAL_1;
  assign system_bus_xbar__EVAL_47 = coupler_to_port_named_ahb_sys_port__EVAL_7;
  assign system_bus_xbar__EVAL_36 = coupler_to_bus_named_cbus__EVAL_17;
  assign clockGroup__EVAL_2 = system_bus_clock_groups__EVAL_3;
  assign coupler_from_bus_named_front_bus__EVAL_0 = system_bus_xbar__EVAL_19;
  assign system_bus_xbar__EVAL_30 = coupler_to_sys_sram_1__EVAL_9;
  assign coupler_to_sys_sram_0__EVAL_26 = system_bus_xbar__EVAL_116;
  assign system_bus_xbar__EVAL_155 = coupler_from_tile_with_no_name__EVAL_45;
  assign coupler_to_sys_sram_1__EVAL_23 = system_bus_xbar__EVAL_81;
  assign system_bus_xbar__EVAL_128 = coupler_from_tile_with_no_name__EVAL_11;
  assign coupler_to_port_named_ahb_sys_port__EVAL_11 = fixedClockNode__EVAL_0;
  assign system_bus_xbar__EVAL_90 = coupler_from_bus_named_front_bus__EVAL_9;
  assign coupler_from_tile_with_no_name__EVAL_82 = _EVAL_103;
  assign system_bus_xbar__EVAL_69 = coupler_from_tile_with_no_name__EVAL_85;
  assign _EVAL_18 = coupler_from_tile_with_no_name__EVAL_51;
  assign system_bus_xbar__EVAL_1 = coupler_from_tile_with_no_name__EVAL_40;
  assign _EVAL_27 = coupler_to_sys_sram_1__EVAL_17;
  assign coupler_to_port_named_ahb_sys_port__EVAL_29 = _EVAL_51;
  assign _EVAL_66 = coupler_to_port_named_ahb_sys_port__EVAL_2;
  assign coupler_to_port_named_ahb_sys_port__EVAL_9 = system_bus_xbar__EVAL_10;
  assign _EVAL_69 = coupler_from_tile_with_no_name__EVAL_94;
  assign coupler_to_bus_named_cbus__EVAL_26 = system_bus_xbar__EVAL_21;
  assign coupler_from_bus_named_front_bus__EVAL_40 = system_bus_xbar__EVAL_131;
  assign system_bus_xbar__EVAL_95 = coupler_to_sys_sram_1__EVAL_25;
  assign coupler_from_bus_named_front_bus__EVAL_35 = _EVAL_0;
  assign coupler_from_bus_named_front_bus__EVAL_36 = _EVAL_112;
  assign coupler_from_tile_with_no_name__EVAL_18 = _EVAL_111;
  assign coupler_from_tile_with_no_name__EVAL_60 = _EVAL_104;
  assign coupler_to_bus_named_cbus__EVAL_21 = system_bus_xbar__EVAL_99;
  assign system_bus_xbar__EVAL_0 = coupler_from_tile_with_no_name__EVAL_7;
  assign coupler_to_bus_named_cbus__EVAL_33 = _EVAL_36;
  assign coupler_from_bus_named_front_bus__EVAL_33 = _EVAL_42;
  assign system_bus_xbar__EVAL_40 = coupler_to_port_named_ahb_sys_port__EVAL_17;
  assign _EVAL_15 = coupler_from_tile_with_no_name__EVAL_74;
  assign system_bus_xbar__EVAL_122 = coupler_from_tile_with_no_name__EVAL_42;
  assign system_bus_xbar__EVAL_124 = coupler_to_port_named_ahb_sys_port__EVAL_19;
  assign _EVAL_89 = coupler_to_sys_sram_0__EVAL_25;
  assign coupler_to_sys_sram_0__EVAL_13 = fixedClockNode__EVAL_2;
  assign system_bus_xbar__EVAL_79 = coupler_from_tile_with_no_name__EVAL_16;
  assign coupler_to_sys_sram_1__EVAL_13 = _EVAL_126;
  assign _EVAL_165 = coupler_to_sys_sram_1__EVAL_10;
  assign coupler_from_tile_with_no_name__EVAL_91 = _EVAL_102;
  assign system_bus_xbar__EVAL_33 = coupler_from_tile_with_no_name__EVAL_80;
  assign coupler_to_bus_named_cbus__EVAL_25 = fixedClockNode__EVAL_0;
  assign _EVAL_157 = coupler_to_sys_sram_1__EVAL_22;
  assign _EVAL_57 = coupler_to_sys_sram_0__EVAL_19;
  assign _EVAL_79 = coupler_to_port_named_ahb_sys_port__EVAL_10;
  assign system_bus_xbar__EVAL_22 = coupler_to_sys_sram_0__EVAL_30;
  assign system_bus_clock_groups__EVAL_12 = _EVAL_158;
  assign coupler_to_sys_sram_0__EVAL_2 = system_bus_xbar__EVAL_82;
  assign coupler_to_port_named_ahb_sys_port__EVAL_1 = system_bus_xbar__EVAL_56;
  assign _EVAL_12 = coupler_to_sys_sram_1__EVAL_19;
  assign _EVAL_47 = coupler_from_tile_with_no_name__EVAL_57;
  assign coupler_from_tile_with_no_name__EVAL_30 = _EVAL_106;
  assign system_bus_xbar__EVAL_152 = coupler_to_bus_named_cbus__EVAL_45;
  assign _EVAL_86 = coupler_from_tile_with_no_name__EVAL_28;
  assign _EVAL_28 = coupler_from_bus_named_front_bus__EVAL_3;
  assign coupler_from_tile_with_no_name__EVAL_15 = system_bus_xbar__EVAL_98;
  assign system_bus_xbar__EVAL_23 = coupler_to_bus_named_cbus__EVAL_23;
  assign _EVAL_156 = system_bus_clock_groups__EVAL_15;
  assign system_bus_xbar__EVAL_115 = coupler_from_tile_with_no_name__EVAL_93;
  assign _EVAL_3 = coupler_to_bus_named_cbus__EVAL_12;
  assign system_bus_xbar__EVAL_109 = coupler_to_bus_named_cbus__EVAL_13;
  assign coupler_from_tile_with_no_name__EVAL_32 = _EVAL_65;
  assign coupler_to_port_named_ahb_sys_port__EVAL_22 = fixedClockNode__EVAL_2;
  assign system_bus_clock_groups__EVAL_1 = _EVAL_153;
  assign coupler_from_tile_with_no_name__EVAL_43 = _EVAL_48;
  assign system_bus_xbar__EVAL_134 = coupler_to_port_named_ahb_sys_port__EVAL_24;
  assign _EVAL_16 = coupler_to_bus_named_cbus__EVAL_10;
  assign system_bus_clock_groups__EVAL_19 = _EVAL_55;
  assign coupler_from_bus_named_front_bus__EVAL_17 = _EVAL_8;
  assign coupler_from_tile_with_no_name__EVAL_17 = _EVAL_87;
  assign coupler_from_bus_named_front_bus__EVAL_7 = _EVAL_151;
  assign coupler_to_sys_sram_0__EVAL_5 = fixedClockNode__EVAL_0;
  assign coupler_to_sys_sram_1__EVAL_5 = system_bus_xbar__EVAL_16;
  assign _EVAL_5 = coupler_from_tile_with_no_name__EVAL_12;
  assign coupler_to_port_named_ahb_sys_port__EVAL_28 = system_bus_xbar__EVAL_68;
  assign system_bus_xbar__EVAL_46 = coupler_from_tile_with_no_name__EVAL_34;
  assign coupler_from_bus_named_front_bus__EVAL_50 = _EVAL_115;
  assign system_bus_clock_groups__EVAL_10 = _EVAL_133;
  assign coupler_to_sys_sram_1__EVAL_31 = _EVAL_109;
  assign _EVAL_24 = coupler_from_bus_named_front_bus__EVAL_31;
  assign system_bus_xbar__EVAL_15 = coupler_to_sys_sram_1__EVAL_11;
  assign coupler_from_tile_with_no_name__EVAL_68 = _EVAL_121;
  assign coupler_to_bus_named_cbus__EVAL_35 = _EVAL_146;
  assign coupler_from_bus_named_front_bus__EVAL_1 = _EVAL_31;
  assign coupler_to_bus_named_cbus__EVAL_44 = system_bus_xbar__EVAL_161;
  assign _EVAL_19 = coupler_to_bus_named_cbus__EVAL_28;
  assign coupler_to_sys_sram_1__EVAL_14 = system_bus_xbar__EVAL_114;
  assign coupler_to_bus_named_cbus__EVAL_27 = system_bus_xbar__EVAL_9;
  assign coupler_to_port_named_ahb_sys_port__EVAL_30 = system_bus_xbar__EVAL_42;
  assign coupler_from_bus_named_front_bus__EVAL_16 = _EVAL_11;
  assign _EVAL_128 = coupler_from_bus_named_front_bus__EVAL_46;
  assign system_bus_xbar__EVAL_13 = coupler_from_tile_with_no_name__EVAL_0;
  assign coupler_from_bus_named_front_bus__EVAL_30 = fixedClockNode__EVAL_2;
  assign coupler_to_bus_named_cbus__EVAL_37 = _EVAL_32;
  assign _EVAL_83 = coupler_to_bus_named_cbus__EVAL_20;
  assign system_bus_xbar__EVAL_111 = coupler_to_port_named_ahb_sys_port__EVAL_21;
  assign coupler_from_tile_with_no_name__EVAL_27 = system_bus_xbar__EVAL_11;
  assign coupler_from_tile_with_no_name__EVAL_9 = _EVAL_113;
  assign coupler_from_bus_named_front_bus__EVAL_37 = _EVAL_159;
  assign coupler_to_sys_sram_1__EVAL_30 = system_bus_xbar__EVAL_35;
endmodule
