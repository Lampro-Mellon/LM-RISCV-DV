//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_178_assert(
  input  [2:0]  _EVAL,
  input  [2:0]  _EVAL_0,
  input  [14:0] _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [3:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input  [1:0]  _EVAL_9,
  input  [1:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13
);
  wire  _EVAL_14;
  wire  _EVAL_15;
  wire [4:0] _EVAL_16;
  wire [1:0] _EVAL_17;
  wire [1:0] _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  reg [2:0] _EVAL_32;
  reg [31:0] _RAND_0;
  reg [4:0] _EVAL_33;
  reg [31:0] _RAND_1;
  wire [7:0] _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire [4:0] _EVAL_37;
  wire  _EVAL_38;
  reg [1:0] _EVAL_39;
  reg [31:0] _RAND_2;
  wire  _EVAL_40;
  wire [1:0] _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire [14:0] _EVAL_47;
  reg [31:0] _EVAL_48;
  reg [31:0] _RAND_3;
  wire  _EVAL_49;
  reg  _EVAL_51;
  reg [31:0] _RAND_4;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  reg [14:0] _EVAL_57;
  reg [31:0] _RAND_5;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire [1:0] _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire [7:0] _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  reg [2:0] _EVAL_73;
  reg [31:0] _RAND_6;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  reg [2:0] _EVAL_78;
  reg [31:0] _RAND_7;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire [15:0] _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  reg  _EVAL_91;
  reg [31:0] _RAND_8;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire [14:0] _EVAL_94;
  reg [2:0] _EVAL_95;
  reg [31:0] _RAND_9;
  reg  _EVAL_96;
  reg [31:0] _RAND_10;
  wire [4:0] _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire [1:0] _EVAL_103;
  wire  _EVAL_104;
  wire [4:0] _EVAL_105;
  wire [15:0] _EVAL_107;
  reg  _EVAL_108;
  reg [31:0] _RAND_11;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire [4:0] _EVAL_114;
  wire  _EVAL_115;
  wire [4:0] _EVAL_116;
  wire [7:0] _EVAL_117;
  wire [3:0] _EVAL_118;
  wire  _EVAL_119;
  wire [1:0] _EVAL_120;
  wire [14:0] _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire [15:0] _EVAL_130;
  wire  _EVAL_132;
  wire  _EVAL_133;
  reg [1:0] _EVAL_134;
  reg [31:0] _RAND_12;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [1:0] _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire [7:0] _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire [32:0] _EVAL_157;
  wire  _EVAL_158;
  reg [2:0] _EVAL_159;
  reg [31:0] _RAND_13;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire [31:0] _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire [3:0] _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire [3:0] _EVAL_189;
  wire [4:0] _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire [1:0] _EVAL_200;
  wire  _EVAL_201;
  wire [3:0] _EVAL_202;
  wire [4:0] _EVAL_203;
  wire  _EVAL_204;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_79 = _EVAL_48 < plusarg_reader_out;
  assign _EVAL_21 = _EVAL_6 & _EVAL_188;
  assign _EVAL_130 = _EVAL_107;
  assign _EVAL_64 = ~_EVAL_60;
  assign _EVAL_198 = _EVAL_33 != 5'h0;
  assign _EVAL_77 = ~_EVAL_158;
  assign _EVAL_157 = _EVAL_48 + 32'h1;
  assign _EVAL_127 = _EVAL_4 == _EVAL_202;
  assign _EVAL_194 = _EVAL <= 3'h3;
  assign _EVAL_173 = ~_EVAL_61;
  assign _EVAL_44 = _EVAL_3 == 3'h5;
  assign _EVAL_181 = _EVAL_3 == 3'h3;
  assign _EVAL_98 = ~_EVAL_12;
  assign _EVAL_61 = _EVAL_9 >= 2'h2;
  assign _EVAL_53 = ~_EVAL_132;
  assign _EVAL_58 = ~_EVAL_63;
  assign _EVAL_202 = {_EVAL_84,_EVAL_166,_EVAL_90,_EVAL_36};
  assign _EVAL_178 = ~_EVAL_4;
  assign _EVAL_195 = ~_EVAL_68;
  assign _EVAL_111 = ~_EVAL_102;
  assign _EVAL_18 = _EVAL_51 - 1'h1;
  assign _EVAL_104 = ~_EVAL_198;
  assign _EVAL_138 = _EVAL_7 == 3'h2;
  assign _EVAL_103 = _EVAL_108 - 1'h1;
  assign _EVAL_46 = _EVAL_7 == 3'h5;
  assign _EVAL_144 = ~_EVAL_91;
  assign _EVAL_26 = _EVAL_165 & _EVAL_170;
  assign _EVAL_68 = ~_EVAL_139;
  assign _EVAL_163 = ~_EVAL_196;
  assign _EVAL_93 = ~_EVAL_43;
  assign _EVAL_186 = _EVAL_6 & _EVAL_101;
  assign _EVAL_162 = ~_EVAL_65;
  assign _EVAL_158 = _EVAL_7 == _EVAL_78;
  assign _EVAL_150 = _EVAL_1[1];
  assign _EVAL_118 = ~_EVAL_202;
  assign _EVAL_199 = _EVAL_83 | _EVAL_67;
  assign _EVAL_151 = _EVAL_112 & _EVAL_122;
  assign _EVAL_189 = _EVAL_4 & _EVAL_118;
  assign _EVAL_72 = ~_EVAL_145;
  assign _EVAL_43 = _EVAL <= 3'h1;
  assign _EVAL_133 = ~_EVAL_185;
  assign _EVAL_14 = _EVAL_5 & _EVAL_177;
  assign _EVAL_121 = _EVAL_1 & _EVAL_94;
  assign _EVAL_120 = _EVAL_41 | 2'h1;
  assign _EVAL_67 = _EVAL_89 & _EVAL_112;
  assign _EVAL_143 = _EVAL_96 - 1'h1;
  assign _EVAL_193 = _EVAL_5 & _EVAL_88;
  assign _EVAL_49 = _EVAL_11 <= 3'h4;
  assign _EVAL_149 = _EVAL_119 | _EVAL_79;
  assign _EVAL_128 = ~_EVAL_31;
  assign _EVAL_140 = ~_EVAL_180;
  assign _EVAL_16 = _EVAL_117[4:0];
  assign _EVAL_179 = _EVAL_24 & _EVAL_147;
  assign _EVAL_154 = _EVAL_83 | _EVAL_148;
  assign _EVAL_161 = _EVAL_5 & _EVAL_135;
  assign _EVAL_152 = _EVAL_5 & _EVAL_141;
  assign _EVAL_126 = ~_EVAL_160;
  assign _EVAL_85 = _EVAL_6 & _EVAL_155;
  assign _EVAL_65 = _EVAL_11 == _EVAL_159;
  assign _EVAL_117 = _EVAL_182 ? _EVAL_70 : 8'h0;
  assign _EVAL_174 = _EVAL_112 & _EVAL_86;
  assign _EVAL_24 = _EVAL_10 <= 2'h2;
  assign _EVAL_54 = ~_EVAL_123;
  assign _EVAL_172 = ~_EVAL_204;
  assign _EVAL_183 = ~_EVAL_127;
  assign _EVAL_180 = _EVAL_7 == 3'h6;
  assign _EVAL_29 = ~_EVAL_187;
  assign _EVAL_132 = _EVAL_1 == _EVAL_57;
  assign _EVAL_30 = ~_EVAL_115;
  assign _EVAL_81 = _EVAL_3 == _EVAL_95;
  assign _EVAL_197 = ~_EVAL_98;
  assign _EVAL_155 = ~_EVAL_69;
  assign _EVAL_99 = _EVAL_6 & _EVAL_138;
  assign _EVAL_177 = _EVAL_3 == 3'h4;
  assign _EVAL_171 = _EVAL_5 & _EVAL_40;
  assign _EVAL_55 = ~_EVAL_81;
  assign _EVAL_76 = _EVAL_150 & _EVAL_122;
  assign _EVAL_203 = _EVAL_105 >> _EVAL_11;
  assign _EVAL_36 = _EVAL_199 | _EVAL_100;
  assign _EVAL_107 = $signed(_EVAL_87) & -16'sh1000;
  assign _EVAL_184 = _EVAL_192 & _EVAL_76;
  assign _EVAL_142 = _EVAL != 3'h0;
  assign _EVAL_42 = _EVAL_59 | _EVAL_165;
  assign _EVAL_17 = _EVAL_97[1:0];
  assign _EVAL_102 = _EVAL == _EVAL_73;
  assign _EVAL_28 = ~_EVAL_179;
  assign _EVAL_191 = _EVAL_165 & _EVAL_69;
  assign _EVAL_135 = _EVAL_3 == 3'h0;
  assign _EVAL_94 = {{13'd0}, _EVAL_66};
  assign _EVAL_204 = _EVAL_0 <= 3'h4;
  assign _EVAL_62 = _EVAL_5 & _EVAL_181;
  assign _EVAL_116 = ~_EVAL_16;
  assign _EVAL_31 = _EVAL_121 == 15'h0;
  assign _EVAL_90 = _EVAL_199 | _EVAL_109;
  assign _EVAL_92 = _EVAL_6 & _EVAL_46;
  assign _EVAL_100 = _EVAL_192 & _EVAL_174;
  assign _EVAL_63 = _EVAL_7 <= 3'h6;
  assign _EVAL_47 = _EVAL_1 ^ 15'h4000;
  assign _EVAL_182 = _EVAL_26 & _EVAL_140;
  assign _EVAL_113 = ~_EVAL_164;
  assign _EVAL_37 = _EVAL_33 >> _EVAL_0;
  assign _EVAL_109 = _EVAL_192 & _EVAL_151;
  assign _EVAL_22 = _EVAL_0 == _EVAL_32;
  assign _EVAL_25 = plusarg_reader_out == 32'h0;
  assign _EVAL_176 = _EVAL_103[0];
  assign _EVAL_123 = _EVAL_9 == _EVAL_39;
  assign _EVAL_122 = _EVAL_1[0];
  assign _EVAL_201 = _EVAL_203[0];
  assign _EVAL_112 = ~_EVAL_150;
  assign _EVAL_83 = _EVAL_10 >= 2'h2;
  assign _EVAL_147 = $signed(_EVAL_130) == 16'sh0;
  assign _EVAL_125 = _EVAL_200[0];
  assign _EVAL_196 = ~_EVAL_96;
  assign _EVAL_153 = ~_EVAL_49;
  assign _EVAL_175 = _EVAL_157[31:0];
  assign _EVAL_114 = _EVAL_34[4:0];
  assign _EVAL_148 = _EVAL_89 & _EVAL_150;
  assign _EVAL_187 = _EVAL <= 3'h2;
  assign _EVAL_38 = _EVAL_6 & _EVAL_23;
  assign _EVAL_15 = _EVAL_5 & _EVAL_82;
  assign _EVAL_170 = ~_EVAL_108;
  assign _EVAL_75 = _EVAL_59 & _EVAL_196;
  assign _EVAL_80 = _EVAL_114 != _EVAL_16;
  assign _EVAL_88 = _EVAL_3 == 3'h6;
  assign _EVAL_82 = _EVAL_3 == 3'h1;
  assign _EVAL_84 = _EVAL_154 | _EVAL_184;
  assign _EVAL_20 = _EVAL_6 & _EVAL_180;
  assign _EVAL_34 = _EVAL_129 ? _EVAL_146 : 8'h0;
  assign _EVAL_56 = ~_EVAL_142;
  assign _EVAL_167 = ~_EVAL_156;
  assign _EVAL_70 = 8'h1 << _EVAL_11;
  assign _EVAL_89 = _EVAL_120[1];
  assign _EVAL_192 = _EVAL_120[0];
  assign _EVAL_66 = ~_EVAL_17;
  assign _EVAL_169 = _EVAL_5 & _EVAL_44;
  assign _EVAL_101 = _EVAL_7 == 3'h1;
  assign _EVAL_23 = _EVAL_7 == 3'h0;
  assign _EVAL_86 = ~_EVAL_122;
  assign _EVAL_156 = _EVAL <= 3'h4;
  assign _EVAL_35 = ~_EVAL_194;
  assign _EVAL_69 = ~_EVAL_51;
  assign _EVAL_60 = _EVAL_178 == 4'h0;
  assign _EVAL_119 = _EVAL_104 | _EVAL_25;
  assign _EVAL_160 = _EVAL_189 == 4'h0;
  assign _EVAL_110 = _EVAL_18[0];
  assign _EVAL_136 = _EVAL_192 & _EVAL_137;
  assign _EVAL_200 = _EVAL_91 - 1'h1;
  assign _EVAL_190 = _EVAL_33 | _EVAL_114;
  assign _EVAL_139 = _EVAL_37[0];
  assign _EVAL_105 = _EVAL_114 | _EVAL_33;
  assign _EVAL_164 = _EVAL_114 != 5'h0;
  assign _EVAL_124 = ~_EVAL_83;
  assign _EVAL_59 = _EVAL_13 & _EVAL_5;
  assign _EVAL_166 = _EVAL_154 | _EVAL_136;
  assign _EVAL_71 = ~_EVAL_201;
  assign _EVAL_188 = _EVAL_7 == 3'h4;
  assign _EVAL_19 = _EVAL_5 & _EVAL_163;
  assign _EVAL_45 = ~_EVAL_22;
  assign _EVAL_87 = {1'b0,$signed(_EVAL_47)};
  assign _EVAL_146 = 8'h1 << _EVAL_0;
  assign _EVAL_129 = _EVAL_59 & _EVAL_144;
  assign _EVAL_141 = _EVAL_3 == 3'h7;
  assign _EVAL_41 = 2'h1 << _EVAL_168;
  assign _EVAL_40 = _EVAL_3 == 3'h2;
  assign _EVAL_74 = ~_EVAL_149;
  assign _EVAL_137 = _EVAL_150 & _EVAL_86;
  assign _EVAL_168 = _EVAL_10[0];
  assign _EVAL_52 = _EVAL_143[0];
  assign _EVAL_165 = _EVAL_2 & _EVAL_6;
  assign _EVAL_115 = _EVAL_10 == _EVAL_134;
  assign _EVAL_145 = _EVAL_80 | _EVAL_113;
  assign _EVAL_97 = 5'h3 << _EVAL_10;
  assign _EVAL_185 = _EVAL == 3'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_32 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_33 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_39 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_48 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_51 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_57 = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_73 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_78 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_91 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_95 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_96 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_108 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_134 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_159 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_8) begin
    if (_EVAL_75) begin
      _EVAL_32 <= _EVAL_0;
    end
    _EVAL_33 <= _EVAL_190 & _EVAL_116;
    if (_EVAL_191) begin
      _EVAL_39 <= _EVAL_9;
    end
    if (_EVAL_42) begin
      _EVAL_48 <= 32'h0;
    end else begin
      _EVAL_48 <= _EVAL_175;
    end
    if (_EVAL_165) begin
      if (_EVAL_69) begin
        _EVAL_51 <= 1'h0;
      end else begin
        _EVAL_51 <= _EVAL_110;
      end
    end
    if (_EVAL_75) begin
      _EVAL_57 <= _EVAL_1;
    end
    if (_EVAL_75) begin
      _EVAL_73 <= _EVAL;
    end
    if (_EVAL_191) begin
      _EVAL_78 <= _EVAL_7;
    end
    if (_EVAL_59) begin
      if (_EVAL_144) begin
        _EVAL_91 <= 1'h0;
      end else begin
        _EVAL_91 <= _EVAL_125;
      end
    end
    if (_EVAL_75) begin
      _EVAL_95 <= _EVAL_3;
    end
    if (_EVAL_59) begin
      if (_EVAL_196) begin
        _EVAL_96 <= 1'h0;
      end else begin
        _EVAL_96 <= _EVAL_52;
      end
    end
    if (_EVAL_165) begin
      if (_EVAL_170) begin
        _EVAL_108 <= 1'h0;
      end else begin
        _EVAL_108 <= _EVAL_176;
      end
    end
    if (_EVAL_75) begin
      _EVAL_134 <= _EVAL_10;
    end
    if (_EVAL_191) begin
      _EVAL_159 <= _EVAL_11;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccf1561b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ae8322f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7bc5bce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba1b75e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11005592)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1cb998a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(900fca35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(428b0ef7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87e983f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca7c1036)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12c23952)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d31429d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23af42bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(205447f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dddfc867)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4144783a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(655caa4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(766ca263)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31668ac4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3fa20ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16db8ef4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(840dc32e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(614c2c58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32b4781e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e8999da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d63897cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c096dfd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8742a04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c444832)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74ea9711)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd91cd68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56818047)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef3e3366)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fab3db20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73eeb965)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81d432d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1971cb10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6e37d56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fe223f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89b2bbb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed4d2b11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3abde3a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc535e0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8cdd93f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa1ec43a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a6a7cf8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99542aca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f5c9cc7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcbce7ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57bf4dbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8eaf14a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd5e1c9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cc28306)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5c490ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6940c86b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f77a0b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3858f8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a440d73b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acd6be12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86076fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7ddbad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74f24815)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84ef941b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f50de34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(694b3aa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(310649e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c07a360c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(719ec368)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbee73ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f20b596)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(487a0621)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6540d3e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27398fe2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
