//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_44(
  input  [1:0]  _EVAL,
  input         _EVAL_0,
  output [2:0]  _EVAL_1,
  output        _EVAL_2,
  output        _EVAL_3,
  input         _EVAL_4,
  input  [31:0] _EVAL_5,
  input         _EVAL_6,
  output [31:0] _EVAL_7,
  input  [2:0]  _EVAL_8,
  output        _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  output [1:0]  _EVAL_12,
  output        _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  output        _EVAL_16,
  output        _EVAL_17,
  input  [3:0]  _EVAL_18,
  output [3:0]  _EVAL_19
);
  wire  _EVAL_20;
  reg [3:0] _EVAL_21 [0:1];
  reg [31:0] _RAND_0;
  wire [3:0] _EVAL_21__EVAL_22_data;
  wire  _EVAL_21__EVAL_22_addr;
  wire [3:0] _EVAL_21__EVAL_23_data;
  wire  _EVAL_21__EVAL_23_addr;
  wire  _EVAL_21__EVAL_23_mask;
  wire  _EVAL_21__EVAL_23_en;
  wire  _EVAL_24;
  reg  _EVAL_25 [0:1];
  reg [31:0] _RAND_1;
  wire  _EVAL_25__EVAL_26_data;
  wire  _EVAL_25__EVAL_26_addr;
  wire  _EVAL_25__EVAL_27_data;
  wire  _EVAL_25__EVAL_27_addr;
  wire  _EVAL_25__EVAL_27_mask;
  wire  _EVAL_25__EVAL_27_en;
  reg  _EVAL_28 [0:1];
  reg [31:0] _RAND_2;
  wire  _EVAL_28__EVAL_29_data;
  wire  _EVAL_28__EVAL_29_addr;
  wire  _EVAL_28__EVAL_30_data;
  wire  _EVAL_28__EVAL_30_addr;
  wire  _EVAL_28__EVAL_30_mask;
  wire  _EVAL_28__EVAL_30_en;
  reg  _EVAL_31;
  reg [31:0] _RAND_3;
  reg  _EVAL_32 [0:1];
  reg [31:0] _RAND_4;
  wire  _EVAL_32__EVAL_33_data;
  wire  _EVAL_32__EVAL_33_addr;
  wire  _EVAL_32__EVAL_34_data;
  wire  _EVAL_32__EVAL_34_addr;
  wire  _EVAL_32__EVAL_34_mask;
  wire  _EVAL_32__EVAL_34_en;
  wire [1:0] _EVAL_35;
  wire  _EVAL_36;
  reg  _EVAL_37 [0:1];
  reg [31:0] _RAND_5;
  wire  _EVAL_37__EVAL_38_data;
  wire  _EVAL_37__EVAL_38_addr;
  wire  _EVAL_37__EVAL_39_data;
  wire  _EVAL_37__EVAL_39_addr;
  wire  _EVAL_37__EVAL_39_mask;
  wire  _EVAL_37__EVAL_39_en;
  wire  _EVAL_41;
  wire [1:0] _EVAL_42;
  reg [1:0] _EVAL_44 [0:1];
  reg [31:0] _RAND_6;
  wire [1:0] _EVAL_44__EVAL_45_data;
  wire  _EVAL_44__EVAL_45_addr;
  wire [1:0] _EVAL_44__EVAL_46_data;
  wire  _EVAL_44__EVAL_46_addr;
  wire  _EVAL_44__EVAL_46_mask;
  wire  _EVAL_44__EVAL_46_en;
  reg  _EVAL_47;
  reg [31:0] _RAND_7;
  wire  _EVAL_48;
  reg  _EVAL_49;
  reg [31:0] _RAND_8;
  wire  _EVAL_50;
  wire  _EVAL_52;
  reg [2:0] _EVAL_53 [0:1];
  reg [31:0] _RAND_9;
  wire [2:0] _EVAL_53__EVAL_54_data;
  wire  _EVAL_53__EVAL_54_addr;
  wire [2:0] _EVAL_53__EVAL_55_data;
  wire  _EVAL_53__EVAL_55_addr;
  wire  _EVAL_53__EVAL_55_mask;
  wire  _EVAL_53__EVAL_55_en;
  wire  _EVAL_56;
  wire  _EVAL_57;
  reg [31:0] _EVAL_58 [0:1];
  reg [31:0] _RAND_10;
  wire [31:0] _EVAL_58__EVAL_59_data;
  wire  _EVAL_58__EVAL_59_addr;
  wire [31:0] _EVAL_58__EVAL_60_data;
  wire  _EVAL_58__EVAL_60_addr;
  wire  _EVAL_58__EVAL_60_mask;
  wire  _EVAL_58__EVAL_60_en;
  assign _EVAL_21__EVAL_22_addr = _EVAL_47;
  assign _EVAL_21__EVAL_22_data = _EVAL_21[_EVAL_21__EVAL_22_addr];
  assign _EVAL_21__EVAL_23_data = _EVAL_18;
  assign _EVAL_21__EVAL_23_addr = _EVAL_49;
  assign _EVAL_21__EVAL_23_mask = 1'h1;
  assign _EVAL_21__EVAL_23_en = _EVAL_13 & _EVAL_10;
  assign _EVAL_25__EVAL_26_addr = _EVAL_47;
  assign _EVAL_25__EVAL_26_data = _EVAL_25[_EVAL_25__EVAL_26_addr];
  assign _EVAL_25__EVAL_27_data = _EVAL_14;
  assign _EVAL_25__EVAL_27_addr = _EVAL_49;
  assign _EVAL_25__EVAL_27_mask = 1'h1;
  assign _EVAL_25__EVAL_27_en = _EVAL_13 & _EVAL_10;
  assign _EVAL_28__EVAL_29_addr = _EVAL_47;
  assign _EVAL_28__EVAL_29_data = _EVAL_28[_EVAL_28__EVAL_29_addr];
  assign _EVAL_28__EVAL_30_data = 1'h0;
  assign _EVAL_28__EVAL_30_addr = _EVAL_49;
  assign _EVAL_28__EVAL_30_mask = 1'h1;
  assign _EVAL_28__EVAL_30_en = _EVAL_13 & _EVAL_10;
  assign _EVAL_32__EVAL_33_addr = _EVAL_47;
  assign _EVAL_32__EVAL_33_data = _EVAL_32[_EVAL_32__EVAL_33_addr];
  assign _EVAL_32__EVAL_34_data = _EVAL_0;
  assign _EVAL_32__EVAL_34_addr = _EVAL_49;
  assign _EVAL_32__EVAL_34_mask = 1'h1;
  assign _EVAL_32__EVAL_34_en = _EVAL_13 & _EVAL_10;
  assign _EVAL_37__EVAL_38_addr = _EVAL_47;
  assign _EVAL_37__EVAL_38_data = _EVAL_37[_EVAL_37__EVAL_38_addr];
  assign _EVAL_37__EVAL_39_data = _EVAL_6;
  assign _EVAL_37__EVAL_39_addr = _EVAL_49;
  assign _EVAL_37__EVAL_39_mask = 1'h1;
  assign _EVAL_37__EVAL_39_en = _EVAL_13 & _EVAL_10;
  assign _EVAL_44__EVAL_45_addr = _EVAL_47;
  assign _EVAL_44__EVAL_45_data = _EVAL_44[_EVAL_44__EVAL_45_addr];
  assign _EVAL_44__EVAL_46_data = _EVAL;
  assign _EVAL_44__EVAL_46_addr = _EVAL_49;
  assign _EVAL_44__EVAL_46_mask = 1'h1;
  assign _EVAL_44__EVAL_46_en = _EVAL_13 & _EVAL_10;
  assign _EVAL_53__EVAL_54_addr = _EVAL_47;
  assign _EVAL_53__EVAL_54_data = _EVAL_53[_EVAL_53__EVAL_54_addr];
  assign _EVAL_53__EVAL_55_data = _EVAL_8;
  assign _EVAL_53__EVAL_55_addr = _EVAL_49;
  assign _EVAL_53__EVAL_55_mask = 1'h1;
  assign _EVAL_53__EVAL_55_en = _EVAL_13 & _EVAL_10;
  assign _EVAL_58__EVAL_59_addr = _EVAL_47;
  assign _EVAL_58__EVAL_59_data = _EVAL_58[_EVAL_58__EVAL_59_addr];
  assign _EVAL_58__EVAL_60_data = _EVAL_5;
  assign _EVAL_58__EVAL_60_addr = _EVAL_49;
  assign _EVAL_58__EVAL_60_mask = 1'h1;
  assign _EVAL_58__EVAL_60_en = _EVAL_13 & _EVAL_10;
  assign _EVAL_24 = _EVAL_41 != _EVAL_56;
  assign _EVAL_42 = _EVAL_47 + 1'h1;
  assign _EVAL_41 = _EVAL_13 & _EVAL_10;
  assign _EVAL_9 = _EVAL_37__EVAL_38_data;
  assign _EVAL_35 = _EVAL_49 + 1'h1;
  assign _EVAL_3 = _EVAL_28__EVAL_29_data;
  assign _EVAL_19 = _EVAL_21__EVAL_22_data;
  assign _EVAL_1 = _EVAL_53__EVAL_54_data;
  assign _EVAL_36 = _EVAL_42[0];
  assign _EVAL_57 = _EVAL_35[0];
  assign _EVAL_13 = ~_EVAL_52;
  assign _EVAL_20 = ~_EVAL_31;
  assign _EVAL_56 = _EVAL_15 & _EVAL_17;
  assign _EVAL_7 = _EVAL_58__EVAL_59_data;
  assign _EVAL_48 = _EVAL_50 & _EVAL_20;
  assign _EVAL_17 = ~_EVAL_48;
  assign _EVAL_50 = _EVAL_49 == _EVAL_47;
  assign _EVAL_12 = _EVAL_44__EVAL_45_data;
  assign _EVAL_2 = _EVAL_25__EVAL_26_data;
  assign _EVAL_16 = _EVAL_32__EVAL_33_data;
  assign _EVAL_52 = _EVAL_50 & _EVAL_31;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_21[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_25[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_28[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_31 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_32[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_37[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_44[initvar] = _RAND_6[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_47 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_49 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_53[initvar] = _RAND_9[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_58[initvar] = _RAND_10[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_11) begin
    if(_EVAL_21__EVAL_23_en & _EVAL_21__EVAL_23_mask) begin
      _EVAL_21[_EVAL_21__EVAL_23_addr] <= _EVAL_21__EVAL_23_data;
    end
    if(_EVAL_25__EVAL_27_en & _EVAL_25__EVAL_27_mask) begin
      _EVAL_25[_EVAL_25__EVAL_27_addr] <= _EVAL_25__EVAL_27_data;
    end
    if(_EVAL_28__EVAL_30_en & _EVAL_28__EVAL_30_mask) begin
      _EVAL_28[_EVAL_28__EVAL_30_addr] <= _EVAL_28__EVAL_30_data;
    end
    if (_EVAL_4) begin
      _EVAL_31 <= 1'h0;
    end else if (_EVAL_24) begin
      _EVAL_31 <= _EVAL_41;
    end
    if(_EVAL_32__EVAL_34_en & _EVAL_32__EVAL_34_mask) begin
      _EVAL_32[_EVAL_32__EVAL_34_addr] <= _EVAL_32__EVAL_34_data;
    end
    if(_EVAL_37__EVAL_39_en & _EVAL_37__EVAL_39_mask) begin
      _EVAL_37[_EVAL_37__EVAL_39_addr] <= _EVAL_37__EVAL_39_data;
    end
    if(_EVAL_44__EVAL_46_en & _EVAL_44__EVAL_46_mask) begin
      _EVAL_44[_EVAL_44__EVAL_46_addr] <= _EVAL_44__EVAL_46_data;
    end
    if (_EVAL_4) begin
      _EVAL_47 <= 1'h0;
    end else if (_EVAL_56) begin
      _EVAL_47 <= _EVAL_36;
    end
    if (_EVAL_4) begin
      _EVAL_49 <= 1'h0;
    end else if (_EVAL_41) begin
      _EVAL_49 <= _EVAL_57;
    end
    if(_EVAL_53__EVAL_55_en & _EVAL_53__EVAL_55_mask) begin
      _EVAL_53[_EVAL_53__EVAL_55_addr] <= _EVAL_53__EVAL_55_data;
    end
    if(_EVAL_58__EVAL_60_en & _EVAL_58__EVAL_60_mask) begin
      _EVAL_58[_EVAL_58__EVAL_60_addr] <= _EVAL_58__EVAL_60_data;
    end
  end
endmodule
