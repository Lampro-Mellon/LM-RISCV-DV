//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_9(
  output        _EVAL,
  output        _EVAL_0,
  output [1:0]  _EVAL_1,
  output        _EVAL_2,
  input  [3:0]  _EVAL_3,
  output [31:0] _EVAL_4,
  output        _EVAL_5,
  output        _EVAL_6,
  output        _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  output        _EVAL_10,
  output [2:0]  _EVAL_11,
  output [1:0]  _EVAL_12,
  input         _EVAL_13,
  output        _EVAL_14,
  input         _EVAL_15,
  output [2:0]  _EVAL_16,
  input  [31:0] _EVAL_17,
  input  [31:0] _EVAL_18,
  output        _EVAL_19,
  output        _EVAL_20,
  output        _EVAL_21,
  input  [2:0]  _EVAL_22,
  input         _EVAL_23,
  output        _EVAL_24,
  input         _EVAL_25,
  output [2:0]  _EVAL_26,
  input  [3:0]  _EVAL_27,
  output [3:0]  _EVAL_28,
  input  [1:0]  _EVAL_29,
  input  [31:0] _EVAL_30,
  output        _EVAL_31,
  input  [3:0]  _EVAL_32,
  input         _EVAL_33,
  output        _EVAL_34,
  output        _EVAL_35,
  output [3:0]  _EVAL_36,
  output        _EVAL_37,
  input         _EVAL_38,
  output        _EVAL_39,
  output        _EVAL_40,
  output [31:0] _EVAL_41,
  output        _EVAL_42,
  input         _EVAL_43,
  input         _EVAL_44,
  output        _EVAL_45,
  input         _EVAL_46,
  input         _EVAL_47,
  output        _EVAL_48,
  output        _EVAL_49,
  input  [31:0] _EVAL_50,
  output        _EVAL_51,
  input         _EVAL_52,
  input         _EVAL_53,
  output        _EVAL_54,
  output        _EVAL_55,
  input         _EVAL_56,
  output [2:0]  _EVAL_57,
  output [3:0]  _EVAL_58,
  output        _EVAL_59,
  input  [31:0] _EVAL_60,
  output [3:0]  _EVAL_61,
  input         _EVAL_62,
  output        _EVAL_63,
  input         _EVAL_64,
  input         _EVAL_65,
  input         _EVAL_66,
  input  [2:0]  _EVAL_67,
  input         _EVAL_68,
  output        _EVAL_69,
  input         _EVAL_70,
  input  [1:0]  _EVAL_71,
  input         _EVAL_72,
  output        _EVAL_73,
  output [31:0] _EVAL_74,
  input  [2:0]  _EVAL_75,
  input         _EVAL_76,
  input  [2:0]  _EVAL_77,
  output        _EVAL_78,
  input  [2:0]  _EVAL_79,
  output        _EVAL_80,
  input         _EVAL_81,
  input         _EVAL_82,
  input         _EVAL_83,
  input         _EVAL_84,
  output        _EVAL_85,
  input         _EVAL_86,
  input         _EVAL_87,
  output [31:0] _EVAL_88,
  output [31:0] _EVAL_89,
  input         _EVAL_90,
  input  [3:0]  _EVAL_91,
  output        _EVAL_92,
  output [3:0]  _EVAL_93,
  output        _EVAL_94,
  input         _EVAL_95,
  input         _EVAL_96,
  output [31:0] _EVAL_97,
  input         _EVAL_98,
  output [2:0]  _EVAL_99,
  output [2:0]  _EVAL_100,
  output [3:0]  _EVAL_101,
  input  [3:0]  _EVAL_102,
  input         _EVAL_103,
  input  [31:0] _EVAL_104,
  input         _EVAL_105,
  input         _EVAL_106,
  input  [3:0]  _EVAL_107,
  input  [2:0]  _EVAL_108
);
  wire  buffer__EVAL;
  wire [2:0] buffer__EVAL_0;
  wire [2:0] buffer__EVAL_1;
  wire  buffer__EVAL_2;
  wire  buffer__EVAL_3;
  wire  buffer__EVAL_4;
  wire  buffer__EVAL_5;
  wire [31:0] buffer__EVAL_6;
  wire  buffer__EVAL_7;
  wire  buffer__EVAL_8;
  wire  buffer__EVAL_9;
  wire [31:0] buffer__EVAL_10;
  wire  buffer__EVAL_11;
  wire  buffer__EVAL_12;
  wire [31:0] buffer__EVAL_13;
  wire  buffer__EVAL_14;
  wire  buffer__EVAL_15;
  wire  buffer__EVAL_16;
  wire [1:0] buffer__EVAL_17;
  wire  buffer__EVAL_18;
  wire  buffer__EVAL_19;
  wire [31:0] buffer__EVAL_20;
  wire  buffer__EVAL_21;
  wire  buffer__EVAL_22;
  wire  buffer__EVAL_23;
  wire [3:0] buffer__EVAL_24;
  wire  buffer__EVAL_25;
  wire [31:0] buffer__EVAL_26;
  wire [3:0] buffer__EVAL_27;
  wire  buffer__EVAL_28;
  wire  buffer__EVAL_29;
  wire  buffer__EVAL_30;
  wire  buffer__EVAL_31;
  wire [1:0] buffer__EVAL_32;
  wire  buffer__EVAL_33;
  wire  buffer__EVAL_34;
  wire [3:0] buffer__EVAL_35;
  wire [2:0] buffer__EVAL_36;
  wire [3:0] buffer__EVAL_37;
  wire  buffer__EVAL_38;
  wire [3:0] buffer__EVAL_39;
  wire  buffer__EVAL_40;
  wire  buffer__EVAL_41;
  wire  buffer__EVAL_42;
  wire [3:0] buffer__EVAL_43;
  wire  buffer__EVAL_44;
  wire [2:0] buffer__EVAL_45;
  wire  buffer__EVAL_46;
  wire  buffer__EVAL_47;
  wire [1:0] buffer__EVAL_48;
  wire  buffer__EVAL_49;
  wire  buffer__EVAL_50;
  wire  buffer__EVAL_51;
  wire [3:0] buffer__EVAL_52;
  wire [31:0] buffer__EVAL_53;
  wire [2:0] buffer__EVAL_54;
  wire  buffer__EVAL_55;
  wire [2:0] buffer__EVAL_56;
  wire  buffer__EVAL_57;
  wire  buffer__EVAL_58;
  wire  buffer__EVAL_59;
  wire  buffer__EVAL_60;
  wire [2:0] buffer__EVAL_61;
  wire  buffer__EVAL_62;
  wire  buffer__EVAL_63;
  wire  buffer__EVAL_64;
  wire  buffer__EVAL_65;
  wire [31:0] buffer__EVAL_66;
  wire [3:0] buffer__EVAL_67;
  wire [2:0] buffer__EVAL_68;
  wire  buffer__EVAL_69;
  wire  buffer__EVAL_70;
  wire  buffer__EVAL_71;
  wire [2:0] buffer__EVAL_72;
  wire [2:0] buffer__EVAL_73;
  wire  buffer__EVAL_74;
  wire [31:0] buffer__EVAL_75;
  wire  buffer__EVAL_76;
  wire  buffer__EVAL_77;
  wire  buffer__EVAL_78;
  wire  buffer__EVAL_79;
  wire  buffer__EVAL_80;
  wire [1:0] buffer__EVAL_81;
  wire  buffer__EVAL_82;
  wire  buffer__EVAL_83;
  wire [31:0] buffer__EVAL_84;
  wire  buffer__EVAL_85;
  wire [3:0] buffer__EVAL_86;
  wire [2:0] buffer__EVAL_87;
  wire  buffer__EVAL_88;
  wire  buffer__EVAL_89;
  wire [3:0] buffer__EVAL_90;
  wire  buffer__EVAL_91;
  wire  buffer__EVAL_92;
  wire [2:0] buffer__EVAL_93;
  wire  buffer__EVAL_94;
  wire  buffer__EVAL_95;
  wire [31:0] buffer__EVAL_96;
  wire  buffer__EVAL_97;
  wire [31:0] buffer__EVAL_98;
  wire  buffer__EVAL_99;
  wire [3:0] buffer__EVAL_100;
  wire  buffer__EVAL_101;
  wire [3:0] buffer__EVAL_102;
  wire  buffer__EVAL_103;
  wire  buffer__EVAL_104;
  wire  buffer__EVAL_105;
  wire [31:0] buffer__EVAL_106;
  wire  buffer__EVAL_107;
  wire  buffer__EVAL_108;
  wire [2:0] fixer__EVAL;
  wire [1:0] fixer__EVAL_0;
  wire  fixer__EVAL_1;
  wire [2:0] fixer__EVAL_2;
  wire  fixer__EVAL_3;
  wire  fixer__EVAL_4;
  wire  fixer__EVAL_5;
  wire  fixer__EVAL_6;
  wire [1:0] fixer__EVAL_7;
  wire  fixer__EVAL_8;
  wire  fixer__EVAL_9;
  wire  fixer__EVAL_10;
  wire [2:0] fixer__EVAL_11;
  wire [3:0] fixer__EVAL_12;
  wire  fixer__EVAL_13;
  wire [2:0] fixer__EVAL_14;
  wire  fixer__EVAL_15;
  wire  fixer__EVAL_16;
  wire  fixer__EVAL_17;
  wire [3:0] fixer__EVAL_18;
  wire [3:0] fixer__EVAL_19;
  wire  fixer__EVAL_20;
  wire  fixer__EVAL_21;
  wire  fixer__EVAL_22;
  wire  fixer__EVAL_23;
  wire  fixer__EVAL_24;
  wire [31:0] fixer__EVAL_25;
  wire  fixer__EVAL_26;
  wire  fixer__EVAL_27;
  wire  fixer__EVAL_28;
  wire  fixer__EVAL_29;
  wire  fixer__EVAL_30;
  wire  fixer__EVAL_31;
  wire  fixer__EVAL_32;
  wire  fixer__EVAL_33;
  wire  fixer__EVAL_34;
  wire  fixer__EVAL_35;
  wire [31:0] fixer__EVAL_36;
  wire  fixer__EVAL_37;
  wire  fixer__EVAL_38;
  wire  fixer__EVAL_39;
  wire  fixer__EVAL_40;
  wire  fixer__EVAL_41;
  wire [2:0] fixer__EVAL_42;
  wire  fixer__EVAL_43;
  wire  fixer__EVAL_44;
  wire [31:0] fixer__EVAL_45;
  wire [2:0] fixer__EVAL_46;
  wire [31:0] fixer__EVAL_47;
  wire [2:0] fixer__EVAL_48;
  wire  fixer__EVAL_49;
  wire [31:0] fixer__EVAL_50;
  wire  fixer__EVAL_51;
  wire [31:0] fixer__EVAL_52;
  wire  fixer__EVAL_53;
  wire  fixer__EVAL_54;
  wire [31:0] fixer__EVAL_55;
  wire [3:0] fixer__EVAL_56;
  wire [2:0] fixer__EVAL_57;
  wire [2:0] fixer__EVAL_58;
  wire [3:0] fixer__EVAL_59;
  wire  fixer__EVAL_60;
  wire [3:0] fixer__EVAL_61;
  wire  fixer__EVAL_62;
  wire [1:0] fixer__EVAL_63;
  wire [3:0] fixer__EVAL_64;
  wire [3:0] fixer__EVAL_65;
  wire  fixer__EVAL_66;
  wire [31:0] fixer__EVAL_67;
  wire  fixer__EVAL_68;
  wire  fixer__EVAL_69;
  wire  fixer__EVAL_70;
  wire  fixer__EVAL_71;
  wire  fixer__EVAL_72;
  wire  fixer__EVAL_73;
  wire  fixer__EVAL_74;
  wire  fixer__EVAL_75;
  wire  fixer__EVAL_76;
  wire  fixer__EVAL_77;
  wire  fixer__EVAL_78;
  wire  fixer__EVAL_79;
  wire [31:0] fixer__EVAL_80;
  wire  fixer__EVAL_81;
  wire  fixer__EVAL_82;
  wire  fixer__EVAL_83;
  wire [2:0] fixer__EVAL_84;
  wire  fixer__EVAL_85;
  wire [3:0] fixer__EVAL_86;
  wire [3:0] fixer__EVAL_87;
  wire  fixer__EVAL_88;
  wire  fixer__EVAL_89;
  wire  fixer__EVAL_90;
  wire  fixer__EVAL_91;
  wire  fixer__EVAL_92;
  wire  fixer__EVAL_93;
  wire [3:0] fixer__EVAL_94;
  wire  fixer__EVAL_95;
  wire  fixer__EVAL_96;
  wire [3:0] fixer__EVAL_97;
  wire  fixer__EVAL_98;
  wire [31:0] fixer__EVAL_99;
  wire [2:0] fixer__EVAL_100;
  wire [31:0] fixer__EVAL_101;
  wire  fixer__EVAL_102;
  wire  fixer__EVAL_103;
  wire [2:0] fixer__EVAL_104;
  wire [31:0] fixer__EVAL_105;
  wire  fixer__EVAL_106;
  wire [1:0] fixer__EVAL_107;
  wire  fixer__EVAL_108;
  _EVAL_6 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32),
    ._EVAL_33(buffer__EVAL_33),
    ._EVAL_34(buffer__EVAL_34),
    ._EVAL_35(buffer__EVAL_35),
    ._EVAL_36(buffer__EVAL_36),
    ._EVAL_37(buffer__EVAL_37),
    ._EVAL_38(buffer__EVAL_38),
    ._EVAL_39(buffer__EVAL_39),
    ._EVAL_40(buffer__EVAL_40),
    ._EVAL_41(buffer__EVAL_41),
    ._EVAL_42(buffer__EVAL_42),
    ._EVAL_43(buffer__EVAL_43),
    ._EVAL_44(buffer__EVAL_44),
    ._EVAL_45(buffer__EVAL_45),
    ._EVAL_46(buffer__EVAL_46),
    ._EVAL_47(buffer__EVAL_47),
    ._EVAL_48(buffer__EVAL_48),
    ._EVAL_49(buffer__EVAL_49),
    ._EVAL_50(buffer__EVAL_50),
    ._EVAL_51(buffer__EVAL_51),
    ._EVAL_52(buffer__EVAL_52),
    ._EVAL_53(buffer__EVAL_53),
    ._EVAL_54(buffer__EVAL_54),
    ._EVAL_55(buffer__EVAL_55),
    ._EVAL_56(buffer__EVAL_56),
    ._EVAL_57(buffer__EVAL_57),
    ._EVAL_58(buffer__EVAL_58),
    ._EVAL_59(buffer__EVAL_59),
    ._EVAL_60(buffer__EVAL_60),
    ._EVAL_61(buffer__EVAL_61),
    ._EVAL_62(buffer__EVAL_62),
    ._EVAL_63(buffer__EVAL_63),
    ._EVAL_64(buffer__EVAL_64),
    ._EVAL_65(buffer__EVAL_65),
    ._EVAL_66(buffer__EVAL_66),
    ._EVAL_67(buffer__EVAL_67),
    ._EVAL_68(buffer__EVAL_68),
    ._EVAL_69(buffer__EVAL_69),
    ._EVAL_70(buffer__EVAL_70),
    ._EVAL_71(buffer__EVAL_71),
    ._EVAL_72(buffer__EVAL_72),
    ._EVAL_73(buffer__EVAL_73),
    ._EVAL_74(buffer__EVAL_74),
    ._EVAL_75(buffer__EVAL_75),
    ._EVAL_76(buffer__EVAL_76),
    ._EVAL_77(buffer__EVAL_77),
    ._EVAL_78(buffer__EVAL_78),
    ._EVAL_79(buffer__EVAL_79),
    ._EVAL_80(buffer__EVAL_80),
    ._EVAL_81(buffer__EVAL_81),
    ._EVAL_82(buffer__EVAL_82),
    ._EVAL_83(buffer__EVAL_83),
    ._EVAL_84(buffer__EVAL_84),
    ._EVAL_85(buffer__EVAL_85),
    ._EVAL_86(buffer__EVAL_86),
    ._EVAL_87(buffer__EVAL_87),
    ._EVAL_88(buffer__EVAL_88),
    ._EVAL_89(buffer__EVAL_89),
    ._EVAL_90(buffer__EVAL_90),
    ._EVAL_91(buffer__EVAL_91),
    ._EVAL_92(buffer__EVAL_92),
    ._EVAL_93(buffer__EVAL_93),
    ._EVAL_94(buffer__EVAL_94),
    ._EVAL_95(buffer__EVAL_95),
    ._EVAL_96(buffer__EVAL_96),
    ._EVAL_97(buffer__EVAL_97),
    ._EVAL_98(buffer__EVAL_98),
    ._EVAL_99(buffer__EVAL_99),
    ._EVAL_100(buffer__EVAL_100),
    ._EVAL_101(buffer__EVAL_101),
    ._EVAL_102(buffer__EVAL_102),
    ._EVAL_103(buffer__EVAL_103),
    ._EVAL_104(buffer__EVAL_104),
    ._EVAL_105(buffer__EVAL_105),
    ._EVAL_106(buffer__EVAL_106),
    ._EVAL_107(buffer__EVAL_107),
    ._EVAL_108(buffer__EVAL_108)
  );
  _EVAL_8 fixer (
    ._EVAL(fixer__EVAL),
    ._EVAL_0(fixer__EVAL_0),
    ._EVAL_1(fixer__EVAL_1),
    ._EVAL_2(fixer__EVAL_2),
    ._EVAL_3(fixer__EVAL_3),
    ._EVAL_4(fixer__EVAL_4),
    ._EVAL_5(fixer__EVAL_5),
    ._EVAL_6(fixer__EVAL_6),
    ._EVAL_7(fixer__EVAL_7),
    ._EVAL_8(fixer__EVAL_8),
    ._EVAL_9(fixer__EVAL_9),
    ._EVAL_10(fixer__EVAL_10),
    ._EVAL_11(fixer__EVAL_11),
    ._EVAL_12(fixer__EVAL_12),
    ._EVAL_13(fixer__EVAL_13),
    ._EVAL_14(fixer__EVAL_14),
    ._EVAL_15(fixer__EVAL_15),
    ._EVAL_16(fixer__EVAL_16),
    ._EVAL_17(fixer__EVAL_17),
    ._EVAL_18(fixer__EVAL_18),
    ._EVAL_19(fixer__EVAL_19),
    ._EVAL_20(fixer__EVAL_20),
    ._EVAL_21(fixer__EVAL_21),
    ._EVAL_22(fixer__EVAL_22),
    ._EVAL_23(fixer__EVAL_23),
    ._EVAL_24(fixer__EVAL_24),
    ._EVAL_25(fixer__EVAL_25),
    ._EVAL_26(fixer__EVAL_26),
    ._EVAL_27(fixer__EVAL_27),
    ._EVAL_28(fixer__EVAL_28),
    ._EVAL_29(fixer__EVAL_29),
    ._EVAL_30(fixer__EVAL_30),
    ._EVAL_31(fixer__EVAL_31),
    ._EVAL_32(fixer__EVAL_32),
    ._EVAL_33(fixer__EVAL_33),
    ._EVAL_34(fixer__EVAL_34),
    ._EVAL_35(fixer__EVAL_35),
    ._EVAL_36(fixer__EVAL_36),
    ._EVAL_37(fixer__EVAL_37),
    ._EVAL_38(fixer__EVAL_38),
    ._EVAL_39(fixer__EVAL_39),
    ._EVAL_40(fixer__EVAL_40),
    ._EVAL_41(fixer__EVAL_41),
    ._EVAL_42(fixer__EVAL_42),
    ._EVAL_43(fixer__EVAL_43),
    ._EVAL_44(fixer__EVAL_44),
    ._EVAL_45(fixer__EVAL_45),
    ._EVAL_46(fixer__EVAL_46),
    ._EVAL_47(fixer__EVAL_47),
    ._EVAL_48(fixer__EVAL_48),
    ._EVAL_49(fixer__EVAL_49),
    ._EVAL_50(fixer__EVAL_50),
    ._EVAL_51(fixer__EVAL_51),
    ._EVAL_52(fixer__EVAL_52),
    ._EVAL_53(fixer__EVAL_53),
    ._EVAL_54(fixer__EVAL_54),
    ._EVAL_55(fixer__EVAL_55),
    ._EVAL_56(fixer__EVAL_56),
    ._EVAL_57(fixer__EVAL_57),
    ._EVAL_58(fixer__EVAL_58),
    ._EVAL_59(fixer__EVAL_59),
    ._EVAL_60(fixer__EVAL_60),
    ._EVAL_61(fixer__EVAL_61),
    ._EVAL_62(fixer__EVAL_62),
    ._EVAL_63(fixer__EVAL_63),
    ._EVAL_64(fixer__EVAL_64),
    ._EVAL_65(fixer__EVAL_65),
    ._EVAL_66(fixer__EVAL_66),
    ._EVAL_67(fixer__EVAL_67),
    ._EVAL_68(fixer__EVAL_68),
    ._EVAL_69(fixer__EVAL_69),
    ._EVAL_70(fixer__EVAL_70),
    ._EVAL_71(fixer__EVAL_71),
    ._EVAL_72(fixer__EVAL_72),
    ._EVAL_73(fixer__EVAL_73),
    ._EVAL_74(fixer__EVAL_74),
    ._EVAL_75(fixer__EVAL_75),
    ._EVAL_76(fixer__EVAL_76),
    ._EVAL_77(fixer__EVAL_77),
    ._EVAL_78(fixer__EVAL_78),
    ._EVAL_79(fixer__EVAL_79),
    ._EVAL_80(fixer__EVAL_80),
    ._EVAL_81(fixer__EVAL_81),
    ._EVAL_82(fixer__EVAL_82),
    ._EVAL_83(fixer__EVAL_83),
    ._EVAL_84(fixer__EVAL_84),
    ._EVAL_85(fixer__EVAL_85),
    ._EVAL_86(fixer__EVAL_86),
    ._EVAL_87(fixer__EVAL_87),
    ._EVAL_88(fixer__EVAL_88),
    ._EVAL_89(fixer__EVAL_89),
    ._EVAL_90(fixer__EVAL_90),
    ._EVAL_91(fixer__EVAL_91),
    ._EVAL_92(fixer__EVAL_92),
    ._EVAL_93(fixer__EVAL_93),
    ._EVAL_94(fixer__EVAL_94),
    ._EVAL_95(fixer__EVAL_95),
    ._EVAL_96(fixer__EVAL_96),
    ._EVAL_97(fixer__EVAL_97),
    ._EVAL_98(fixer__EVAL_98),
    ._EVAL_99(fixer__EVAL_99),
    ._EVAL_100(fixer__EVAL_100),
    ._EVAL_101(fixer__EVAL_101),
    ._EVAL_102(fixer__EVAL_102),
    ._EVAL_103(fixer__EVAL_103),
    ._EVAL_104(fixer__EVAL_104),
    ._EVAL_105(fixer__EVAL_105),
    ._EVAL_106(fixer__EVAL_106),
    ._EVAL_107(fixer__EVAL_107),
    ._EVAL_108(fixer__EVAL_108)
  );
  assign fixer__EVAL_49 = buffer__EVAL_94;
  assign _EVAL_14 = buffer__EVAL_99;
  assign _EVAL_99 = buffer__EVAL_68;
  assign fixer__EVAL_75 = _EVAL_86;
  assign fixer__EVAL_58 = buffer__EVAL_45;
  assign buffer__EVAL_81 = _EVAL_29;
  assign fixer__EVAL_98 = buffer__EVAL_59;
  assign fixer__EVAL_32 = buffer__EVAL_57;
  assign _EVAL_20 = fixer__EVAL_53;
  assign _EVAL_69 = buffer__EVAL_15;
  assign fixer__EVAL_0 = buffer__EVAL_32;
  assign fixer__EVAL_30 = _EVAL_83;
  assign buffer__EVAL_38 = fixer__EVAL_102;
  assign buffer__EVAL_31 = fixer__EVAL_54;
  assign fixer__EVAL_101 = _EVAL_30;
  assign buffer__EVAL_34 = fixer__EVAL_81;
  assign fixer__EVAL_106 = _EVAL_9;
  assign _EVAL_0 = buffer__EVAL_83;
  assign buffer__EVAL_13 = _EVAL_104;
  assign fixer__EVAL_1 = _EVAL_62;
  assign buffer__EVAL_75 = fixer__EVAL_55;
  assign fixer__EVAL_70 = buffer__EVAL_4;
  assign fixer__EVAL_56 = buffer__EVAL_102;
  assign buffer__EVAL_69 = fixer__EVAL_5;
  assign buffer__EVAL_2 = fixer__EVAL_43;
  assign fixer__EVAL_7 = buffer__EVAL_48;
  assign buffer__EVAL_51 = fixer__EVAL_29;
  assign fixer__EVAL_103 = _EVAL_106;
  assign _EVAL_94 = fixer__EVAL_89;
  assign _EVAL_37 = fixer__EVAL_83;
  assign buffer__EVAL_63 = fixer__EVAL_91;
  assign buffer__EVAL_91 = _EVAL_72;
  assign buffer__EVAL_29 = fixer__EVAL_4;
  assign fixer__EVAL_76 = _EVAL_96;
  assign fixer__EVAL_20 = _EVAL_95;
  assign _EVAL_34 = buffer__EVAL_8;
  assign fixer__EVAL_3 = _EVAL_8;
  assign _EVAL_39 = buffer__EVAL_70;
  assign fixer__EVAL_17 = _EVAL_103;
  assign fixer__EVAL_68 = _EVAL_98;
  assign buffer__EVAL_18 = fixer__EVAL_37;
  assign _EVAL_51 = fixer__EVAL_31;
  assign buffer__EVAL_40 = _EVAL_98;
  assign fixer__EVAL_48 = _EVAL_79;
  assign _EVAL_63 = fixer__EVAL_28;
  assign fixer__EVAL_100 = _EVAL_108;
  assign fixer__EVAL_36 = buffer__EVAL_98;
  assign fixer__EVAL_108 = _EVAL_38;
  assign buffer__EVAL_56 = fixer__EVAL_46;
  assign _EVAL_55 = buffer__EVAL_47;
  assign buffer__EVAL_33 = _EVAL_62;
  assign _EVAL_101 = buffer__EVAL_24;
  assign buffer__EVAL_78 = fixer__EVAL_92;
  assign _EVAL_28 = fixer__EVAL_64;
  assign fixer__EVAL_22 = _EVAL_87;
  assign buffer__EVAL_1 = fixer__EVAL_2;
  assign fixer__EVAL_9 = buffer__EVAL_101;
  assign fixer__EVAL_10 = buffer__EVAL_7;
  assign buffer__EVAL_73 = fixer__EVAL_84;
  assign buffer__EVAL_0 = fixer__EVAL_11;
  assign fixer__EVAL_57 = _EVAL_75;
  assign buffer__EVAL_74 = fixer__EVAL_27;
  assign buffer__EVAL_100 = fixer__EVAL_19;
  assign fixer__EVAL_12 = _EVAL_107;
  assign _EVAL_16 = buffer__EVAL_36;
  assign fixer__EVAL_21 = buffer__EVAL_28;
  assign _EVAL_48 = fixer__EVAL_79;
  assign fixer__EVAL_16 = _EVAL_68;
  assign buffer__EVAL_97 = _EVAL_52;
  assign _EVAL_58 = buffer__EVAL_52;
  assign buffer__EVAL_61 = _EVAL_67;
  assign fixer__EVAL_87 = _EVAL_91;
  assign _EVAL_31 = buffer__EVAL_23;
  assign fixer__EVAL_62 = buffer__EVAL_55;
  assign fixer__EVAL_71 = buffer__EVAL_46;
  assign _EVAL_49 = buffer__EVAL_60;
  assign buffer__EVAL_85 = fixer__EVAL_8;
  assign buffer__EVAL_108 = fixer__EVAL_24;
  assign _EVAL_4 = buffer__EVAL_20;
  assign buffer__EVAL_54 = _EVAL_77;
  assign _EVAL_1 = fixer__EVAL_107;
  assign buffer__EVAL_92 = fixer__EVAL_35;
  assign _EVAL_19 = fixer__EVAL_60;
  assign _EVAL_35 = buffer__EVAL_64;
  assign buffer__EVAL_66 = fixer__EVAL_80;
  assign _EVAL_7 = buffer__EVAL_71;
  assign _EVAL_78 = fixer__EVAL_88;
  assign fixer__EVAL_14 = _EVAL_22;
  assign fixer__EVAL_104 = buffer__EVAL_72;
  assign buffer__EVAL_89 = _EVAL_105;
  assign _EVAL_5 = fixer__EVAL_15;
  assign fixer__EVAL_50 = _EVAL_17;
  assign _EVAL_74 = fixer__EVAL_52;
  assign _EVAL_88 = buffer__EVAL_106;
  assign _EVAL_85 = buffer__EVAL_95;
  assign buffer__EVAL_49 = fixer__EVAL_85;
  assign fixer__EVAL_94 = _EVAL_102;
  assign _EVAL_100 = buffer__EVAL_87;
  assign fixer__EVAL_51 = buffer__EVAL_19;
  assign buffer__EVAL_103 = _EVAL_66;
  assign _EVAL = buffer__EVAL_9;
  assign buffer__EVAL_16 = _EVAL_76;
  assign _EVAL_57 = fixer__EVAL_42;
  assign buffer__EVAL_96 = _EVAL_50;
  assign _EVAL_73 = buffer__EVAL_104;
  assign buffer__EVAL = fixer__EVAL_78;
  assign buffer__EVAL_90 = fixer__EVAL_18;
  assign buffer__EVAL_86 = fixer__EVAL_59;
  assign fixer__EVAL_26 = _EVAL_82;
  assign fixer__EVAL_90 = _EVAL_47;
  assign _EVAL_40 = buffer__EVAL_80;
  assign fixer__EVAL_96 = _EVAL_46;
  assign fixer__EVAL_40 = _EVAL_13;
  assign _EVAL_26 = fixer__EVAL;
  assign buffer__EVAL_43 = fixer__EVAL_61;
  assign _EVAL_2 = fixer__EVAL_82;
  assign _EVAL_6 = buffer__EVAL_11;
  assign _EVAL_12 = fixer__EVAL_63;
  assign buffer__EVAL_53 = fixer__EVAL_67;
  assign _EVAL_93 = buffer__EVAL_39;
  assign fixer__EVAL_34 = _EVAL_43;
  assign buffer__EVAL_76 = fixer__EVAL_39;
  assign _EVAL_36 = buffer__EVAL_35;
  assign fixer__EVAL_99 = _EVAL_18;
  assign buffer__EVAL_17 = _EVAL_71;
  assign fixer__EVAL_105 = buffer__EVAL_26;
  assign _EVAL_61 = fixer__EVAL_65;
  assign fixer__EVAL_23 = _EVAL_65;
  assign fixer__EVAL_38 = _EVAL_33;
  assign fixer__EVAL_33 = buffer__EVAL_88;
  assign _EVAL_11 = buffer__EVAL_93;
  assign _EVAL_10 = buffer__EVAL_3;
  assign fixer__EVAL_69 = _EVAL_64;
  assign fixer__EVAL_74 = _EVAL_53;
  assign fixer__EVAL_66 = buffer__EVAL_77;
  assign buffer__EVAL_25 = fixer__EVAL_13;
  assign _EVAL_97 = buffer__EVAL_84;
  assign _EVAL_42 = buffer__EVAL_22;
  assign buffer__EVAL_5 = fixer__EVAL_93;
  assign fixer__EVAL_86 = _EVAL_32;
  assign _EVAL_89 = buffer__EVAL_6;
  assign buffer__EVAL_67 = _EVAL_27;
  assign _EVAL_45 = buffer__EVAL_14;
  assign fixer__EVAL_97 = buffer__EVAL_27;
  assign _EVAL_59 = fixer__EVAL_73;
  assign buffer__EVAL_58 = _EVAL_23;
  assign buffer__EVAL_42 = _EVAL_56;
  assign buffer__EVAL_10 = fixer__EVAL_25;
  assign _EVAL_21 = buffer__EVAL_50;
  assign buffer__EVAL_30 = _EVAL_90;
  assign buffer__EVAL_44 = _EVAL_15;
  assign _EVAL_54 = fixer__EVAL_44;
  assign fixer__EVAL_72 = _EVAL_84;
  assign _EVAL_24 = buffer__EVAL_21;
  assign buffer__EVAL_79 = fixer__EVAL_95;
  assign buffer__EVAL_65 = _EVAL_44;
  assign buffer__EVAL_12 = _EVAL_70;
  assign _EVAL_92 = buffer__EVAL_107;
  assign buffer__EVAL_82 = fixer__EVAL_41;
  assign buffer__EVAL_105 = fixer__EVAL_77;
  assign _EVAL_80 = buffer__EVAL_62;
  assign fixer__EVAL_6 = _EVAL_25;
  assign buffer__EVAL_41 = _EVAL_81;
  assign _EVAL_41 = fixer__EVAL_45;
  assign buffer__EVAL_37 = _EVAL_3;
  assign fixer__EVAL_47 = _EVAL_60;
endmodule
