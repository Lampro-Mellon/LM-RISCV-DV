//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_180(
  input        _EVAL,
  input        _EVAL_0,
  output       _EVAL_1,
  output       _EVAL_2,
  output       _EVAL_3,
  input        _EVAL_4,
  input  [1:0] _EVAL_5,
  input        _EVAL_6,
  input        _EVAL_7,
  input        _EVAL_8
);
  reg  _EVAL_9;
  reg [31:0] _RAND_0;
  reg  _EVAL_10;
  reg [31:0] _RAND_1;
  wire  _EVAL_11;
  wire  _EVAL_12;
  wire  _EVAL_16;
  reg  _EVAL_20;
  reg [31:0] _RAND_2;
  wire  _EVAL_22;
  wire  _EVAL_23;
  reg  _EVAL_25;
  reg [31:0] _RAND_3;
  reg  _EVAL_26;
  reg [31:0] _RAND_4;
  wire [7:0] _EVAL_29;
  wire [31:0] _EVAL_33;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire [15:0] _EVAL_38;
  reg  _EVAL_40;
  reg [31:0] _RAND_5;
  wire  _EVAL_42;
  wire  _EVAL_44;
  reg  _EVAL_45;
  reg [31:0] _RAND_6;
  reg  _EVAL_51;
  reg [31:0] _RAND_7;
  reg  _EVAL_53;
  reg [31:0] _RAND_8;
  reg  _EVAL_54;
  reg [31:0] _RAND_9;
  wire  _EVAL_55;
  reg  _EVAL_56;
  reg [31:0] _RAND_10;
  reg  _EVAL_59;
  reg [31:0] _RAND_11;
  reg  _EVAL_60;
  reg [31:0] _RAND_12;
  wire  _EVAL_62;
  reg  _EVAL_63;
  reg [31:0] _RAND_13;
  reg  _EVAL_64;
  reg [31:0] _RAND_14;
  reg  _EVAL_65;
  reg [31:0] _RAND_15;
  wire  _EVAL_67;
  reg  _EVAL_68;
  reg [31:0] _RAND_16;
  reg  _EVAL_70;
  reg [31:0] _RAND_17;
  wire  _EVAL_75;
  reg  _EVAL_76;
  reg [31:0] _RAND_18;
  wire  _EVAL_77;
  reg  _EVAL_80;
  reg [31:0] _RAND_19;
  reg  _EVAL_83;
  reg [31:0] _RAND_20;
  wire  _EVAL_84;
  wire  _EVAL_90;
  wire  _EVAL_94;
  wire  _EVAL_96;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  reg  _EVAL_103;
  reg [31:0] _RAND_21;
  wire  _EVAL_106;
  reg  _EVAL_109;
  reg [31:0] _RAND_22;
  reg  _EVAL_110;
  reg [31:0] _RAND_23;
  reg  _EVAL_112;
  reg [31:0] _RAND_24;
  wire  _EVAL_115;
  reg  _EVAL_117;
  reg [31:0] _RAND_25;
  wire  _EVAL_118;
  reg  _EVAL_119;
  reg [31:0] _RAND_26;
  wire [7:0] _EVAL_120;
  wire  _EVAL_123;
  wire  _EVAL_128;
  wire  _EVAL_131;
  reg  _EVAL_132;
  reg [31:0] _RAND_27;
  wire [31:0] _EVAL_139;
  wire  _EVAL_140;
  reg  _EVAL_142;
  reg [31:0] _RAND_28;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  reg  _EVAL_146;
  reg [31:0] _RAND_29;
  wire  _EVAL_150;
  reg  _EVAL_152;
  reg [31:0] _RAND_30;
  reg  _EVAL_153;
  reg [31:0] _RAND_31;
  assign _EVAL_98 = _EVAL_33[12];
  assign _EVAL_150 = _EVAL_33[17];
  assign _EVAL_16 = _EVAL_33[16];
  assign _EVAL_62 = _EVAL_33[31];
  assign _EVAL_106 = _EVAL_33[10];
  assign _EVAL_115 = _EVAL_33[5];
  assign _EVAL_44 = _EVAL_33[22];
  assign _EVAL_140 = _EVAL_33[6];
  assign _EVAL_145 = _EVAL_33[2];
  assign _EVAL_38 = {_EVAL_119,_EVAL_63,_EVAL_83,_EVAL_153,_EVAL_64,_EVAL_152,_EVAL_54,_EVAL_146,_EVAL_29};
  assign _EVAL_94 = _EVAL_33[25];
  assign _EVAL_23 = _EVAL_33[24];
  assign _EVAL_131 = _EVAL_33[11];
  assign _EVAL_12 = _EVAL_33[7];
  assign _EVAL_22 = _EVAL_33[20];
  assign _EVAL_29 = {_EVAL_80,_EVAL_110,_EVAL_56,_EVAL_25,_EVAL_9,_EVAL_20,_EVAL_45,_EVAL_26};
  assign _EVAL_77 = _EVAL_33[9];
  assign _EVAL_11 = _EVAL_33[14];
  assign _EVAL_123 = _EVAL_33[3];
  assign _EVAL_42 = _EVAL_33[21];
  assign _EVAL_67 = _EVAL_33[28];
  assign _EVAL_55 = _EVAL_33[26];
  assign _EVAL_84 = _EVAL_33[19];
  assign _EVAL_120 = {_EVAL_10,_EVAL_59,_EVAL_70,_EVAL_68,_EVAL_112,_EVAL_132,_EVAL_65,_EVAL_60};
  assign _EVAL_100 = _EVAL_33[8];
  assign _EVAL_99 = _EVAL_33[15];
  assign _EVAL_144 = _EVAL_33[29];
  assign _EVAL_118 = _EVAL_33[18];
  assign _EVAL_90 = _EVAL_33[1];
  assign _EVAL_33 = {20'h5,_EVAL_5,6'h7,4'h1};
  assign _EVAL_75 = _EVAL_33[0];
  assign _EVAL_3 = _EVAL_8 ? 1'h0 : _EVAL_4;
  assign _EVAL_143 = _EVAL_33[27];
  assign _EVAL_1 = _EVAL_26;
  assign _EVAL_96 = _EVAL_33[13];
  assign _EVAL_128 = _EVAL_33[30];
  assign _EVAL_2 = _EVAL_139[16];
  assign _EVAL_139 = {_EVAL_103,_EVAL_117,_EVAL_51,_EVAL_142,_EVAL_40,_EVAL_109,_EVAL_76,_EVAL_53,_EVAL_120,_EVAL_38};
  assign _EVAL_36 = _EVAL_33[23];
  assign _EVAL_37 = _EVAL_33[4];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_9 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_10 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_20 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_25 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_26 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_40 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_45 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_51 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_53 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_54 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_56 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_59 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_60 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_63 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_64 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_65 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_68 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_70 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_76 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_80 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_83 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_103 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_109 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_110 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _EVAL_112 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _EVAL_117 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _EVAL_119 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _EVAL_132 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _EVAL_142 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _EVAL_146 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _EVAL_152 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _EVAL_153 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL) begin
    if (_EVAL_8) begin
      _EVAL_9 <= _EVAL_123;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_9 <= _EVAL_25;
      end
    end
    if (_EVAL_8) begin
      _EVAL_10 <= _EVAL_36;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_10 <= _EVAL_53;
      end
    end
    if (_EVAL_8) begin
      _EVAL_20 <= _EVAL_145;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_20 <= _EVAL_9;
      end
    end
    if (_EVAL_8) begin
      _EVAL_25 <= _EVAL_37;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_25 <= _EVAL_56;
      end
    end
    if (_EVAL_8) begin
      _EVAL_26 <= _EVAL_75;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_26 <= _EVAL_45;
      end
    end
    if (_EVAL_8) begin
      _EVAL_40 <= _EVAL_143;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_40 <= _EVAL_142;
      end
    end
    if (_EVAL_8) begin
      _EVAL_45 <= _EVAL_90;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_45 <= _EVAL_20;
      end
    end
    if (_EVAL_8) begin
      _EVAL_51 <= _EVAL_144;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_51 <= _EVAL_117;
      end
    end
    if (_EVAL_8) begin
      _EVAL_53 <= _EVAL_23;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_53 <= _EVAL_76;
      end
    end
    if (_EVAL_8) begin
      _EVAL_54 <= _EVAL_77;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_54 <= _EVAL_152;
      end
    end
    if (_EVAL_8) begin
      _EVAL_56 <= _EVAL_115;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_56 <= _EVAL_110;
      end
    end
    if (_EVAL_8) begin
      _EVAL_59 <= _EVAL_44;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_59 <= _EVAL_10;
      end
    end
    if (_EVAL_8) begin
      _EVAL_60 <= _EVAL_16;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_60 <= _EVAL_65;
      end
    end
    if (_EVAL_8) begin
      _EVAL_63 <= _EVAL_11;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_63 <= _EVAL_119;
      end
    end
    if (_EVAL_8) begin
      _EVAL_64 <= _EVAL_131;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_64 <= _EVAL_153;
      end
    end
    if (_EVAL_8) begin
      _EVAL_65 <= _EVAL_150;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_65 <= _EVAL_132;
      end
    end
    if (_EVAL_8) begin
      _EVAL_68 <= _EVAL_22;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_68 <= _EVAL_70;
      end
    end
    if (_EVAL_8) begin
      _EVAL_70 <= _EVAL_42;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_70 <= _EVAL_59;
      end
    end
    if (_EVAL_8) begin
      _EVAL_76 <= _EVAL_94;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_76 <= _EVAL_109;
      end
    end
    if (_EVAL_8) begin
      _EVAL_80 <= _EVAL_12;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_80 <= _EVAL_146;
      end
    end
    if (_EVAL_8) begin
      _EVAL_83 <= _EVAL_96;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_83 <= _EVAL_63;
      end
    end
    if (_EVAL_8) begin
      _EVAL_103 <= _EVAL_62;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_103 <= _EVAL_6;
      end
    end
    if (_EVAL_8) begin
      _EVAL_109 <= _EVAL_55;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_109 <= _EVAL_40;
      end
    end
    if (_EVAL_8) begin
      _EVAL_110 <= _EVAL_140;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_110 <= _EVAL_80;
      end
    end
    if (_EVAL_8) begin
      _EVAL_112 <= _EVAL_84;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_112 <= _EVAL_68;
      end
    end
    if (_EVAL_8) begin
      _EVAL_117 <= _EVAL_128;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_117 <= _EVAL_103;
      end
    end
    if (_EVAL_8) begin
      _EVAL_119 <= _EVAL_99;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_119 <= _EVAL_60;
      end
    end
    if (_EVAL_8) begin
      _EVAL_132 <= _EVAL_118;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_132 <= _EVAL_112;
      end
    end
    if (_EVAL_8) begin
      _EVAL_142 <= _EVAL_67;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_142 <= _EVAL_51;
      end
    end
    if (_EVAL_8) begin
      _EVAL_146 <= _EVAL_100;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_146 <= _EVAL_54;
      end
    end
    if (_EVAL_8) begin
      _EVAL_152 <= _EVAL_106;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_152 <= _EVAL_64;
      end
    end
    if (_EVAL_8) begin
      _EVAL_153 <= _EVAL_98;
    end else if (!(_EVAL_4)) begin
      if (_EVAL_7) begin
        _EVAL_153 <= _EVAL_83;
      end
    end
  end
endmodule
