//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_114_assert(
  input  [2:0]  _EVAL,
  input  [1:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input  [3:0]  _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [25:0] _EVAL_5,
  input  [1:0]  _EVAL_6,
  input         _EVAL_7,
  input  [2:0]  _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [2:0]  _EVAL_13,
  input         _EVAL_14
);
  wire [4:0] _EVAL_15;
  wire  _EVAL_16;
  wire [1:0] _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire [1:0] _EVAL_21;
  wire [4:0] _EVAL_22;
  wire  _EVAL_23;
  wire [1:0] _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  reg  _EVAL_27;
  reg [31:0] _RAND_0;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  reg  _EVAL_32;
  reg [31:0] _RAND_1;
  wire [26:0] _EVAL_33;
  wire  _EVAL_34;
  wire [1:0] _EVAL_35;
  reg [1:0] _EVAL_36;
  reg [31:0] _RAND_2;
  wire  _EVAL_37;
  wire  _EVAL_38;
  reg [4:0] _EVAL_39;
  reg [31:0] _RAND_3;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire [7:0] _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_46;
  wire [7:0] _EVAL_47;
  wire [26:0] _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire [3:0] _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire [1:0] _EVAL_58;
  wire  _EVAL_59;
  wire [1:0] _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  reg [2:0] _EVAL_64;
  reg [31:0] _RAND_4;
  wire [4:0] _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  reg [2:0] _EVAL_82;
  reg [31:0] _RAND_5;
  wire  _EVAL_83;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire [1:0] _EVAL_91;
  wire  _EVAL_92;
  wire [32:0] _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire [4:0] _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire [4:0] _EVAL_99;
  wire  _EVAL_100;
  reg [2:0] _EVAL_101;
  reg [31:0] _RAND_6;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  reg  _EVAL_114;
  reg [31:0] _RAND_7;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  reg [2:0] _EVAL_126;
  reg [31:0] _RAND_8;
  wire  _EVAL_127;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire [1:0] _EVAL_142;
  wire [7:0] _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire [26:0] _EVAL_146;
  wire [3:0] _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire [4:0] _EVAL_153;
  wire  _EVAL_154;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  reg [2:0] _EVAL_160;
  reg [31:0] _RAND_9;
  wire [25:0] _EVAL_161;
  wire  _EVAL_162;
  reg  _EVAL_163;
  reg [31:0] _RAND_10;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire [4:0] _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire [25:0] _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire [25:0] _EVAL_200;
  reg [31:0] _EVAL_201;
  reg [31:0] _RAND_11;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire [3:0] _EVAL_206;
  reg [1:0] _EVAL_207;
  reg [31:0] _RAND_12;
  wire  _EVAL_208;
  wire [7:0] _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire [4:0] _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire [3:0] _EVAL_221;
  wire  _EVAL_222;
  wire [31:0] _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  reg [25:0] _EVAL_232;
  reg [31:0] _RAND_13;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire [4:0] _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_241;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_123 = _EVAL_39 != 5'h0;
  assign _EVAL_88 = ~_EVAL_66;
  assign _EVAL_174 = _EVAL_9 & _EVAL_199;
  assign _EVAL_190 = _EVAL_55 == 4'h0;
  assign _EVAL_198 = _EVAL_97 | _EVAL_7;
  assign _EVAL_89 = _EVAL_228 | _EVAL_7;
  assign _EVAL_99 = _EVAL_96 >> _EVAL_8;
  assign _EVAL_113 = ~_EVAL_109;
  assign _EVAL_26 = _EVAL_85 | _EVAL_7;
  assign _EVAL_107 = ~_EVAL_222;
  assign _EVAL_53 = ~_EVAL_158;
  assign _EVAL_78 = ~_EVAL_164;
  assign _EVAL_168 = _EVAL_209[4:0];
  assign _EVAL_231 = _EVAL == 3'h5;
  assign _EVAL_228 = _EVAL_4 <= 3'h2;
  assign _EVAL_97 = _EVAL == _EVAL_64;
  assign _EVAL_109 = _EVAL_162 | _EVAL_7;
  assign _EVAL_142 = 2'h1 << _EVAL_132;
  assign _EVAL_46 = _EVAL_9 & _EVAL_37;
  assign _EVAL_102 = _EVAL_178 & _EVAL_151;
  assign _EVAL_145 = _EVAL_204 & _EVAL_216;
  assign _EVAL_224 = _EVAL_186 | _EVAL_7;
  assign _EVAL_209 = _EVAL_59 ? _EVAL_47 : 8'h0;
  assign _EVAL_151 = _EVAL_238 & _EVAL_211;
  assign _EVAL_241 = _EVAL_13 <= 3'h4;
  assign _EVAL_121 = _EVAL_149 | _EVAL_7;
  assign _EVAL_29 = ~_EVAL_177;
  assign _EVAL_86 = _EVAL_13 == _EVAL_126;
  assign _EVAL_172 = ~_EVAL_63;
  assign _EVAL_66 = _EVAL_182 | _EVAL_7;
  assign _EVAL_127 = _EVAL_12 <= 3'h6;
  assign _EVAL_69 = _EVAL_21[0];
  assign _EVAL_196 = _EVAL_8 <= 3'h4;
  assign _EVAL_54 = _EVAL == 3'h7;
  assign _EVAL_184 = $signed(_EVAL_146) == 27'sh0;
  assign _EVAL_43 = _EVAL_9 & _EVAL_110;
  assign _EVAL_148 = _EVAL_5[1];
  assign _EVAL_17 = _EVAL_114 - 1'h1;
  assign _EVAL_226 = ~_EVAL_111;
  assign _EVAL_41 = _EVAL_86 | _EVAL_7;
  assign _EVAL_208 = _EVAL_12 == 3'h6;
  assign _EVAL_193 = _EVAL_9 & _EVAL_175;
  assign _EVAL_176 = ~_EVAL_141;
  assign _EVAL_171 = ~_EVAL_233;
  assign _EVAL_162 = _EVAL_4 == _EVAL_101;
  assign _EVAL_140 = _EVAL_168 != _EVAL_153;
  assign _EVAL_125 = _EVAL_50 | _EVAL_7;
  assign _EVAL_44 = _EVAL == 3'h1;
  assign _EVAL_183 = _EVAL_106 | _EVAL_7;
  assign _EVAL_62 = _EVAL_119 | _EVAL_7;
  assign _EVAL_161 = _EVAL_5 & _EVAL_173;
  assign _EVAL_191 = _EVAL_17[0];
  assign _EVAL_170 = ~_EVAL_179;
  assign _EVAL_81 = ~_EVAL_62;
  assign _EVAL_25 = _EVAL_12 == 3'h1;
  assign _EVAL_230 = _EVAL_11 & _EVAL_214;
  assign _EVAL_51 = ~_EVAL_67;
  assign _EVAL_115 = plusarg_reader_out == 32'h0;
  assign _EVAL_177 = _EVAL_196 | _EVAL_7;
  assign _EVAL_77 = _EVAL_11 & _EVAL_28;
  assign _EVAL_52 = _EVAL_6 <= 2'h2;
  assign _EVAL_136 = _EVAL_9 & _EVAL_44;
  assign _EVAL_20 = _EVAL_192 & _EVAL_238;
  assign _EVAL_72 = _EVAL_241 | _EVAL_7;
  assign _EVAL_200 = _EVAL_5 ^ 26'h2000000;
  assign _EVAL_217 = 5'h3 << _EVAL_6;
  assign _EVAL_212 = _EVAL_91[0];
  assign _EVAL_37 = _EVAL == 3'h3;
  assign _EVAL_175 = _EVAL == 3'h0;
  assign _EVAL_57 = _EVAL_227 | _EVAL_7;
  assign _EVAL_154 = _EVAL_166 | _EVAL_7;
  assign _EVAL_35 = ~_EVAL_58;
  assign _EVAL_103 = _EVAL_130 | _EVAL_20;
  assign _EVAL_238 = ~_EVAL_148;
  assign _EVAL_138 = _EVAL_103 | _EVAL_112;
  assign _EVAL_65 = _EVAL_39 | _EVAL_168;
  assign _EVAL_237 = _EVAL_65 & _EVAL_22;
  assign _EVAL_75 = _EVAL_3 == _EVAL_147;
  assign _EVAL_71 = ~_EVAL_154;
  assign _EVAL_83 = _EVAL_238 & _EVAL_49;
  assign _EVAL_111 = _EVAL_18 | _EVAL_7;
  assign _EVAL_188 = _EVAL_31 & _EVAL_104;
  assign _EVAL_159 = _EVAL_178 & _EVAL_117;
  assign _EVAL_166 = _EVAL_4 <= 3'h1;
  assign _EVAL_122 = ~_EVAL_123;
  assign _EVAL_22 = ~_EVAL_153;
  assign _EVAL_195 = _EVAL_168 != 5'h0;
  assign _EVAL_194 = ~_EVAL_89;
  assign _EVAL_173 = {{24'd0}, _EVAL_35};
  assign _EVAL_219 = ~_EVAL_80;
  assign _EVAL_63 = _EVAL_75 | _EVAL_7;
  assign _EVAL_117 = _EVAL_148 & _EVAL_211;
  assign _EVAL_34 = ~_EVAL_152;
  assign _EVAL_48 = $signed(_EVAL_33) & -27'sh1000000;
  assign _EVAL_150 = ~_EVAL_183;
  assign _EVAL_116 = _EVAL_148 & _EVAL_49;
  assign _EVAL_165 = _EVAL_205 | _EVAL_108;
  assign _EVAL_47 = 8'h1 << _EVAL_13;
  assign _EVAL_31 = _EVAL_14 & _EVAL_11;
  assign _EVAL_169 = _EVAL_11 & _EVAL_208;
  assign _EVAL_181 = ~_EVAL_57;
  assign _EVAL_15 = _EVAL_39 >> _EVAL_13;
  assign _EVAL_50 = _EVAL_0 == _EVAL_36;
  assign _EVAL_94 = _EVAL_157 | _EVAL_7;
  assign _EVAL_93 = _EVAL_201 + 32'h1;
  assign _EVAL_110 = ~_EVAL_216;
  assign _EVAL_55 = _EVAL_3 & _EVAL_221;
  assign _EVAL_106 = _EVAL_140 | _EVAL_124;
  assign _EVAL_61 = _EVAL_11 & _EVAL_70;
  assign _EVAL_85 = _EVAL_0 >= 2'h2;
  assign _EVAL_157 = _EVAL_206 == 4'h0;
  assign _EVAL_143 = 8'h1 << _EVAL_8;
  assign _EVAL_206 = ~_EVAL_3;
  assign _EVAL_178 = _EVAL_60[0];
  assign _EVAL_24 = _EVAL_27 - 1'h1;
  assign _EVAL_225 = _EVAL_103 | _EVAL_102;
  assign _EVAL_234 = ~_EVAL_72;
  assign _EVAL_95 = _EVAL_192 & _EVAL_148;
  assign _EVAL_104 = ~_EVAL_163;
  assign _EVAL_147 = {_EVAL_202,_EVAL_165,_EVAL_225,_EVAL_138};
  assign _EVAL_76 = _EVAL_4 <= 3'h3;
  assign _EVAL_164 = _EVAL_130 | _EVAL_7;
  assign _EVAL_21 = _EVAL_32 - 1'h1;
  assign _EVAL_223 = _EVAL_93[31:0];
  assign _EVAL_130 = _EVAL_6 >= 2'h2;
  assign _EVAL_120 = _EVAL_9 & _EVAL_54;
  assign _EVAL_28 = _EVAL_12 == 3'h5;
  assign _EVAL_129 = ~_EVAL_7;
  assign _EVAL_40 = _EVAL == 3'h4;
  assign _EVAL_23 = _EVAL_127 | _EVAL_7;
  assign _EVAL_118 = ~_EVAL_208;
  assign _EVAL_199 = _EVAL == 3'h2;
  assign _EVAL_204 = _EVAL_10 & _EVAL_9;
  assign _EVAL_124 = ~_EVAL_195;
  assign _EVAL_203 = ~_EVAL_32;
  assign _EVAL_80 = _EVAL_105 | _EVAL_7;
  assign _EVAL_215 = _EVAL_6 == _EVAL_207;
  assign _EVAL_59 = _EVAL_204 & _EVAL_139;
  assign _EVAL_137 = _EVAL_11 & _EVAL_25;
  assign _EVAL_220 = _EVAL_9 & _EVAL_98;
  assign _EVAL_152 = _EVAL_156 | _EVAL_7;
  assign _EVAL_30 = _EVAL_134 | _EVAL_7;
  assign _EVAL_179 = _EVAL_213 | _EVAL_7;
  assign _EVAL_211 = _EVAL_5[0];
  assign _EVAL_216 = ~_EVAL_27;
  assign _EVAL_229 = ~_EVAL_121;
  assign _EVAL_189 = _EVAL_12 == 3'h2;
  assign _EVAL_16 = ~_EVAL_30;
  assign _EVAL_202 = _EVAL_205 | _EVAL_159;
  assign _EVAL_92 = _EVAL_9 & _EVAL_40;
  assign _EVAL_134 = _EVAL_4 != 3'h0;
  assign _EVAL_108 = _EVAL_178 & _EVAL_116;
  assign _EVAL_105 = _EVAL_8 == _EVAL_160;
  assign _EVAL_33 = {1'b0,$signed(_EVAL_200)};
  assign _EVAL_236 = ~_EVAL_1;
  assign _EVAL_112 = _EVAL_178 & _EVAL_83;
  assign _EVAL_67 = _EVAL_167 | _EVAL_7;
  assign _EVAL_214 = _EVAL_12 == 3'h0;
  assign _EVAL_131 = _EVAL_12 == 3'h4;
  assign _EVAL_167 = _EVAL_4 <= 3'h4;
  assign _EVAL_56 = _EVAL_11 & _EVAL_189;
  assign _EVAL_144 = _EVAL_204 | _EVAL_31;
  assign _EVAL_156 = _EVAL_5 == _EVAL_232;
  assign _EVAL_205 = _EVAL_130 | _EVAL_95;
  assign _EVAL_19 = _EVAL_24[0];
  assign _EVAL_233 = _EVAL_76 | _EVAL_7;
  assign _EVAL_141 = _EVAL_190 | _EVAL_7;
  assign _EVAL_68 = ~_EVAL_224;
  assign _EVAL_139 = ~_EVAL_114;
  assign _EVAL_180 = _EVAL_11 & _EVAL_131;
  assign _EVAL_58 = _EVAL_217[1:0];
  assign _EVAL_222 = _EVAL_215 | _EVAL_7;
  assign _EVAL_158 = _EVAL_236 | _EVAL_7;
  assign _EVAL_221 = ~_EVAL_147;
  assign _EVAL_91 = _EVAL_163 - 1'h1;
  assign _EVAL_185 = ~_EVAL_198;
  assign _EVAL_149 = ~_EVAL_133;
  assign _EVAL_227 = _EVAL_4 == 3'h0;
  assign _EVAL_213 = _EVAL_52 & _EVAL_184;
  assign _EVAL_192 = _EVAL_60[1];
  assign _EVAL_38 = ~_EVAL_41;
  assign _EVAL_218 = _EVAL_122 | _EVAL_115;
  assign _EVAL_146 = _EVAL_48;
  assign _EVAL_70 = ~_EVAL_203;
  assign _EVAL_197 = ~_EVAL_94;
  assign _EVAL_187 = ~_EVAL_26;
  assign _EVAL_155 = ~_EVAL_125;
  assign _EVAL_98 = _EVAL == 3'h6;
  assign _EVAL_182 = _EVAL_161 == 26'h0;
  assign _EVAL_210 = _EVAL_201 < plusarg_reader_out;
  assign _EVAL_96 = _EVAL_168 | _EVAL_39;
  assign _EVAL_87 = ~_EVAL_23;
  assign _EVAL_100 = _EVAL_9 & _EVAL_231;
  assign _EVAL_186 = _EVAL_12 == _EVAL_82;
  assign _EVAL_153 = _EVAL_42[4:0];
  assign _EVAL_132 = _EVAL_6[0];
  assign _EVAL_79 = _EVAL_31 & _EVAL_203;
  assign _EVAL_60 = _EVAL_142 | 2'h1;
  assign _EVAL_235 = _EVAL_188 & _EVAL_118;
  assign _EVAL_42 = _EVAL_235 ? _EVAL_143 : 8'h0;
  assign _EVAL_18 = _EVAL_99[0];
  assign _EVAL_133 = _EVAL_15[0];
  assign _EVAL_119 = _EVAL_218 | _EVAL_210;
  assign _EVAL_49 = ~_EVAL_211;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_27 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_32 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_36 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_39 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_64 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_82 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_101 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_114 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_126 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_160 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_163 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_201 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_207 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_232 = _RAND_13[25:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_2) begin
    if (_EVAL_7) begin
      _EVAL_27 <= 1'h0;
    end else if (_EVAL_204) begin
      if (_EVAL_216) begin
        _EVAL_27 <= 1'h0;
      end else begin
        _EVAL_27 <= _EVAL_19;
      end
    end
    if (_EVAL_7) begin
      _EVAL_32 <= 1'h0;
    end else if (_EVAL_31) begin
      if (_EVAL_203) begin
        _EVAL_32 <= 1'h0;
      end else begin
        _EVAL_32 <= _EVAL_69;
      end
    end
    if (_EVAL_79) begin
      _EVAL_36 <= _EVAL_0;
    end
    if (_EVAL_7) begin
      _EVAL_39 <= 5'h0;
    end else begin
      _EVAL_39 <= _EVAL_237;
    end
    if (_EVAL_145) begin
      _EVAL_64 <= _EVAL;
    end
    if (_EVAL_79) begin
      _EVAL_82 <= _EVAL_12;
    end
    if (_EVAL_145) begin
      _EVAL_101 <= _EVAL_4;
    end
    if (_EVAL_7) begin
      _EVAL_114 <= 1'h0;
    end else if (_EVAL_204) begin
      if (_EVAL_139) begin
        _EVAL_114 <= 1'h0;
      end else begin
        _EVAL_114 <= _EVAL_191;
      end
    end
    if (_EVAL_145) begin
      _EVAL_126 <= _EVAL_13;
    end
    if (_EVAL_79) begin
      _EVAL_160 <= _EVAL_8;
    end
    if (_EVAL_7) begin
      _EVAL_163 <= 1'h0;
    end else if (_EVAL_31) begin
      if (_EVAL_104) begin
        _EVAL_163 <= 1'h0;
      end else begin
        _EVAL_163 <= _EVAL_212;
      end
    end
    if (_EVAL_7) begin
      _EVAL_201 <= 32'h0;
    end else if (_EVAL_144) begin
      _EVAL_201 <= 32'h0;
    end else begin
      _EVAL_201 <= _EVAL_223;
    end
    if (_EVAL_145) begin
      _EVAL_207 <= _EVAL_6;
    end
    if (_EVAL_145) begin
      _EVAL_232 <= _EVAL_5;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae80f7af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71d73540)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74147629)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4704700c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ab7a1e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de6fde31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc4070ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6fccb9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fef715e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ced0571)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abad51ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(752eabab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23f4d11a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61dae4a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff12e8a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(944091)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b74616ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9358a263)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6442543)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddd60903)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c34288d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(767e12a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5728ce06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6489a64a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(896d69c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_16) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99a9e578)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34ef7c49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(984b065d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8796bab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b7e619)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba944d55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fc3677a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71d2630)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e32e690)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(510e88c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f18260c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(695e7e5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_16) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(660e194f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92e6253d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39ed4189)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eda7db81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12e3667f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5b36697)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(698dea1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b9815a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1acab565)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(832efffd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e6ba534)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0555d2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6fb9dc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba17ca29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a63f8ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63f8106a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(250d82e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9a8fa3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65240eab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d91b004)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c25c181)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d02b52e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dc5a233)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e2264d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c4d6ecd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1323d6cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44236504)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75408ea6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f184f8ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b56a075)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e4c3c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(347827ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee49fd02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a5f0980)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e83e55a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12216baf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
