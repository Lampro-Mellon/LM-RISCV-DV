//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_21(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  output        _EVAL_2,
  output [1:0]  _EVAL_3,
  input         _EVAL_4,
  output        _EVAL_5,
  input  [2:0]  _EVAL_6,
  output        _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  output [2:0]  _EVAL_10,
  output [2:0]  _EVAL_11,
  output [2:0]  _EVAL_12,
  input  [31:0] _EVAL_13,
  output        _EVAL_14,
  input         _EVAL_15,
  output        _EVAL_16,
  input  [2:0]  _EVAL_17,
  output [31:0] _EVAL_18
);
  reg [2:0] _EVAL_20 [0:1];
  reg [31:0] _RAND_0;
  wire [2:0] _EVAL_20__EVAL_21_data;
  wire  _EVAL_20__EVAL_21_addr;
  wire [2:0] _EVAL_20__EVAL_22_data;
  wire  _EVAL_20__EVAL_22_addr;
  wire  _EVAL_20__EVAL_22_mask;
  wire  _EVAL_20__EVAL_22_en;
  wire  _EVAL_23;
  wire  _EVAL_24;
  reg  _EVAL_25;
  reg [31:0] _RAND_1;
  reg [2:0] _EVAL_27 [0:1];
  reg [31:0] _RAND_2;
  wire [2:0] _EVAL_27__EVAL_28_data;
  wire  _EVAL_27__EVAL_28_addr;
  wire [2:0] _EVAL_27__EVAL_29_data;
  wire  _EVAL_27__EVAL_29_addr;
  wire  _EVAL_27__EVAL_29_mask;
  wire  _EVAL_27__EVAL_29_en;
  reg  _EVAL_30;
  reg [31:0] _RAND_3;
  reg  _EVAL_31 [0:1];
  reg [31:0] _RAND_4;
  wire  _EVAL_31__EVAL_32_data;
  wire  _EVAL_31__EVAL_32_addr;
  wire  _EVAL_31__EVAL_33_data;
  wire  _EVAL_31__EVAL_33_addr;
  wire  _EVAL_31__EVAL_33_mask;
  wire  _EVAL_31__EVAL_33_en;
  wire  _EVAL_34;
  wire [1:0] _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  reg [31:0] _EVAL_41 [0:1];
  reg [31:0] _RAND_5;
  wire [31:0] _EVAL_41__EVAL_42_data;
  wire  _EVAL_41__EVAL_42_addr;
  wire [31:0] _EVAL_41__EVAL_43_data;
  wire  _EVAL_41__EVAL_43_addr;
  wire  _EVAL_41__EVAL_43_mask;
  wire  _EVAL_41__EVAL_43_en;
  reg  _EVAL_44;
  reg [31:0] _RAND_6;
  wire  _EVAL_45;
  reg [1:0] _EVAL_46 [0:1];
  reg [31:0] _RAND_7;
  wire [1:0] _EVAL_46__EVAL_47_data;
  wire  _EVAL_46__EVAL_47_addr;
  wire [1:0] _EVAL_46__EVAL_48_data;
  wire  _EVAL_46__EVAL_48_addr;
  wire  _EVAL_46__EVAL_48_mask;
  wire  _EVAL_46__EVAL_48_en;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  reg [2:0] _EVAL_52 [0:1];
  reg [31:0] _RAND_8;
  wire [2:0] _EVAL_52__EVAL_53_data;
  wire  _EVAL_52__EVAL_53_addr;
  wire [2:0] _EVAL_52__EVAL_54_data;
  wire  _EVAL_52__EVAL_54_addr;
  wire  _EVAL_52__EVAL_54_mask;
  wire  _EVAL_52__EVAL_54_en;
  wire  _EVAL_55;
  wire  _EVAL_56;
  reg  _EVAL_57 [0:1];
  reg [31:0] _RAND_9;
  wire  _EVAL_57__EVAL_58_data;
  wire  _EVAL_57__EVAL_58_addr;
  wire  _EVAL_57__EVAL_59_data;
  wire  _EVAL_57__EVAL_59_addr;
  wire  _EVAL_57__EVAL_59_mask;
  wire  _EVAL_57__EVAL_59_en;
  reg  _EVAL_60 [0:1];
  reg [31:0] _RAND_10;
  wire  _EVAL_60__EVAL_61_data;
  wire  _EVAL_60__EVAL_61_addr;
  wire  _EVAL_60__EVAL_62_data;
  wire  _EVAL_60__EVAL_62_addr;
  wire  _EVAL_60__EVAL_62_mask;
  wire  _EVAL_60__EVAL_62_en;
  wire [1:0] _EVAL_63;
  assign _EVAL_20__EVAL_21_addr = _EVAL_25;
  assign _EVAL_20__EVAL_21_data = _EVAL_20[_EVAL_20__EVAL_21_addr];
  assign _EVAL_20__EVAL_22_data = _EVAL_6;
  assign _EVAL_20__EVAL_22_addr = _EVAL_30;
  assign _EVAL_20__EVAL_22_mask = 1'h1;
  assign _EVAL_20__EVAL_22_en = _EVAL_50 ? _EVAL_40 : _EVAL_49;
  assign _EVAL_27__EVAL_28_addr = _EVAL_25;
  assign _EVAL_27__EVAL_28_data = _EVAL_27[_EVAL_27__EVAL_28_addr];
  assign _EVAL_27__EVAL_29_data = _EVAL_17;
  assign _EVAL_27__EVAL_29_addr = _EVAL_30;
  assign _EVAL_27__EVAL_29_mask = 1'h1;
  assign _EVAL_27__EVAL_29_en = _EVAL_50 ? _EVAL_40 : _EVAL_49;
  assign _EVAL_31__EVAL_32_addr = _EVAL_25;
  assign _EVAL_31__EVAL_32_data = _EVAL_31[_EVAL_31__EVAL_32_addr];
  assign _EVAL_31__EVAL_33_data = 1'h0;
  assign _EVAL_31__EVAL_33_addr = _EVAL_30;
  assign _EVAL_31__EVAL_33_mask = 1'h1;
  assign _EVAL_31__EVAL_33_en = _EVAL_50 ? _EVAL_40 : _EVAL_49;
  assign _EVAL_41__EVAL_42_addr = _EVAL_25;
  assign _EVAL_41__EVAL_42_data = _EVAL_41[_EVAL_41__EVAL_42_addr];
  assign _EVAL_41__EVAL_43_data = _EVAL_13;
  assign _EVAL_41__EVAL_43_addr = _EVAL_30;
  assign _EVAL_41__EVAL_43_mask = 1'h1;
  assign _EVAL_41__EVAL_43_en = _EVAL_50 ? _EVAL_40 : _EVAL_49;
  assign _EVAL_46__EVAL_47_addr = _EVAL_25;
  assign _EVAL_46__EVAL_47_data = _EVAL_46[_EVAL_46__EVAL_47_addr];
  assign _EVAL_46__EVAL_48_data = 2'h0;
  assign _EVAL_46__EVAL_48_addr = _EVAL_30;
  assign _EVAL_46__EVAL_48_mask = 1'h1;
  assign _EVAL_46__EVAL_48_en = _EVAL_50 ? _EVAL_40 : _EVAL_49;
  assign _EVAL_52__EVAL_53_addr = _EVAL_25;
  assign _EVAL_52__EVAL_53_data = _EVAL_52[_EVAL_52__EVAL_53_addr];
  assign _EVAL_52__EVAL_54_data = _EVAL;
  assign _EVAL_52__EVAL_54_addr = _EVAL_30;
  assign _EVAL_52__EVAL_54_mask = 1'h1;
  assign _EVAL_52__EVAL_54_en = _EVAL_50 ? _EVAL_40 : _EVAL_49;
  assign _EVAL_57__EVAL_58_addr = _EVAL_25;
  assign _EVAL_57__EVAL_58_data = _EVAL_57[_EVAL_57__EVAL_58_addr];
  assign _EVAL_57__EVAL_59_data = _EVAL_15;
  assign _EVAL_57__EVAL_59_addr = _EVAL_30;
  assign _EVAL_57__EVAL_59_mask = 1'h1;
  assign _EVAL_57__EVAL_59_en = _EVAL_50 ? _EVAL_40 : _EVAL_49;
  assign _EVAL_60__EVAL_61_addr = _EVAL_25;
  assign _EVAL_60__EVAL_61_data = _EVAL_60[_EVAL_60__EVAL_61_addr];
  assign _EVAL_60__EVAL_62_data = _EVAL_8;
  assign _EVAL_60__EVAL_62_addr = _EVAL_30;
  assign _EVAL_60__EVAL_62_mask = 1'h1;
  assign _EVAL_60__EVAL_62_en = _EVAL_50 ? _EVAL_40 : _EVAL_49;
  assign _EVAL_35 = _EVAL_30 + 1'h1;
  assign _EVAL_40 = _EVAL_4 ? 1'h0 : _EVAL_49;
  assign _EVAL_55 = ~_EVAL_50;
  assign _EVAL_10 = _EVAL_50 ? _EVAL_17 : _EVAL_27__EVAL_28_data;
  assign _EVAL_39 = _EVAL_30 == _EVAL_25;
  assign _EVAL_16 = _EVAL_50 ? 1'h0 : _EVAL_31__EVAL_32_data;
  assign _EVAL_7 = _EVAL_1 | _EVAL_55;
  assign _EVAL_14 = _EVAL_50 ? _EVAL_8 : _EVAL_60__EVAL_61_data;
  assign _EVAL_63 = _EVAL_25 + 1'h1;
  assign _EVAL_24 = _EVAL_4 & _EVAL_7;
  assign _EVAL_12 = _EVAL_50 ? _EVAL_6 : _EVAL_20__EVAL_21_data;
  assign _EVAL_34 = _EVAL_45 != _EVAL_56;
  assign _EVAL_2 = _EVAL_50 ? _EVAL_15 : _EVAL_57__EVAL_58_data;
  assign _EVAL_38 = _EVAL_35[0];
  assign _EVAL_45 = _EVAL_50 ? _EVAL_40 : _EVAL_49;
  assign _EVAL_11 = _EVAL_50 ? _EVAL : _EVAL_52__EVAL_53_data;
  assign _EVAL_50 = _EVAL_39 & _EVAL_36;
  assign _EVAL_51 = _EVAL_63[0];
  assign _EVAL_56 = _EVAL_50 ? 1'h0 : _EVAL_24;
  assign _EVAL_49 = _EVAL_5 & _EVAL_1;
  assign _EVAL_23 = _EVAL_39 & _EVAL_44;
  assign _EVAL_3 = _EVAL_50 ? 2'h0 : _EVAL_46__EVAL_47_data;
  assign _EVAL_36 = ~_EVAL_44;
  assign _EVAL_5 = ~_EVAL_23;
  assign _EVAL_18 = _EVAL_50 ? _EVAL_13 : _EVAL_41__EVAL_42_data;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_20[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_25 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_27[initvar] = _RAND_2[2:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_30 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_31[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_41[initvar] = _RAND_5[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_44 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_46[initvar] = _RAND_7[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_52[initvar] = _RAND_8[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_57[initvar] = _RAND_9[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _EVAL_60[initvar] = _RAND_10[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_9) begin
    if(_EVAL_20__EVAL_22_en & _EVAL_20__EVAL_22_mask) begin
      _EVAL_20[_EVAL_20__EVAL_22_addr] <= _EVAL_20__EVAL_22_data;
    end
    if (_EVAL_0) begin
      _EVAL_25 <= 1'h0;
    end else if (_EVAL_56) begin
      _EVAL_25 <= _EVAL_51;
    end
    if(_EVAL_27__EVAL_29_en & _EVAL_27__EVAL_29_mask) begin
      _EVAL_27[_EVAL_27__EVAL_29_addr] <= _EVAL_27__EVAL_29_data;
    end
    if (_EVAL_0) begin
      _EVAL_30 <= 1'h0;
    end else if (_EVAL_45) begin
      _EVAL_30 <= _EVAL_38;
    end
    if(_EVAL_31__EVAL_33_en & _EVAL_31__EVAL_33_mask) begin
      _EVAL_31[_EVAL_31__EVAL_33_addr] <= _EVAL_31__EVAL_33_data;
    end
    if(_EVAL_41__EVAL_43_en & _EVAL_41__EVAL_43_mask) begin
      _EVAL_41[_EVAL_41__EVAL_43_addr] <= _EVAL_41__EVAL_43_data;
    end
    if (_EVAL_0) begin
      _EVAL_44 <= 1'h0;
    end else if (_EVAL_34) begin
      if (_EVAL_50) begin
        if (_EVAL_4) begin
          _EVAL_44 <= 1'h0;
        end else begin
          _EVAL_44 <= _EVAL_49;
        end
      end else begin
        _EVAL_44 <= _EVAL_49;
      end
    end
    if(_EVAL_46__EVAL_48_en & _EVAL_46__EVAL_48_mask) begin
      _EVAL_46[_EVAL_46__EVAL_48_addr] <= _EVAL_46__EVAL_48_data;
    end
    if(_EVAL_52__EVAL_54_en & _EVAL_52__EVAL_54_mask) begin
      _EVAL_52[_EVAL_52__EVAL_54_addr] <= _EVAL_52__EVAL_54_data;
    end
    if(_EVAL_57__EVAL_59_en & _EVAL_57__EVAL_59_mask) begin
      _EVAL_57[_EVAL_57__EVAL_59_addr] <= _EVAL_57__EVAL_59_data;
    end
    if(_EVAL_60__EVAL_62_en & _EVAL_60__EVAL_62_mask) begin
      _EVAL_60[_EVAL_60__EVAL_62_addr] <= _EVAL_60__EVAL_62_data;
    end
  end
endmodule
