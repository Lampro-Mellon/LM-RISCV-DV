//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_96(
  output [3:0]  _EVAL,
  input         _EVAL_0,
  output [2:0]  _EVAL_1,
  output [2:0]  _EVAL_2,
  input  [31:0] _EVAL_3,
  input  [2:0]  _EVAL_4,
  output [1:0]  _EVAL_5,
  output [31:0] _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input  [1:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  output        _EVAL_15,
  output        _EVAL_16,
  output [1:0]  _EVAL_17,
  output [31:0] _EVAL_18,
  input         _EVAL_19,
  input  [31:0] _EVAL_20,
  output        _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  output [1:0]  _EVAL_24,
  input         _EVAL_25,
  output [2:0]  _EVAL_26,
  output [29:0] _EVAL_27,
  input  [29:0] _EVAL_28,
  output        _EVAL_29,
  output        _EVAL_30,
  output        _EVAL_31,
  input  [2:0]  _EVAL_32,
  input  [3:0]  _EVAL_33
);
  wire  fragmenter__EVAL;
  wire [2:0] fragmenter__EVAL_0;
  wire [2:0] fragmenter__EVAL_1;
  wire  fragmenter__EVAL_2;
  wire [2:0] fragmenter__EVAL_3;
  wire [2:0] fragmenter__EVAL_4;
  wire [2:0] fragmenter__EVAL_5;
  wire [3:0] fragmenter__EVAL_6;
  wire  fragmenter__EVAL_7;
  wire [2:0] fragmenter__EVAL_8;
  wire  fragmenter__EVAL_9;
  wire [1:0] fragmenter__EVAL_10;
  wire  fragmenter__EVAL_11;
  wire [31:0] fragmenter__EVAL_12;
  wire [31:0] fragmenter__EVAL_13;
  wire  fragmenter__EVAL_14;
  wire [2:0] fragmenter__EVAL_15;
  wire  fragmenter__EVAL_16;
  wire [2:0] fragmenter__EVAL_17;
  wire  fragmenter__EVAL_18;
  wire [1:0] fragmenter__EVAL_19;
  wire  fragmenter__EVAL_20;
  wire  fragmenter__EVAL_21;
  wire  fragmenter__EVAL_22;
  wire [2:0] fragmenter__EVAL_23;
  wire  fragmenter__EVAL_24;
  wire [1:0] fragmenter__EVAL_25;
  wire  fragmenter__EVAL_26;
  wire  fragmenter__EVAL_27;
  wire  fragmenter__EVAL_28;
  wire [31:0] fragmenter__EVAL_29;
  wire [29:0] fragmenter__EVAL_30;
  wire [1:0] fragmenter__EVAL_31;
  wire [1:0] fragmenter__EVAL_32;
  wire  fragmenter__EVAL_33;
  wire  fragmenter__EVAL_34;
  wire  fragmenter__EVAL_35;
  wire  fragmenter__EVAL_36;
  wire [3:0] fragmenter__EVAL_37;
  wire  fragmenter__EVAL_38;
  wire  fragmenter__EVAL_39;
  wire  fragmenter__EVAL_40;
  wire  fragmenter__EVAL_41;
  wire [29:0] fragmenter__EVAL_42;
  wire [2:0] fragmenter__EVAL_43;
  wire [31:0] fragmenter__EVAL_44;
  wire  fragmenter__EVAL_45;
  wire [1:0] fragmenter__EVAL_46;
  wire  fragmenter__EVAL_47;
  wire  fragmenter__EVAL_48;
  wire  buffer__EVAL;
  wire [1:0] buffer__EVAL_0;
  wire [2:0] buffer__EVAL_1;
  wire [3:0] buffer__EVAL_2;
  wire  buffer__EVAL_3;
  wire [3:0] buffer__EVAL_4;
  wire  buffer__EVAL_5;
  wire  buffer__EVAL_6;
  wire  buffer__EVAL_7;
  wire [1:0] buffer__EVAL_8;
  wire  buffer__EVAL_9;
  wire  buffer__EVAL_10;
  wire  buffer__EVAL_11;
  wire [2:0] buffer__EVAL_12;
  wire  buffer__EVAL_13;
  wire  buffer__EVAL_14;
  wire  buffer__EVAL_15;
  wire  buffer__EVAL_16;
  wire  buffer__EVAL_17;
  wire  buffer__EVAL_18;
  wire [1:0] buffer__EVAL_19;
  wire [2:0] buffer__EVAL_20;
  wire  buffer__EVAL_21;
  wire [2:0] buffer__EVAL_22;
  wire [1:0] buffer__EVAL_23;
  wire [1:0] buffer__EVAL_24;
  wire [2:0] buffer__EVAL_25;
  wire [2:0] buffer__EVAL_26;
  wire  buffer__EVAL_27;
  wire  buffer__EVAL_28;
  wire  buffer__EVAL_29;
  wire [1:0] buffer__EVAL_30;
  wire [31:0] buffer__EVAL_31;
  wire [29:0] buffer__EVAL_32;
  wire  buffer__EVAL_33;
  wire [31:0] buffer__EVAL_34;
  wire [2:0] buffer__EVAL_35;
  wire  buffer__EVAL_36;
  wire  buffer__EVAL_37;
  wire  buffer__EVAL_38;
  wire  buffer__EVAL_39;
  wire [2:0] buffer__EVAL_40;
  wire  buffer__EVAL_41;
  wire  buffer__EVAL_42;
  wire [2:0] buffer__EVAL_43;
  wire [31:0] buffer__EVAL_44;
  wire [29:0] buffer__EVAL_45;
  wire [31:0] buffer__EVAL_46;
  wire [2:0] buffer__EVAL_47;
  wire  buffer__EVAL_48;
  wire [2:0] widget__EVAL;
  wire  widget__EVAL_0;
  wire [1:0] widget__EVAL_1;
  wire  widget__EVAL_2;
  wire  widget__EVAL_3;
  wire  widget__EVAL_4;
  wire [29:0] widget__EVAL_5;
  wire [2:0] widget__EVAL_6;
  wire [31:0] widget__EVAL_7;
  wire  widget__EVAL_8;
  wire  widget__EVAL_9;
  wire [1:0] widget__EVAL_10;
  wire  widget__EVAL_11;
  wire  widget__EVAL_12;
  wire  widget__EVAL_13;
  wire  widget__EVAL_14;
  wire [31:0] widget__EVAL_15;
  wire [1:0] widget__EVAL_16;
  wire [2:0] widget__EVAL_17;
  wire  widget__EVAL_18;
  wire [1:0] widget__EVAL_19;
  wire  widget__EVAL_20;
  wire  widget__EVAL_21;
  wire  widget__EVAL_22;
  wire  widget__EVAL_23;
  wire  widget__EVAL_24;
  wire [2:0] widget__EVAL_25;
  wire [31:0] widget__EVAL_26;
  wire  widget__EVAL_27;
  wire [2:0] widget__EVAL_28;
  wire  widget__EVAL_29;
  wire [31:0] widget__EVAL_30;
  wire [3:0] widget__EVAL_31;
  wire [2:0] widget__EVAL_32;
  wire  widget__EVAL_33;
  wire  widget__EVAL_34;
  wire [2:0] widget__EVAL_35;
  wire  widget__EVAL_36;
  wire  widget__EVAL_37;
  wire [3:0] widget__EVAL_38;
  wire [29:0] widget__EVAL_39;
  wire  widget__EVAL_40;
  wire [2:0] widget__EVAL_41;
  wire [1:0] widget__EVAL_42;
  wire  widget__EVAL_43;
  wire [1:0] widget__EVAL_44;
  wire  widget__EVAL_45;
  wire [2:0] widget__EVAL_46;
  wire  widget__EVAL_47;
  wire [2:0] widget__EVAL_48;
  wire [31:0] tl2ahb__EVAL;
  wire  tl2ahb__EVAL_0;
  wire  tl2ahb__EVAL_1;
  wire [2:0] tl2ahb__EVAL_2;
  wire [2:0] tl2ahb__EVAL_3;
  wire  tl2ahb__EVAL_4;
  wire  tl2ahb__EVAL_5;
  wire [29:0] tl2ahb__EVAL_6;
  wire [2:0] tl2ahb__EVAL_7;
  wire  tl2ahb__EVAL_8;
  wire  tl2ahb__EVAL_9;
  wire  tl2ahb__EVAL_10;
  wire [31:0] tl2ahb__EVAL_11;
  wire [2:0] tl2ahb__EVAL_12;
  wire  tl2ahb__EVAL_13;
  wire [31:0] tl2ahb__EVAL_14;
  wire  tl2ahb__EVAL_15;
  wire [3:0] tl2ahb__EVAL_16;
  wire [1:0] tl2ahb__EVAL_17;
  wire  tl2ahb__EVAL_18;
  wire  tl2ahb__EVAL_19;
  wire  tl2ahb__EVAL_20;
  wire [1:0] tl2ahb__EVAL_21;
  wire  tl2ahb__EVAL_22;
  wire [2:0] tl2ahb__EVAL_23;
  wire  tl2ahb__EVAL_24;
  wire [31:0] tl2ahb__EVAL_25;
  wire  tl2ahb__EVAL_26;
  wire [29:0] tl2ahb__EVAL_27;
  wire [1:0] tl2ahb__EVAL_28;
  wire  tl2ahb__EVAL_29;
  wire [3:0] tl2ahb__EVAL_30;
  wire [2:0] tl2ahb__EVAL_31;
  wire  tl2ahb__EVAL_32;
  wire [1:0] tl2ahb__EVAL_33;
  wire [1:0] buffer_1__EVAL;
  wire  buffer_1__EVAL_0;
  wire  buffer_1__EVAL_1;
  wire  buffer_1__EVAL_2;
  wire  buffer_1__EVAL_3;
  wire  buffer_1__EVAL_4;
  wire [3:0] buffer_1__EVAL_5;
  wire [2:0] buffer_1__EVAL_6;
  wire [31:0] buffer_1__EVAL_7;
  wire [31:0] buffer_1__EVAL_8;
  wire  buffer_1__EVAL_9;
  wire [2:0] buffer_1__EVAL_10;
  wire  buffer_1__EVAL_11;
  wire  buffer_1__EVAL_12;
  wire [29:0] buffer_1__EVAL_13;
  wire [1:0] buffer_1__EVAL_14;
  wire  buffer_1__EVAL_15;
  wire [2:0] buffer_1__EVAL_16;
  wire  buffer_1__EVAL_17;
  wire [29:0] buffer_1__EVAL_18;
  wire  buffer_1__EVAL_19;
  wire [2:0] buffer_1__EVAL_20;
  wire [1:0] buffer_1__EVAL_21;
  wire [2:0] buffer_1__EVAL_22;
  wire  buffer_1__EVAL_23;
  wire [3:0] buffer_1__EVAL_24;
  wire  buffer_1__EVAL_25;
  wire  buffer_1__EVAL_26;
  wire [31:0] buffer_1__EVAL_27;
  wire  buffer_1__EVAL_28;
  wire  buffer_1__EVAL_29;
  wire  buffer_1__EVAL_30;
  wire  buffer_1__EVAL_31;
  wire [2:0] buffer_1__EVAL_32;
  wire  buffer_1__EVAL_33;
  wire  buffer_1__EVAL_34;
  wire [2:0] buffer_1__EVAL_35;
  wire  buffer_1__EVAL_36;
  wire [1:0] buffer_1__EVAL_37;
  wire [2:0] buffer_1__EVAL_38;
  wire  buffer_1__EVAL_39;
  wire [1:0] buffer_1__EVAL_40;
  wire [1:0] buffer_1__EVAL_41;
  wire  buffer_1__EVAL_42;
  wire  buffer_1__EVAL_43;
  wire  buffer_1__EVAL_44;
  wire [2:0] buffer_1__EVAL_45;
  wire [31:0] buffer_1__EVAL_46;
  wire [2:0] buffer_1__EVAL_47;
  wire  buffer_1__EVAL_48;
  _EVAL_91 fragmenter (
    ._EVAL(fragmenter__EVAL),
    ._EVAL_0(fragmenter__EVAL_0),
    ._EVAL_1(fragmenter__EVAL_1),
    ._EVAL_2(fragmenter__EVAL_2),
    ._EVAL_3(fragmenter__EVAL_3),
    ._EVAL_4(fragmenter__EVAL_4),
    ._EVAL_5(fragmenter__EVAL_5),
    ._EVAL_6(fragmenter__EVAL_6),
    ._EVAL_7(fragmenter__EVAL_7),
    ._EVAL_8(fragmenter__EVAL_8),
    ._EVAL_9(fragmenter__EVAL_9),
    ._EVAL_10(fragmenter__EVAL_10),
    ._EVAL_11(fragmenter__EVAL_11),
    ._EVAL_12(fragmenter__EVAL_12),
    ._EVAL_13(fragmenter__EVAL_13),
    ._EVAL_14(fragmenter__EVAL_14),
    ._EVAL_15(fragmenter__EVAL_15),
    ._EVAL_16(fragmenter__EVAL_16),
    ._EVAL_17(fragmenter__EVAL_17),
    ._EVAL_18(fragmenter__EVAL_18),
    ._EVAL_19(fragmenter__EVAL_19),
    ._EVAL_20(fragmenter__EVAL_20),
    ._EVAL_21(fragmenter__EVAL_21),
    ._EVAL_22(fragmenter__EVAL_22),
    ._EVAL_23(fragmenter__EVAL_23),
    ._EVAL_24(fragmenter__EVAL_24),
    ._EVAL_25(fragmenter__EVAL_25),
    ._EVAL_26(fragmenter__EVAL_26),
    ._EVAL_27(fragmenter__EVAL_27),
    ._EVAL_28(fragmenter__EVAL_28),
    ._EVAL_29(fragmenter__EVAL_29),
    ._EVAL_30(fragmenter__EVAL_30),
    ._EVAL_31(fragmenter__EVAL_31),
    ._EVAL_32(fragmenter__EVAL_32),
    ._EVAL_33(fragmenter__EVAL_33),
    ._EVAL_34(fragmenter__EVAL_34),
    ._EVAL_35(fragmenter__EVAL_35),
    ._EVAL_36(fragmenter__EVAL_36),
    ._EVAL_37(fragmenter__EVAL_37),
    ._EVAL_38(fragmenter__EVAL_38),
    ._EVAL_39(fragmenter__EVAL_39),
    ._EVAL_40(fragmenter__EVAL_40),
    ._EVAL_41(fragmenter__EVAL_41),
    ._EVAL_42(fragmenter__EVAL_42),
    ._EVAL_43(fragmenter__EVAL_43),
    ._EVAL_44(fragmenter__EVAL_44),
    ._EVAL_45(fragmenter__EVAL_45),
    ._EVAL_46(fragmenter__EVAL_46),
    ._EVAL_47(fragmenter__EVAL_47),
    ._EVAL_48(fragmenter__EVAL_48)
  );
  _EVAL_89 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32),
    ._EVAL_33(buffer__EVAL_33),
    ._EVAL_34(buffer__EVAL_34),
    ._EVAL_35(buffer__EVAL_35),
    ._EVAL_36(buffer__EVAL_36),
    ._EVAL_37(buffer__EVAL_37),
    ._EVAL_38(buffer__EVAL_38),
    ._EVAL_39(buffer__EVAL_39),
    ._EVAL_40(buffer__EVAL_40),
    ._EVAL_41(buffer__EVAL_41),
    ._EVAL_42(buffer__EVAL_42),
    ._EVAL_43(buffer__EVAL_43),
    ._EVAL_44(buffer__EVAL_44),
    ._EVAL_45(buffer__EVAL_45),
    ._EVAL_46(buffer__EVAL_46),
    ._EVAL_47(buffer__EVAL_47),
    ._EVAL_48(buffer__EVAL_48)
  );
  _EVAL_93 widget (
    ._EVAL(widget__EVAL),
    ._EVAL_0(widget__EVAL_0),
    ._EVAL_1(widget__EVAL_1),
    ._EVAL_2(widget__EVAL_2),
    ._EVAL_3(widget__EVAL_3),
    ._EVAL_4(widget__EVAL_4),
    ._EVAL_5(widget__EVAL_5),
    ._EVAL_6(widget__EVAL_6),
    ._EVAL_7(widget__EVAL_7),
    ._EVAL_8(widget__EVAL_8),
    ._EVAL_9(widget__EVAL_9),
    ._EVAL_10(widget__EVAL_10),
    ._EVAL_11(widget__EVAL_11),
    ._EVAL_12(widget__EVAL_12),
    ._EVAL_13(widget__EVAL_13),
    ._EVAL_14(widget__EVAL_14),
    ._EVAL_15(widget__EVAL_15),
    ._EVAL_16(widget__EVAL_16),
    ._EVAL_17(widget__EVAL_17),
    ._EVAL_18(widget__EVAL_18),
    ._EVAL_19(widget__EVAL_19),
    ._EVAL_20(widget__EVAL_20),
    ._EVAL_21(widget__EVAL_21),
    ._EVAL_22(widget__EVAL_22),
    ._EVAL_23(widget__EVAL_23),
    ._EVAL_24(widget__EVAL_24),
    ._EVAL_25(widget__EVAL_25),
    ._EVAL_26(widget__EVAL_26),
    ._EVAL_27(widget__EVAL_27),
    ._EVAL_28(widget__EVAL_28),
    ._EVAL_29(widget__EVAL_29),
    ._EVAL_30(widget__EVAL_30),
    ._EVAL_31(widget__EVAL_31),
    ._EVAL_32(widget__EVAL_32),
    ._EVAL_33(widget__EVAL_33),
    ._EVAL_34(widget__EVAL_34),
    ._EVAL_35(widget__EVAL_35),
    ._EVAL_36(widget__EVAL_36),
    ._EVAL_37(widget__EVAL_37),
    ._EVAL_38(widget__EVAL_38),
    ._EVAL_39(widget__EVAL_39),
    ._EVAL_40(widget__EVAL_40),
    ._EVAL_41(widget__EVAL_41),
    ._EVAL_42(widget__EVAL_42),
    ._EVAL_43(widget__EVAL_43),
    ._EVAL_44(widget__EVAL_44),
    ._EVAL_45(widget__EVAL_45),
    ._EVAL_46(widget__EVAL_46),
    ._EVAL_47(widget__EVAL_47),
    ._EVAL_48(widget__EVAL_48)
  );
  _EVAL_85 tl2ahb (
    ._EVAL(tl2ahb__EVAL),
    ._EVAL_0(tl2ahb__EVAL_0),
    ._EVAL_1(tl2ahb__EVAL_1),
    ._EVAL_2(tl2ahb__EVAL_2),
    ._EVAL_3(tl2ahb__EVAL_3),
    ._EVAL_4(tl2ahb__EVAL_4),
    ._EVAL_5(tl2ahb__EVAL_5),
    ._EVAL_6(tl2ahb__EVAL_6),
    ._EVAL_7(tl2ahb__EVAL_7),
    ._EVAL_8(tl2ahb__EVAL_8),
    ._EVAL_9(tl2ahb__EVAL_9),
    ._EVAL_10(tl2ahb__EVAL_10),
    ._EVAL_11(tl2ahb__EVAL_11),
    ._EVAL_12(tl2ahb__EVAL_12),
    ._EVAL_13(tl2ahb__EVAL_13),
    ._EVAL_14(tl2ahb__EVAL_14),
    ._EVAL_15(tl2ahb__EVAL_15),
    ._EVAL_16(tl2ahb__EVAL_16),
    ._EVAL_17(tl2ahb__EVAL_17),
    ._EVAL_18(tl2ahb__EVAL_18),
    ._EVAL_19(tl2ahb__EVAL_19),
    ._EVAL_20(tl2ahb__EVAL_20),
    ._EVAL_21(tl2ahb__EVAL_21),
    ._EVAL_22(tl2ahb__EVAL_22),
    ._EVAL_23(tl2ahb__EVAL_23),
    ._EVAL_24(tl2ahb__EVAL_24),
    ._EVAL_25(tl2ahb__EVAL_25),
    ._EVAL_26(tl2ahb__EVAL_26),
    ._EVAL_27(tl2ahb__EVAL_27),
    ._EVAL_28(tl2ahb__EVAL_28),
    ._EVAL_29(tl2ahb__EVAL_29),
    ._EVAL_30(tl2ahb__EVAL_30),
    ._EVAL_31(tl2ahb__EVAL_31),
    ._EVAL_32(tl2ahb__EVAL_32),
    ._EVAL_33(tl2ahb__EVAL_33)
  );
  _EVAL_95 buffer_1 (
    ._EVAL(buffer_1__EVAL),
    ._EVAL_0(buffer_1__EVAL_0),
    ._EVAL_1(buffer_1__EVAL_1),
    ._EVAL_2(buffer_1__EVAL_2),
    ._EVAL_3(buffer_1__EVAL_3),
    ._EVAL_4(buffer_1__EVAL_4),
    ._EVAL_5(buffer_1__EVAL_5),
    ._EVAL_6(buffer_1__EVAL_6),
    ._EVAL_7(buffer_1__EVAL_7),
    ._EVAL_8(buffer_1__EVAL_8),
    ._EVAL_9(buffer_1__EVAL_9),
    ._EVAL_10(buffer_1__EVAL_10),
    ._EVAL_11(buffer_1__EVAL_11),
    ._EVAL_12(buffer_1__EVAL_12),
    ._EVAL_13(buffer_1__EVAL_13),
    ._EVAL_14(buffer_1__EVAL_14),
    ._EVAL_15(buffer_1__EVAL_15),
    ._EVAL_16(buffer_1__EVAL_16),
    ._EVAL_17(buffer_1__EVAL_17),
    ._EVAL_18(buffer_1__EVAL_18),
    ._EVAL_19(buffer_1__EVAL_19),
    ._EVAL_20(buffer_1__EVAL_20),
    ._EVAL_21(buffer_1__EVAL_21),
    ._EVAL_22(buffer_1__EVAL_22),
    ._EVAL_23(buffer_1__EVAL_23),
    ._EVAL_24(buffer_1__EVAL_24),
    ._EVAL_25(buffer_1__EVAL_25),
    ._EVAL_26(buffer_1__EVAL_26),
    ._EVAL_27(buffer_1__EVAL_27),
    ._EVAL_28(buffer_1__EVAL_28),
    ._EVAL_29(buffer_1__EVAL_29),
    ._EVAL_30(buffer_1__EVAL_30),
    ._EVAL_31(buffer_1__EVAL_31),
    ._EVAL_32(buffer_1__EVAL_32),
    ._EVAL_33(buffer_1__EVAL_33),
    ._EVAL_34(buffer_1__EVAL_34),
    ._EVAL_35(buffer_1__EVAL_35),
    ._EVAL_36(buffer_1__EVAL_36),
    ._EVAL_37(buffer_1__EVAL_37),
    ._EVAL_38(buffer_1__EVAL_38),
    ._EVAL_39(buffer_1__EVAL_39),
    ._EVAL_40(buffer_1__EVAL_40),
    ._EVAL_41(buffer_1__EVAL_41),
    ._EVAL_42(buffer_1__EVAL_42),
    ._EVAL_43(buffer_1__EVAL_43),
    ._EVAL_44(buffer_1__EVAL_44),
    ._EVAL_45(buffer_1__EVAL_45),
    ._EVAL_46(buffer_1__EVAL_46),
    ._EVAL_47(buffer_1__EVAL_47),
    ._EVAL_48(buffer_1__EVAL_48)
  );
  assign _EVAL_6 = tl2ahb__EVAL_11;
  assign buffer__EVAL_14 = _EVAL_8;
  assign buffer__EVAL_47 = fragmenter__EVAL_17;
  assign fragmenter__EVAL_36 = buffer__EVAL_37;
  assign _EVAL_15 = tl2ahb__EVAL_4;
  assign fragmenter__EVAL_3 = buffer__EVAL_12;
  assign _EVAL_30 = buffer_1__EVAL_0;
  assign buffer__EVAL_44 = tl2ahb__EVAL_25;
  assign widget__EVAL_28 = fragmenter__EVAL_1;
  assign buffer__EVAL_23 = tl2ahb__EVAL_28;
  assign buffer_1__EVAL_27 = widget__EVAL_7;
  assign buffer__EVAL_28 = _EVAL_12;
  assign _EVAL_16 = buffer_1__EVAL_25;
  assign buffer__EVAL_45 = fragmenter__EVAL_30;
  assign widget__EVAL_27 = fragmenter__EVAL_2;
  assign buffer__EVAL_17 = tl2ahb__EVAL_5;
  assign buffer__EVAL_29 = fragmenter__EVAL_21;
  assign _EVAL_24 = buffer_1__EVAL_14;
  assign widget__EVAL_4 = buffer_1__EVAL_33;
  assign buffer__EVAL_36 = fragmenter__EVAL_33;
  assign buffer__EVAL_11 = tl2ahb__EVAL_22;
  assign tl2ahb__EVAL_12 = buffer__EVAL_26;
  assign widget__EVAL_5 = buffer_1__EVAL_18;
  assign tl2ahb__EVAL_0 = buffer__EVAL_5;
  assign _EVAL_18 = buffer_1__EVAL_46;
  assign fragmenter__EVAL_23 = widget__EVAL_48;
  assign tl2ahb__EVAL_23 = buffer__EVAL_1;
  assign buffer_1__EVAL_1 = _EVAL_12;
  assign widget__EVAL_3 = buffer_1__EVAL_44;
  assign fragmenter__EVAL_29 = widget__EVAL_30;
  assign buffer_1__EVAL_43 = _EVAL_25;
  assign buffer__EVAL_25 = tl2ahb__EVAL_31;
  assign _EVAL_27 = tl2ahb__EVAL_27;
  assign buffer__EVAL_19 = fragmenter__EVAL_10;
  assign buffer_1__EVAL_32 = _EVAL_32;
  assign widget__EVAL_31 = buffer_1__EVAL_5;
  assign buffer__EVAL_7 = fragmenter__EVAL_34;
  assign _EVAL_29 = buffer_1__EVAL_11;
  assign buffer_1__EVAL_21 = _EVAL_11;
  assign _EVAL_17 = buffer_1__EVAL_37;
  assign buffer_1__EVAL_26 = widget__EVAL_47;
  assign widget__EVAL_6 = buffer_1__EVAL_10;
  assign buffer_1__EVAL_35 = _EVAL_7;
  assign tl2ahb__EVAL_2 = buffer__EVAL_35;
  assign buffer__EVAL_2 = fragmenter__EVAL_37;
  assign fragmenter__EVAL_27 = widget__EVAL_29;
  assign fragmenter__EVAL_8 = buffer__EVAL_43;
  assign widget__EVAL_44 = fragmenter__EVAL_31;
  assign buffer_1__EVAL_40 = widget__EVAL_42;
  assign buffer__EVAL_20 = fragmenter__EVAL_5;
  assign fragmenter__EVAL_11 = buffer__EVAL_3;
  assign buffer__EVAL_6 = tl2ahb__EVAL_10;
  assign tl2ahb__EVAL_29 = _EVAL_8;
  assign buffer_1__EVAL_20 = widget__EVAL_35;
  assign buffer_1__EVAL_7 = _EVAL_20;
  assign buffer_1__EVAL_12 = _EVAL_22;
  assign widget__EVAL_36 = fragmenter__EVAL_7;
  assign buffer__EVAL_9 = tl2ahb__EVAL_18;
  assign fragmenter__EVAL_6 = widget__EVAL_38;
  assign widget__EVAL_9 = buffer_1__EVAL_36;
  assign fragmenter__EVAL = widget__EVAL_22;
  assign buffer_1__EVAL_41 = widget__EVAL_16;
  assign buffer__EVAL_10 = fragmenter__EVAL_35;
  assign buffer_1__EVAL_17 = _EVAL_8;
  assign tl2ahb__EVAL_1 = buffer__EVAL_42;
  assign fragmenter__EVAL_46 = buffer__EVAL_30;
  assign widget__EVAL_46 = buffer_1__EVAL_16;
  assign fragmenter__EVAL_32 = buffer__EVAL_0;
  assign _EVAL_2 = buffer_1__EVAL_45;
  assign buffer_1__EVAL_28 = widget__EVAL_14;
  assign buffer__EVAL_21 = tl2ahb__EVAL_15;
  assign fragmenter__EVAL_9 = widget__EVAL_45;
  assign tl2ahb__EVAL_24 = buffer__EVAL_41;
  assign tl2ahb__EVAL_32 = _EVAL_10;
  assign buffer_1__EVAL_39 = widget__EVAL_23;
  assign tl2ahb__EVAL_14 = buffer__EVAL_34;
  assign buffer_1__EVAL_31 = _EVAL_0;
  assign widget__EVAL_26 = buffer_1__EVAL_8;
  assign widget__EVAL = buffer_1__EVAL_22;
  assign _EVAL = tl2ahb__EVAL_30;
  assign widget__EVAL_11 = buffer_1__EVAL_23;
  assign widget__EVAL_34 = _EVAL_12;
  assign fragmenter__EVAL_26 = widget__EVAL_20;
  assign buffer_1__EVAL_6 = widget__EVAL_32;
  assign fragmenter__EVAL_38 = _EVAL_12;
  assign fragmenter__EVAL_18 = widget__EVAL_13;
  assign tl2ahb__EVAL_13 = buffer__EVAL_15;
  assign buffer__EVAL_13 = fragmenter__EVAL_45;
  assign _EVAL_31 = buffer_1__EVAL_48;
  assign tl2ahb__EVAL_21 = buffer__EVAL_8;
  assign tl2ahb__EVAL_20 = buffer__EVAL_39;
  assign fragmenter__EVAL_19 = widget__EVAL_10;
  assign tl2ahb__EVAL_16 = buffer__EVAL_4;
  assign fragmenter__EVAL_16 = buffer__EVAL_27;
  assign buffer__EVAL_38 = fragmenter__EVAL_22;
  assign _EVAL_5 = tl2ahb__EVAL_33;
  assign widget__EVAL_1 = fragmenter__EVAL_25;
  assign widget__EVAL_12 = fragmenter__EVAL_47;
  assign tl2ahb__EVAL_9 = _EVAL_12;
  assign widget__EVAL_19 = buffer_1__EVAL;
  assign fragmenter__EVAL_39 = widget__EVAL_43;
  assign buffer_1__EVAL_13 = _EVAL_28;
  assign fragmenter__EVAL_48 = widget__EVAL_33;
  assign tl2ahb__EVAL_26 = buffer__EVAL_33;
  assign tl2ahb__EVAL_8 = _EVAL_23;
  assign fragmenter__EVAL_28 = buffer__EVAL;
  assign _EVAL_1 = tl2ahb__EVAL_7;
  assign buffer__EVAL_24 = tl2ahb__EVAL_17;
  assign widget__EVAL_18 = fragmenter__EVAL_41;
  assign buffer_1__EVAL_34 = _EVAL_13;
  assign tl2ahb__EVAL = _EVAL_3;
  assign fragmenter__EVAL_0 = widget__EVAL_41;
  assign buffer_1__EVAL_9 = _EVAL_19;
  assign buffer_1__EVAL_4 = widget__EVAL_2;
  assign buffer__EVAL_22 = fragmenter__EVAL_15;
  assign fragmenter__EVAL_42 = widget__EVAL_39;
  assign buffer__EVAL_40 = tl2ahb__EVAL_3;
  assign tl2ahb__EVAL_6 = buffer__EVAL_32;
  assign buffer_1__EVAL_29 = _EVAL_14;
  assign widget__EVAL_40 = _EVAL_8;
  assign widget__EVAL_8 = buffer_1__EVAL_42;
  assign fragmenter__EVAL_14 = _EVAL_8;
  assign buffer_1__EVAL_47 = _EVAL_4;
  assign fragmenter__EVAL_44 = buffer__EVAL_31;
  assign buffer_1__EVAL_24 = _EVAL_33;
  assign widget__EVAL_15 = fragmenter__EVAL_13;
  assign buffer__EVAL_48 = fragmenter__EVAL_24;
  assign buffer_1__EVAL_30 = widget__EVAL_24;
  assign fragmenter__EVAL_20 = buffer__EVAL_16;
  assign buffer_1__EVAL_2 = _EVAL_9;
  assign widget__EVAL_21 = buffer_1__EVAL_19;
  assign fragmenter__EVAL_4 = widget__EVAL_25;
  assign widget__EVAL_37 = buffer_1__EVAL_15;
  assign tl2ahb__EVAL_19 = buffer__EVAL_18;
  assign _EVAL_26 = buffer_1__EVAL_38;
  assign _EVAL_21 = buffer_1__EVAL_3;
  assign widget__EVAL_0 = fragmenter__EVAL_40;
  assign widget__EVAL_17 = fragmenter__EVAL_43;
  assign buffer__EVAL_46 = fragmenter__EVAL_12;
endmodule
