//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_116_assert(
  input           _EVAL_11,
  input           _EVAL_24,
  input  [2:0]    _EVAL_25,
  input  [1:0]    _EVAL_26,
  input           _EVAL_34,
  input  [2:0]    _EVAL_77,
  input  [2:0]    _EVAL_88,
  input           _EVAL_106,
  input           _EVAL_112,
  input  [3:0]    _EVAL_124,
  input  [25:0]   _EVAL_131,
  input           _EVAL_156,
  input           _EVAL_158,
  input           _EVAL_174,
  input           _EVAL_176,
  input           _EVAL_197,
  input           _EVAL_203,
  input           _EVAL_212,
  input           _EVAL_234,
  input           _EVAL_236,
  input           _EVAL_245,
  input           _EVAL_277,
  input           _EVAL_281,
  input           _EVAL_283,
  input           _EVAL_289,
  input           _EVAL_300,
  input           _EVAL_306,
  input           _EVAL_315,
  input           _EVAL_317,
  input           _EVAL_340,
  input  [7:0]    _EVAL_350,
  input           _EVAL_355,
  input           _EVAL_356,
  input           _EVAL_367,
  input           _EVAL_381,
  input           _EVAL_397,
  input           _EVAL_406,
  input           _EVAL_444,
  input           _EVAL_454,
  input           _EVAL_455,
  input           _EVAL_463,
  input           _EVAL_465,
  input           _EVAL_471,
  input           _EVAL_484,
  input           _EVAL_487,
  input           _EVAL_488,
  input           _EVAL_489,
  input           _EVAL_506,
  input           _EVAL_507,
  input           _EVAL_527,
  input           _EVAL_543,
  input           _EVAL_546,
  input           _EVAL_547,
  input           _EVAL_550,
  input           _EVAL_553,
  input           _EVAL_556,
  input           _EVAL_557,
  input           _EVAL_560,
  input           _EVAL_571,
  input           _EVAL_582,
  input           _EVAL_601,
  input           _EVAL_603,
  input           _EVAL_606,
  input           _EVAL_616,
  input           _EVAL_618,
  input           _EVAL_624,
  input           _EVAL_628,
  input           _EVAL_643,
  input           _EVAL_644,
  input           _EVAL_650,
  input           _EVAL_658,
  input           _EVAL_661,
  input           _EVAL_666,
  input           _EVAL_669,
  input           _EVAL_671,
  input           _EVAL_673,
  input           _EVAL_676,
  input           _EVAL_678,
  input           _EVAL_690,
  input           _EVAL_691,
  input           _EVAL_696,
  input           _EVAL_697,
  input           _EVAL_724,
  input           _EVAL_727,
  input           _EVAL_747,
  input           _EVAL_756,
  input           _EVAL_759,
  input           _EVAL_760,
  input           _EVAL_765,
  input           _EVAL_783,
  input           _EVAL_786,
  input           _EVAL_788,
  input           _EVAL_791,
  input           _EVAL_810,
  input           _EVAL_813,
  input           _EVAL_824,
  input           _EVAL_844,
  input           _EVAL_847,
  input           _EVAL_864,
  input           _EVAL_874,
  input           _EVAL_879,
  input           _EVAL_880,
  input           _EVAL_887,
  input           _EVAL_889,
  input           _EVAL_891,
  input           _EVAL_892,
  input           _EVAL_893,
  input           _EVAL_896,
  input           _EVAL_906,
  input           _EVAL_913,
  input           _EVAL_916,
  input           _EVAL_923,
  input           _EVAL_934,
  input           _EVAL_943,
  input           _EVAL_948,
  input           _EVAL_968,
  input           _EVAL_970,
  input           _EVAL_978,
  input           _EVAL_1005,
  input           _EVAL_1024,
  input           _EVAL_1031,
  input           _EVAL_1040,
  input           _EVAL_1041,
  input           _EVAL_1057,
  input           _EVAL_1059,
  input           _EVAL_1066,
  input           _EVAL_1072,
  input           _EVAL_1073,
  input           _EVAL_1087,
  input           _EVAL_1089,
  input           _EVAL_1093,
  input           _EVAL_1100,
  input           _EVAL_1111,
  input           _EVAL_1117,
  input           _EVAL_1121,
  input           _EVAL_1131,
  input           _EVAL_1147,
  input           _EVAL_1150,
  input  [31:0]   _EVAL_1159,
  input           _EVAL_1163,
  input           _EVAL_1166,
  input           _EVAL_1178,
  input           _EVAL_1187,
  input           _EVAL_1188,
  input           _EVAL_1200,
  input           _EVAL_1206,
  input           _EVAL_1211,
  input           _EVAL_1215,
  input           _EVAL_1225,
  input           _EVAL_1229,
  input           _EVAL_1235,
  input           _EVAL_1240,
  input           _EVAL_1245,
  input           _EVAL_1247,
  input           _EVAL_1250,
  input           _EVAL_1251,
  input           _EVAL_1255,
  input           _EVAL_1261,
  input           _EVAL_1278,
  input           _EVAL_1287,
  input           _EVAL_1293,
  input           _EVAL_1301,
  input           _EVAL_1307,
  input           _EVAL_1311,
  input           _EVAL_1314,
  input           _EVAL_1325,
  input           _EVAL_1331,
  input           _EVAL_1333,
  input           _EVAL_1342,
  input           _EVAL_1352,
  input           _EVAL_1367,
  input           _EVAL_1383,
  input           _EVAL_1388,
  input           _EVAL_1396,
  input           _EVAL_1407,
  input           _EVAL_1408,
  input           _EVAL_1409,
  input           _EVAL_1415,
  input           _EVAL_1444,
  input           _EVAL_1451,
  input           _EVAL_1454,
  input           _EVAL_1462,
  input           _EVAL_1464,
  input           _EVAL_1465,
  input           _EVAL_1493,
  input           _EVAL_1506,
  input           _EVAL_1510,
  input           _EVAL_1524,
  input           _EVAL_1532,
  input           _EVAL_1537,
  input           _EVAL_1544,
  input           _EVAL_1551,
  input           _EVAL_1565,
  input           _EVAL_1575,
  input           _EVAL_1589,
  input           _EVAL_1592,
  input           _EVAL_1593,
  input           _EVAL_1595,
  input           _EVAL_1602,
  input           _EVAL_1618,
  input           _EVAL_1637,
  input           _EVAL_1641,
  input           _EVAL_1645,
  input           _EVAL_1664,
  input           _EVAL_1665,
  input           _EVAL_1666,
  input           _EVAL_1669,
  input           _EVAL_1670,
  input           _EVAL_1671,
  input           _EVAL_1682,
  input           _EVAL_1699,
  input           _EVAL_1706,
  input           _EVAL_1714,
  input           _EVAL_1730,
  input           _EVAL_1762,
  input  [3:0]    _EVAL_1763,
  input           _EVAL_1765,
  input           _EVAL_1777,
  input           _EVAL_1779,
  input           _EVAL_1809,
  input           _EVAL_1820,
  input           _EVAL_1826,
  input           _EVAL_1831,
  input           _EVAL_1834,
  input           _EVAL_1844,
  input           _EVAL_1851,
  input           _EVAL_1864,
  input           _EVAL_1871,
  input           _EVAL_1875,
  input           _EVAL_1877,
  input           _EVAL_1880,
  input           _EVAL_1901,
  input           _EVAL_1907,
  input           _EVAL_1917,
  input           _EVAL_1922,
  input           _EVAL_1929,
  input           _EVAL_1934,
  input           _EVAL_1942,
  input           _EVAL_1949,
  input           _EVAL_1982,
  input           _EVAL_1990,
  input           _EVAL_1999,
  input           _EVAL_2009,
  input           _EVAL_2013,
  input           _EVAL_2020,
  input           _EVAL_2022,
  input           _EVAL_2025,
  input           _EVAL_2052,
  input           _EVAL_2057,
  input           _EVAL_2063,
  input           _EVAL_2065,
  input           _EVAL_2070,
  input           _EVAL_2074,
  input           _EVAL_2077,
  input           _EVAL_2081,
  input           _EVAL_2086,
  input           _EVAL_2091,
  input           _EVAL_2096,
  input           _EVAL_2105,
  input           _EVAL_2108,
  input           _EVAL_2119,
  input           _EVAL_2130,
  input           _EVAL_2141,
  input           _EVAL_2148,
  input           _EVAL_2154,
  input           _EVAL_2160,
  input           _EVAL_2162,
  input           _EVAL_2168,
  input           _EVAL_2176,
  input           _EVAL_2177,
  input           _EVAL_2198,
  input           _EVAL_2202,
  input           _EVAL_2203,
  input           _EVAL_2215,
  input           _EVAL_2216,
  input           _EVAL_2229,
  input           _EVAL_2233,
  input           _EVAL_2239,
  input           _EVAL_2244,
  input           _EVAL_2247,
  input           _EVAL_2249,
  input           _EVAL_2259,
  input           _EVAL_2265,
  input           _EVAL_2277,
  input           _EVAL_2281,
  input           _EVAL_2289,
  input           _EVAL_2291,
  input           _EVAL_2300,
  input           _EVAL_2301,
  input           _EVAL_2308,
  input           _EVAL_2311,
  input           _EVAL_2312,
  input           _EVAL_2324,
  input           _EVAL_2339,
  input           _EVAL_2341,
  input           _EVAL_2343,
  input           _EVAL_2346,
  input           _EVAL_2357,
  input           _EVAL_2360,
  input           _EVAL_2366,
  input           _EVAL_2377,
  input           _EVAL_2381,
  input           _EVAL_2392,
  input           _EVAL_2394,
  input           _EVAL_2400,
  input           _EVAL_2406,
  input           _EVAL_2407,
  input           _EVAL_2413,
  input           _EVAL_2417,
  input           _EVAL_2421,
  input           _EVAL_2422,
  input           _EVAL_2444,
  input           _EVAL_2457,
  input           _EVAL_2484,
  input           _EVAL_2489,
  input           _EVAL_2495,
  input           _EVAL_2499,
  input           _EVAL_2503,
  input           _EVAL_2510,
  input           _EVAL_2515,
  input           _EVAL_2516,
  input           _EVAL_2519,
  input           _EVAL_2520,
  input           _EVAL_2521,
  input           _EVAL_2523,
  input           _EVAL_2528,
  input           _EVAL_2530,
  input           _EVAL_2575,
  input           _EVAL_2577,
  input           _EVAL_2578,
  input           _EVAL_2580,
  input           _EVAL_2583,
  input           _EVAL_2589,
  input           _EVAL_2598,
  input           _EVAL_2605,
  input           _EVAL_2611,
  input           _EVAL_2616,
  input           _EVAL_2622,
  input           _EVAL_2630,
  input           _EVAL_2635,
  input           _EVAL_2660,
  input           _EVAL_2661,
  input           _EVAL_2666,
  input           _EVAL_2668,
  input           _EVAL_2669,
  input           _EVAL_2674,
  input           _EVAL_2690,
  input           _EVAL_2693,
  input           _EVAL_2706,
  input           _EVAL_2711,
  input           _EVAL_2714,
  input           _EVAL_2717,
  input           _EVAL_2737,
  input           _EVAL_2740,
  input           _EVAL_2741,
  input           _EVAL_2755,
  input           _EVAL_2758,
  input           _EVAL_2760,
  input           _EVAL_2766,
  input           _EVAL_2778,
  input           _EVAL_2782,
  input           _EVAL_2804,
  input           _EVAL_2815,
  input           _EVAL_2825,
  input           _EVAL_2828,
  input           _EVAL_2829,
  input           _EVAL_2837,
  input           _EVAL_2841,
  input           _EVAL_2847,
  input           _EVAL_2851,
  input           _EVAL_2861,
  input           _EVAL_2864,
  input           _EVAL_2876,
  input           _EVAL_2884,
  input           _EVAL_2895,
  input           _EVAL_2898,
  input           _EVAL_2905,
  input           _EVAL_2910,
  input           _EVAL_2914,
  input           _EVAL_2915,
  input           _EVAL_2918,
  input           _EVAL_2922,
  input           _EVAL_2929,
  input           _EVAL_2935,
  input           _EVAL_2952,
  input           _EVAL_2988,
  input           _EVAL_2993,
  input           _EVAL_3001,
  input           _EVAL_3030,
  input           _EVAL_3044,
  input  [3:0]    _EVAL_3047,
  input  [7:0]    _EVAL_3048,
  input           _EVAL_3051,
  input           _EVAL_3053,
  input           _EVAL_3056,
  input  [7:0]    _EVAL_3058,
  input           _EVAL_3087,
  input           _EVAL_3094,
  input           _EVAL_3104,
  input           _EVAL_3129,
  input           _EVAL_3133,
  input           _EVAL_3145,
  input           _EVAL_3152,
  input           _EVAL_3154,
  input           _EVAL_3158,
  input           _EVAL_3169,
  input           _EVAL_3171,
  input           _EVAL_3181,
  input           _EVAL_3193,
  input           _EVAL_3194,
  input           _EVAL_3196,
  input           _EVAL_3197,
  input           _EVAL_3200,
  input           _EVAL_3203,
  input           _EVAL_3207,
  input           _EVAL_3211,
  input           _EVAL_3213,
  input           _EVAL_3225,
  input           _EVAL_3230,
  input           _EVAL_3234,
  input           _EVAL_3266,
  input           _EVAL_3280,
  input           _EVAL_3285,
  input           _EVAL_3286,
  input           _EVAL_3290,
  input           _EVAL_3294,
  input           _EVAL_3298,
  input           _EVAL_3311,
  input           _EVAL_3327,
  input           _EVAL_3336,
  input           _EVAL_3345,
  input           _EVAL_3358,
  input           _EVAL_3363,
  input           _EVAL_3365,
  input           _EVAL_3374,
  input           _EVAL_3389,
  input           _EVAL_3390,
  input           _EVAL_3391,
  input           _EVAL_3410,
  input           _EVAL_3422,
  input  [3:0]    _EVAL_3427,
  input           _EVAL_3434,
  input           _EVAL_3435,
  input           _EVAL_3438,
  input           _EVAL_3439,
  input           _EVAL_3441,
  input           _EVAL_3443,
  input           _EVAL_3450,
  input           _EVAL_3456,
  input           _EVAL_3466,
  input           _EVAL_3472,
  input           _EVAL_3475,
  input           _EVAL_3479,
  input           _EVAL_3487,
  input           _EVAL_3493,
  input           _EVAL_3501,
  input           _EVAL_3502,
  input           _EVAL_3516,
  input           _EVAL_3517,
  input           _EVAL_3530,
  input           _EVAL_3535,
  input           _EVAL_3537,
  input           _EVAL_3542,
  input           _EVAL_3561,
  input           _EVAL_3564,
  input           _EVAL_3580,
  input           _EVAL_3584,
  input           _EVAL_3589,
  input           _EVAL_3590,
  input           _EVAL_3594,
  input           _EVAL_3603,
  input           _EVAL_3607,
  input           _EVAL_3609,
  input           _EVAL_3613,
  input           _EVAL_3620,
  input           _EVAL_3629,
  input           _EVAL_3634,
  input           _EVAL_3636,
  input           _EVAL_3639,
  input           _EVAL_3641,
  input           _EVAL_3642,
  input           _EVAL_3644,
  input           _EVAL_3646,
  input           _EVAL_3652,
  input           _EVAL_3683,
  input           _EVAL_3705,
  input           _EVAL_3716,
  input           _EVAL_3735,
  input           _EVAL_3737,
  input           _EVAL_3739,
  input           _EVAL_3748,
  input           _EVAL_3753,
  input           _EVAL_3757,
  input           _EVAL_3758,
  input           _EVAL_3783,
  input           _EVAL_3789,
  input           _EVAL_3795,
  input           _EVAL_3799,
  input           _EVAL_3805,
  input           _EVAL_3831,
  input           _EVAL_3843,
  input           _EVAL_3847,
  input           _EVAL_3854,
  input           _EVAL_3861,
  input           _EVAL_3866,
  input           _EVAL_3876,
  input           _EVAL_3887,
  input           _EVAL_3892,
  input           _EVAL_3899,
  input           _EVAL_3911,
  input           _EVAL_3914,
  input           _EVAL_3922,
  input           _EVAL_3939,
  input           _EVAL_3940,
  input           _EVAL_3944,
  input  [3:0]    _EVAL_3945,
  input           _EVAL_3946,
  input           _EVAL_3958,
  input           _EVAL_3962,
  input           _EVAL_3965,
  input           _EVAL_3967,
  input           _EVAL_3977,
  input           _EVAL_3980,
  input           _EVAL_3983,
  input           _EVAL_3985,
  input           _EVAL_3986,
  input           _EVAL_3999,
  input           _EVAL_4005,
  input           _EVAL_4007,
  input           _EVAL_4008,
  input           _EVAL_4013,
  input           _EVAL_4014,
  input           _EVAL_4025,
  input           _EVAL_4045,
  input           _EVAL_4051,
  input           _EVAL_4053,
  input           _EVAL_4065,
  input           _EVAL_4068,
  input           _EVAL_4080,
  input           _EVAL_4085,
  input           _EVAL_4087,
  input           _EVAL_4096,
  input           _EVAL_4103,
  input           _EVAL_4115,
  input           _EVAL_4117,
  input           _EVAL_4119,
  input           _EVAL_4162,
  input           _EVAL_4164,
  input           _EVAL_4167,
  input           _EVAL_4168,
  input           _EVAL_4174,
  input           _EVAL_4184,
  input  [3:0]    _EVAL_4213,
  input           _EVAL_4233,
  input           _EVAL_4236,
  input           _EVAL_4242,
  input           _EVAL_4246,
  input           _EVAL_4255,
  input           _EVAL_4271,
  input           _EVAL_4282,
  input           _EVAL_4291,
  input           _EVAL_4297,
  input           _EVAL_4301,
  input           _EVAL_4308,
  input           _EVAL_4336,
  input           _EVAL_4338,
  input           _EVAL_4339,
  input           _EVAL_4344,
  input           _EVAL_4348,
  input           _EVAL_4367,
  input           _EVAL_4374,
  input           _EVAL_4382,
  input           _EVAL_4386,
  input           _EVAL_4397,
  input           _EVAL_4398,
  input           _EVAL_4403,
  input           _EVAL_4406,
  input           _EVAL_4414,
  input           _EVAL_4437,
  input           _EVAL_4440,
  input           _EVAL_4441,
  input           _EVAL_4443,
  input           _EVAL_4449,
  input           _EVAL_4467,
  input           _EVAL_4476,
  input           _EVAL_4477,
  input           _EVAL_4480,
  input           _EVAL_4500,
  input           _EVAL_4532,
  input           _EVAL_4547,
  input           _EVAL_4554,
  input           _EVAL_4566,
  input           _EVAL_4584,
  input           _EVAL_4588,
  input           _EVAL_4599,
  input           _EVAL_4610,
  input           _EVAL_4612,
  input           _EVAL_4620,
  input           _EVAL_4650,
  input           _EVAL_4662,
  input           _EVAL_4676,
  input           _EVAL_4684,
  input           _EVAL_4696,
  input           _EVAL_4732,
  input           _EVAL_4738,
  input           _EVAL_4742,
  input           _EVAL_4753,
  input           _EVAL_4779,
  input           _EVAL_4785,
  input           _EVAL_4791,
  input           _EVAL_4797,
  input           _EVAL_4807,
  input           _EVAL_4808,
  input           _EVAL_4810,
  input           _EVAL_4815,
  input           _EVAL_4819,
  input           _EVAL_4822,
  input           _EVAL_4839,
  input           _EVAL_4843,
  input           _EVAL_4876,
  input           _EVAL_4878,
  input           _EVAL_4882,
  input           _EVAL_4901,
  input           _EVAL_4922,
  input           _EVAL_4932,
  input           _EVAL_4937,
  input           _EVAL_4942,
  input           _EVAL_4944,
  input           _EVAL_4955,
  input           _EVAL_4956,
  input           _EVAL_4959,
  input           _EVAL_4965,
  input           _EVAL_4968,
  input  [23:0]   _EVAL_4986,
  input           _EVAL_4992,
  input  [7:0]    _EVAL_5000,
  input           _EVAL_5002,
  input           _EVAL_5012,
  input           _EVAL_5014,
  input           _EVAL_5022,
  input           _EVAL_5024,
  input           _EVAL_5029,
  input           _EVAL_5030,
  input           _EVAL_5034,
  input           _EVAL_5041,
  input           _EVAL_5046,
  input  [1023:0] _EVAL_5068,
  input           _EVAL_5086,
  input           _EVAL_5101,
  input           _EVAL_5108,
  input           _EVAL_5111,
  input           _EVAL_5115,
  input           _EVAL_5131,
  input           _EVAL_5147,
  input           _EVAL_5150,
  input           _EVAL_5154,
  input           _EVAL_5163,
  input           _EVAL_5168,
  input           _EVAL_5169,
  input           _EVAL_5172,
  input           _EVAL_5188,
  input           _EVAL_5190,
  input           _EVAL_5195,
  input           _EVAL_5203,
  input           _EVAL_5221,
  input           _EVAL_5225,
  input           _EVAL_5232,
  input           _EVAL_5249,
  input           _EVAL_5255,
  input           _EVAL_5266,
  input           _EVAL_5267,
  input           _EVAL_5269,
  input           _EVAL_5288,
  input           _EVAL_5293,
  input           _EVAL_5294,
  input           _EVAL_5300,
  input           _EVAL_5307,
  input           _EVAL_5309,
  input           _EVAL_5315,
  input           _EVAL_5326,
  input           _EVAL_5331,
  input           _EVAL_5340,
  input           _EVAL_5345,
  input           _EVAL_5348,
  input           _EVAL_5350,
  input           _EVAL_5363,
  input           _EVAL_5369,
  input           _EVAL_5386,
  input           _EVAL_5390,
  input           _EVAL_5391,
  input           _EVAL_5405,
  input           _EVAL_5409,
  input           _EVAL_5411,
  input           _EVAL_5421,
  input           _EVAL_5448,
  input           _EVAL_5469,
  input           _EVAL_5479,
  input           _EVAL_5481,
  input           _EVAL_5484,
  input           _EVAL_5491,
  input           _EVAL_5506,
  input           _EVAL_5516,
  input           _EVAL_5521,
  input           _EVAL_5535,
  input           _EVAL_5539,
  input           _EVAL_5546,
  input           _EVAL_5556,
  input           _EVAL_5557,
  input           _EVAL_5558,
  input           _EVAL_5582,
  input           _EVAL_5591,
  input           _EVAL_5597,
  input           _EVAL_5600,
  input           _EVAL_5603,
  input           _EVAL_5608,
  input           _EVAL_5609,
  input           _EVAL_5619,
  input           _EVAL_5627,
  input           _EVAL_5629,
  input           _EVAL_5637,
  input           _EVAL_5646,
  input           _EVAL_5657,
  input           _EVAL_5682,
  input           _EVAL_5684,
  input           _EVAL_5696,
  input           _EVAL_5699,
  input           _EVAL_5711,
  input           _EVAL_5730,
  input           _EVAL_5735,
  input           _EVAL_5741,
  input           _EVAL_5743,
  input           _EVAL_5745,
  input           _EVAL_5748,
  input           _EVAL_5759,
  input           _EVAL_5771,
  input           _EVAL_5781,
  input           _EVAL_5782,
  input           _EVAL_5800,
  input           _EVAL_5802,
  input           _EVAL_5813,
  input           _EVAL_5818,
  input           _EVAL_5829,
  input           _EVAL_5833,
  input           _EVAL_5841,
  input           _EVAL_5846,
  input           _EVAL_5851,
  input           _EVAL_5860,
  input           _EVAL_5862,
  input           _EVAL_5878,
  input           _EVAL_5890,
  input           _EVAL_5894,
  input  [3:0]    _EVAL_5905,
  input           _EVAL_5907,
  input           _EVAL_5909,
  input  [3:0]    _EVAL_5913,
  input           _EVAL_5916,
  input           _EVAL_5924,
  input           _EVAL_5940,
  input           _EVAL_5957,
  input           _EVAL_5966,
  input           _EVAL_5984,
  input           _EVAL_5985,
  input           _EVAL_5993,
  input           _EVAL_5997,
  input           _EVAL_6004,
  input           _EVAL_6009,
  input           _EVAL_6014,
  input           _EVAL_6021,
  input           _EVAL_6023,
  input           _EVAL_6030,
  input           _EVAL_6042,
  input           _EVAL_6043,
  input           _EVAL_6046,
  input           _EVAL_6060,
  input           _EVAL_6071,
  input           _EVAL_6074,
  input           _EVAL_6081,
  input           _EVAL_6092,
  input           _EVAL_6098,
  input           _EVAL_6101,
  input  [1:0]    Queue__EVAL_11,
  input  [2:0]    Queue__EVAL_0,
  input           Queue__EVAL_9,
  input           Queue__EVAL_14,
  input           Queue__EVAL_2
);
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_157;
  wire  _EVAL_159;
  wire  _EVAL_162;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_175;
  wire  _EVAL_177;
  wire  _EVAL_179;
  wire  _EVAL_181;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_187;
  wire  _EVAL_191;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_196;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_231;
  wire  _EVAL_233;
  wire  _EVAL_235;
  wire  _EVAL_237;
  wire  _EVAL_239;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_271;
  wire  _EVAL_275;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_282;
  wire  _EVAL_284;
  wire  _EVAL_287;
  wire  _EVAL_290;
  wire  _EVAL_292;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_307;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_314;
  wire  _EVAL_316;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_321;
  wire  _EVAL_322;
  wire [3:0] _EVAL_323;
  wire  _EVAL_326;
  wire  _EVAL_327;
  wire  _EVAL_328;
  wire  _EVAL_330;
  wire  _EVAL_331;
  wire  _EVAL_332;
  wire [7:0] _EVAL_334;
  wire  _EVAL_335;
  wire  _EVAL_339;
  wire  _EVAL_341;
  wire  _EVAL_342;
  wire  _EVAL_345;
  wire  _EVAL_346;
  wire  _EVAL_347;
  wire  _EVAL_348;
  wire  _EVAL_351;
  wire  _EVAL_352;
  wire  _EVAL_354;
  wire  _EVAL_357;
  wire  _EVAL_358;
  wire  _EVAL_360;
  wire  _EVAL_361;
  wire  _EVAL_362;
  wire  _EVAL_363;
  wire  _EVAL_364;
  wire  _EVAL_365;
  wire  _EVAL_369;
  wire  _EVAL_370;
  wire  _EVAL_372;
  wire  _EVAL_373;
  wire  _EVAL_374;
  wire  _EVAL_375;
  wire  _EVAL_376;
  wire  _EVAL_377;
  wire  _EVAL_378;
  wire  _EVAL_380;
  wire [1:0] _EVAL_383;
  wire  _EVAL_385;
  wire  _EVAL_386;
  wire  _EVAL_387;
  wire  _EVAL_388;
  wire  _EVAL_389;
  wire  _EVAL_390;
  wire  _EVAL_391;
  wire  _EVAL_392;
  wire  _EVAL_395;
  wire  _EVAL_396;
  wire  _EVAL_398;
  wire  _EVAL_402;
  wire  _EVAL_407;
  wire [6:0] _EVAL_408;
  wire  _EVAL_409;
  wire  _EVAL_410;
  wire  _EVAL_413;
  wire  _EVAL_415;
  wire  _EVAL_418;
  wire  _EVAL_421;
  wire  _EVAL_422;
  wire  _EVAL_424;
  wire  _EVAL_428;
  wire  _EVAL_429;
  wire  _EVAL_434;
  wire  _EVAL_435;
  wire  _EVAL_440;
  wire  _EVAL_441;
  wire  _EVAL_442;
  wire  _EVAL_446;
  wire  _EVAL_449;
  wire  _EVAL_451;
  wire  _EVAL_453;
  wire  _EVAL_457;
  wire  _EVAL_458;
  wire  _EVAL_460;
  wire  _EVAL_461;
  wire  _EVAL_462;
  wire  _EVAL_464;
  wire  _EVAL_467;
  wire  _EVAL_469;
  wire  _EVAL_470;
  wire  _EVAL_473;
  wire  _EVAL_474;
  wire  _EVAL_475;
  wire  _EVAL_476;
  wire  _EVAL_477;
  wire  _EVAL_478;
  wire  _EVAL_479;
  wire  _EVAL_480;
  wire  _EVAL_481;
  wire  _EVAL_482;
  wire  _EVAL_486;
  wire  _EVAL_490;
  wire  _EVAL_491;
  wire  _EVAL_492;
  wire  _EVAL_496;
  wire  _EVAL_503;
  wire  _EVAL_504;
  wire  _EVAL_508;
  wire  _EVAL_509;
  wire  _EVAL_510;
  wire  _EVAL_512;
  wire  _EVAL_513;
  wire  _EVAL_515;
  wire  _EVAL_521;
  wire [7:0] _EVAL_523;
  wire  _EVAL_528;
  wire  _EVAL_529;
  wire  _EVAL_530;
  wire  _EVAL_532;
  wire  _EVAL_534;
  wire  _EVAL_535;
  wire  _EVAL_536;
  wire  _EVAL_537;
  wire  _EVAL_538;
  wire  _EVAL_539;
  wire  _EVAL_540;
  wire  _EVAL_541;
  wire  _EVAL_544;
  wire  _EVAL_549;
  wire  _EVAL_551;
  wire  _EVAL_552;
  wire  _EVAL_554;
  wire  _EVAL_555;
  wire  _EVAL_562;
  wire  _EVAL_564;
  wire  _EVAL_565;
  wire  _EVAL_566;
  wire [3:0] _EVAL_568;
  wire  _EVAL_570;
  wire  _EVAL_572;
  wire  _EVAL_573;
  wire  _EVAL_574;
  wire  _EVAL_577;
  wire  _EVAL_578;
  wire  _EVAL_579;
  wire  _EVAL_580;
  wire  _EVAL_581;
  wire  _EVAL_583;
  wire  _EVAL_584;
  wire  _EVAL_585;
  wire  _EVAL_586;
  wire  _EVAL_587;
  wire  _EVAL_588;
  wire  _EVAL_589;
  wire  _EVAL_590;
  wire  _EVAL_591;
  wire  _EVAL_594;
  wire  _EVAL_596;
  wire  _EVAL_599;
  wire  _EVAL_600;
  wire  _EVAL_608;
  wire  _EVAL_610;
  wire  _EVAL_612;
  wire  _EVAL_613;
  wire  _EVAL_617;
  wire  _EVAL_619;
  wire  _EVAL_620;
  wire  _EVAL_621;
  wire  _EVAL_622;
  wire  _EVAL_623;
  wire  _EVAL_625;
  wire  _EVAL_626;
  wire  _EVAL_627;
  wire  _EVAL_629;
  wire  _EVAL_630;
  wire  _EVAL_631;
  wire  _EVAL_633;
  wire  _EVAL_635;
  wire  _EVAL_637;
  wire  _EVAL_638;
  wire  _EVAL_641;
  wire  _EVAL_645;
  wire  _EVAL_646;
  wire  _EVAL_649;
  wire  _EVAL_651;
  wire  _EVAL_652;
  wire  _EVAL_654;
  wire  _EVAL_656;
  wire  _EVAL_659;
  wire  _EVAL_660;
  wire  _EVAL_663;
  wire  _EVAL_668;
  wire  _EVAL_670;
  wire  _EVAL_679;
  wire  _EVAL_680;
  wire  _EVAL_682;
  wire  _EVAL_684;
  wire  _EVAL_686;
  wire  _EVAL_688;
  wire  _EVAL_692;
  wire  _EVAL_694;
  wire  _EVAL_695;
  wire  _EVAL_698;
  wire  _EVAL_699;
  wire  _EVAL_701;
  wire  _EVAL_704;
  wire  _EVAL_708;
  wire [6:0] _EVAL_709;
  wire  _EVAL_710;
  wire  _EVAL_711;
  wire  _EVAL_712;
  wire  _EVAL_713;
  wire  _EVAL_714;
  wire  _EVAL_721;
  wire  _EVAL_722;
  wire  _EVAL_725;
  wire  _EVAL_726;
  wire  _EVAL_731;
  wire  _EVAL_734;
  wire  _EVAL_735;
  wire  _EVAL_739;
  wire  _EVAL_740;
  wire  _EVAL_744;
  wire  _EVAL_745;
  wire  _EVAL_746;
  wire  _EVAL_748;
  wire  _EVAL_751;
  wire  _EVAL_752;
  wire  _EVAL_754;
  wire  _EVAL_755;
  wire  _EVAL_757;
  wire  _EVAL_758;
  wire  _EVAL_761;
  wire  _EVAL_764;
  wire  _EVAL_767;
  wire  _EVAL_768;
  wire  _EVAL_769;
  wire  _EVAL_770;
  wire  _EVAL_771;
  wire  _EVAL_773;
  wire  _EVAL_774;
  wire  _EVAL_775;
  wire  _EVAL_776;
  wire  _EVAL_777;
  wire  _EVAL_778;
  wire  _EVAL_779;
  wire  _EVAL_781;
  wire  _EVAL_787;
  wire  _EVAL_789;
  wire  _EVAL_790;
  wire  _EVAL_792;
  wire  _EVAL_793;
  wire  _EVAL_797;
  wire  _EVAL_798;
  wire  _EVAL_799;
  wire  _EVAL_800;
  wire  _EVAL_801;
  wire  _EVAL_802;
  wire  _EVAL_803;
  wire  _EVAL_804;
  wire  _EVAL_807;
  wire  _EVAL_808;
  wire  _EVAL_809;
  wire  _EVAL_814;
  wire  _EVAL_816;
  wire  _EVAL_817;
  wire  _EVAL_818;
  wire  _EVAL_819;
  wire  _EVAL_820;
  wire  _EVAL_821;
  wire  _EVAL_825;
  wire  _EVAL_826;
  wire  _EVAL_827;
  wire  _EVAL_828;
  wire  _EVAL_829;
  wire  _EVAL_830;
  wire  _EVAL_831;
  wire  _EVAL_832;
  wire  _EVAL_836;
  wire  _EVAL_837;
  wire  _EVAL_839;
  wire  _EVAL_842;
  wire  _EVAL_843;
  wire  _EVAL_845;
  wire  _EVAL_849;
  wire  _EVAL_854;
  wire  _EVAL_856;
  wire  _EVAL_857;
  wire  _EVAL_859;
  wire  _EVAL_860;
  wire  _EVAL_862;
  wire  _EVAL_865;
  wire  _EVAL_867;
  wire  _EVAL_868;
  wire  _EVAL_869;
  wire  _EVAL_870;
  wire  _EVAL_871;
  wire  _EVAL_873;
  wire  _EVAL_875;
  wire  _EVAL_876;
  wire  _EVAL_877;
  wire  _EVAL_878;
  wire  _EVAL_882;
  wire  _EVAL_884;
  wire  _EVAL_885;
  wire  _EVAL_886;
  wire  _EVAL_888;
  wire  _EVAL_894;
  wire  _EVAL_895;
  wire  _EVAL_897;
  wire  _EVAL_900;
  wire  _EVAL_904;
  wire  _EVAL_905;
  wire  _EVAL_908;
  wire  _EVAL_909;
  wire  _EVAL_910;
  wire  _EVAL_911;
  wire  _EVAL_914;
  wire  _EVAL_917;
  wire  _EVAL_920;
  wire  _EVAL_921;
  wire  _EVAL_922;
  wire  _EVAL_925;
  wire  _EVAL_926;
  wire  _EVAL_927;
  wire  _EVAL_928;
  wire  _EVAL_931;
  wire  _EVAL_932;
  wire  _EVAL_933;
  wire  _EVAL_935;
  wire  _EVAL_936;
  wire  _EVAL_937;
  wire  _EVAL_938;
  wire  _EVAL_940;
  wire  _EVAL_941;
  wire  _EVAL_944;
  wire  _EVAL_946;
  wire  _EVAL_947;
  wire  _EVAL_949;
  wire  _EVAL_950;
  wire  _EVAL_951;
  wire  _EVAL_952;
  wire  _EVAL_954;
  wire  _EVAL_955;
  wire  _EVAL_956;
  wire  _EVAL_957;
  wire  _EVAL_961;
  wire  _EVAL_963;
  wire  _EVAL_964;
  wire  _EVAL_965;
  wire  _EVAL_967;
  wire  _EVAL_971;
  wire  _EVAL_972;
  wire  _EVAL_973;
  wire  _EVAL_974;
  wire  _EVAL_975;
  wire  _EVAL_976;
  wire  _EVAL_982;
  wire  _EVAL_983;
  wire  _EVAL_984;
  wire  _EVAL_985;
  wire  _EVAL_987;
  wire  _EVAL_989;
  wire  _EVAL_996;
  wire  _EVAL_997;
  wire  _EVAL_998;
  wire  _EVAL_1000;
  wire  _EVAL_1001;
  wire  _EVAL_1003;
  wire  _EVAL_1004;
  wire  _EVAL_1006;
  wire  _EVAL_1007;
  wire  _EVAL_1008;
  wire  _EVAL_1009;
  wire  _EVAL_1010;
  wire  _EVAL_1012;
  wire  _EVAL_1014;
  wire  _EVAL_1015;
  wire  _EVAL_1016;
  wire  _EVAL_1017;
  wire  _EVAL_1019;
  wire  _EVAL_1022;
  wire  _EVAL_1025;
  wire  _EVAL_1029;
  wire  _EVAL_1033;
  wire  _EVAL_1034;
  wire  _EVAL_1036;
  wire  _EVAL_1037;
  wire  _EVAL_1038;
  wire  _EVAL_1039;
  wire  _EVAL_1043;
  wire  _EVAL_1044;
  wire  _EVAL_1045;
  wire  _EVAL_1046;
  wire  _EVAL_1047;
  wire  _EVAL_1049;
  wire  _EVAL_1050;
  wire  _EVAL_1051;
  wire  _EVAL_1053;
  wire  _EVAL_1055;
  wire  _EVAL_1058;
  wire  _EVAL_1061;
  wire  _EVAL_1062;
  wire  _EVAL_1063;
  wire  _EVAL_1064;
  wire  _EVAL_1065;
  wire  _EVAL_1067;
  wire  _EVAL_1068;
  wire  _EVAL_1069;
  wire  _EVAL_1070;
  wire  _EVAL_1071;
  wire  _EVAL_1076;
  wire  _EVAL_1077;
  wire  _EVAL_1078;
  wire  _EVAL_1079;
  wire  _EVAL_1081;
  wire  _EVAL_1082;
  wire  _EVAL_1083;
  wire  _EVAL_1084;
  wire  _EVAL_1085;
  wire  _EVAL_1086;
  wire  _EVAL_1088;
  wire  _EVAL_1090;
  wire  _EVAL_1094;
  wire  _EVAL_1095;
  wire  _EVAL_1096;
  wire  _EVAL_1097;
  wire  _EVAL_1099;
  wire  _EVAL_1102;
  wire  _EVAL_1103;
  wire  _EVAL_1104;
  wire  _EVAL_1105;
  wire  _EVAL_1107;
  wire  _EVAL_1108;
  wire  _EVAL_1109;
  wire  _EVAL_1116;
  wire  _EVAL_1118;
  wire  _EVAL_1122;
  wire  _EVAL_1125;
  wire  _EVAL_1126;
  wire  _EVAL_1127;
  wire  _EVAL_1133;
  wire  _EVAL_1134;
  wire  _EVAL_1136;
  wire  _EVAL_1137;
  wire  _EVAL_1139;
  wire  _EVAL_1142;
  wire  _EVAL_1144;
  wire [1023:0] _EVAL_1145;
  wire  _EVAL_1146;
  wire  _EVAL_1149;
  wire  _EVAL_1151;
  wire  _EVAL_1152;
  wire  _EVAL_1155;
  wire  _EVAL_1158;
  wire  _EVAL_1161;
  wire  _EVAL_1162;
  wire  _EVAL_1165;
  wire  _EVAL_1167;
  wire  _EVAL_1169;
  wire  _EVAL_1170;
  wire  _EVAL_1171;
  wire  _EVAL_1173;
  wire  _EVAL_1175;
  wire  _EVAL_1176;
  wire  _EVAL_1179;
  wire  _EVAL_1180;
  wire  _EVAL_1182;
  wire  _EVAL_1183;
  wire  _EVAL_1185;
  wire  _EVAL_1189;
  wire  _EVAL_1193;
  wire  _EVAL_1194;
  wire  _EVAL_1195;
  wire  _EVAL_1196;
  wire  _EVAL_1197;
  wire  _EVAL_1198;
  wire  _EVAL_1199;
  wire  _EVAL_1201;
  wire  _EVAL_1202;
  wire  _EVAL_1203;
  wire  _EVAL_1207;
  wire  _EVAL_1209;
  wire  _EVAL_1210;
  wire  _EVAL_1212;
  wire  _EVAL_1213;
  wire  _EVAL_1214;
  wire  _EVAL_1223;
  wire  _EVAL_1224;
  wire  _EVAL_1226;
  wire  _EVAL_1227;
  wire  _EVAL_1231;
  wire  _EVAL_1233;
  wire  _EVAL_1234;
  wire  _EVAL_1241;
  wire  _EVAL_1242;
  wire  _EVAL_1243;
  wire  _EVAL_1244;
  wire  _EVAL_1246;
  wire  _EVAL_1254;
  wire  _EVAL_1256;
  wire  _EVAL_1259;
  wire  _EVAL_1262;
  wire  _EVAL_1266;
  wire  _EVAL_1268;
  wire  _EVAL_1269;
  wire  _EVAL_1270;
  wire  _EVAL_1272;
  wire  _EVAL_1274;
  wire  _EVAL_1277;
  wire  _EVAL_1281;
  wire  _EVAL_1283;
  wire  _EVAL_1285;
  wire  _EVAL_1290;
  wire  _EVAL_1291;
  wire  _EVAL_1294;
  wire  _EVAL_1296;
  wire  _EVAL_1297;
  wire  _EVAL_1299;
  wire  _EVAL_1300;
  wire  _EVAL_1302;
  wire  _EVAL_1305;
  wire  _EVAL_1310;
  wire  _EVAL_1312;
  wire  _EVAL_1313;
  wire [31:0] _EVAL_1316;
  wire  _EVAL_1317;
  wire  _EVAL_1319;
  wire  _EVAL_1322;
  wire  _EVAL_1324;
  wire  _EVAL_1326;
  wire  _EVAL_1327;
  wire  _EVAL_1328;
  wire  _EVAL_1329;
  wire  _EVAL_1332;
  wire  _EVAL_1334;
  wire  _EVAL_1338;
  wire  _EVAL_1340;
  wire  _EVAL_1341;
  wire  _EVAL_1343;
  wire  _EVAL_1344;
  wire  _EVAL_1346;
  wire  _EVAL_1348;
  wire  _EVAL_1349;
  wire  _EVAL_1350;
  wire  _EVAL_1355;
  wire  _EVAL_1358;
  wire  _EVAL_1360;
  wire  _EVAL_1361;
  wire  _EVAL_1363;
  wire  _EVAL_1364;
  wire  _EVAL_1365;
  wire  _EVAL_1366;
  wire  _EVAL_1369;
  wire  _EVAL_1370;
  wire  _EVAL_1371;
  wire  _EVAL_1373;
  wire  _EVAL_1375;
  wire  _EVAL_1376;
  wire  _EVAL_1380;
  wire  _EVAL_1384;
  wire  _EVAL_1385;
  wire  _EVAL_1386;
  wire  _EVAL_1387;
  wire  _EVAL_1389;
  wire  _EVAL_1391;
  wire  _EVAL_1392;
  wire  _EVAL_1393;
  wire  _EVAL_1394;
  wire  _EVAL_1395;
  wire  _EVAL_1399;
  wire  _EVAL_1401;
  wire  _EVAL_1402;
  wire  _EVAL_1404;
  wire  _EVAL_1405;
  wire  _EVAL_1406;
  wire  _EVAL_1411;
  wire  _EVAL_1412;
  wire  _EVAL_1413;
  wire  _EVAL_1418;
  wire  _EVAL_1419;
  wire  _EVAL_1420;
  wire  _EVAL_1421;
  wire  _EVAL_1424;
  wire  _EVAL_1426;
  wire  _EVAL_1428;
  wire  _EVAL_1432;
  wire  _EVAL_1434;
  wire  _EVAL_1439;
  wire  _EVAL_1443;
  wire  _EVAL_1446;
  wire  _EVAL_1447;
  wire  _EVAL_1448;
  wire  _EVAL_1449;
  wire  _EVAL_1450;
  wire  _EVAL_1452;
  wire  _EVAL_1453;
  wire  _EVAL_1455;
  wire  _EVAL_1458;
  wire  _EVAL_1459;
  wire  _EVAL_1463;
  wire  _EVAL_1467;
  wire  _EVAL_1468;
  wire [3:0] _EVAL_1470;
  wire  _EVAL_1471;
  wire [7:0] _EVAL_1475;
  wire  _EVAL_1478;
  wire  _EVAL_1479;
  wire  _EVAL_1480;
  wire  _EVAL_1482;
  wire  _EVAL_1483;
  wire  _EVAL_1485;
  wire  _EVAL_1487;
  wire  _EVAL_1488;
  wire  _EVAL_1489;
  wire  _EVAL_1490;
  wire  _EVAL_1491;
  wire  _EVAL_1494;
  wire  _EVAL_1499;
  wire  _EVAL_1500;
  wire  _EVAL_1501;
  wire  _EVAL_1505;
  wire  _EVAL_1509;
  wire  _EVAL_1511;
  wire  _EVAL_1512;
  wire  _EVAL_1513;
  wire  _EVAL_1514;
  wire  _EVAL_1516;
  wire  _EVAL_1518;
  wire  _EVAL_1521;
  wire  _EVAL_1523;
  wire  _EVAL_1525;
  wire  _EVAL_1526;
  wire  _EVAL_1528;
  wire  _EVAL_1529;
  wire  _EVAL_1530;
  wire  _EVAL_1533;
  wire  _EVAL_1535;
  wire  _EVAL_1536;
  wire  _EVAL_1538;
  wire  _EVAL_1539;
  wire  _EVAL_1541;
  wire  _EVAL_1542;
  wire  _EVAL_1543;
  wire  _EVAL_1545;
  wire  _EVAL_1546;
  wire  _EVAL_1547;
  wire  _EVAL_1548;
  wire  _EVAL_1553;
  wire  _EVAL_1555;
  wire  _EVAL_1557;
  wire  _EVAL_1558;
  wire  _EVAL_1559;
  wire  _EVAL_1561;
  wire  _EVAL_1562;
  wire  _EVAL_1563;
  wire  _EVAL_1567;
  wire  _EVAL_1568;
  wire  _EVAL_1570;
  wire  _EVAL_1574;
  wire  _EVAL_1578;
  wire  _EVAL_1579;
  wire  _EVAL_1580;
  wire  _EVAL_1582;
  wire  _EVAL_1584;
  wire  _EVAL_1585;
  wire  _EVAL_1586;
  wire  _EVAL_1588;
  wire  _EVAL_1590;
  wire  _EVAL_1591;
  wire  _EVAL_1594;
  wire  _EVAL_1596;
  wire  _EVAL_1599;
  wire  _EVAL_1600;
  wire  _EVAL_1601;
  wire  _EVAL_1603;
  wire  _EVAL_1604;
  wire  _EVAL_1605;
  wire  _EVAL_1606;
  wire  _EVAL_1607;
  wire  _EVAL_1611;
  wire  _EVAL_1612;
  wire  _EVAL_1615;
  wire  _EVAL_1616;
  wire [6:0] _EVAL_1619;
  wire  _EVAL_1620;
  wire  _EVAL_1622;
  wire  _EVAL_1624;
  wire  _EVAL_1625;
  wire  _EVAL_1627;
  wire  _EVAL_1628;
  wire  _EVAL_1631;
  wire  _EVAL_1633;
  wire  _EVAL_1634;
  wire  _EVAL_1635;
  wire  _EVAL_1638;
  wire  _EVAL_1639;
  wire  _EVAL_1640;
  wire  _EVAL_1642;
  wire  _EVAL_1647;
  wire  _EVAL_1649;
  wire  _EVAL_1650;
  wire  _EVAL_1651;
  wire  _EVAL_1652;
  wire  _EVAL_1653;
  wire  _EVAL_1655;
  wire  _EVAL_1657;
  wire  _EVAL_1658;
  wire  _EVAL_1660;
  wire  _EVAL_1661;
  wire  _EVAL_1663;
  wire  _EVAL_1667;
  wire  _EVAL_1673;
  wire  _EVAL_1675;
  wire  _EVAL_1677;
  wire  _EVAL_1679;
  wire  _EVAL_1684;
  wire  _EVAL_1685;
  wire  _EVAL_1687;
  wire  _EVAL_1689;
  wire  _EVAL_1691;
  wire  _EVAL_1692;
  wire  _EVAL_1694;
  wire  _EVAL_1695;
  wire  _EVAL_1696;
  wire  _EVAL_1697;
  wire  _EVAL_1700;
  wire  _EVAL_1701;
  wire  _EVAL_1702;
  wire  _EVAL_1703;
  wire  _EVAL_1707;
  wire  _EVAL_1708;
  wire  _EVAL_1709;
  wire  _EVAL_1711;
  wire  _EVAL_1715;
  wire  _EVAL_1716;
  wire  _EVAL_1717;
  wire  _EVAL_1718;
  wire  _EVAL_1719;
  wire  _EVAL_1721;
  wire  _EVAL_1722;
  wire  _EVAL_1723;
  wire  _EVAL_1724;
  wire  _EVAL_1725;
  wire  _EVAL_1727;
  wire  _EVAL_1728;
  wire  _EVAL_1729;
  wire [1:0] _EVAL_1731;
  wire  _EVAL_1733;
  wire  _EVAL_1734;
  wire  _EVAL_1735;
  wire  _EVAL_1736;
  wire  _EVAL_1739;
  wire  _EVAL_1741;
  wire  _EVAL_1742;
  wire  _EVAL_1743;
  wire  _EVAL_1745;
  wire  _EVAL_1747;
  wire  _EVAL_1750;
  wire  _EVAL_1752;
  wire  _EVAL_1754;
  wire  _EVAL_1755;
  wire  _EVAL_1756;
  wire  _EVAL_1757;
  wire  _EVAL_1764;
  wire  _EVAL_1767;
  wire  _EVAL_1769;
  wire  _EVAL_1772;
  wire  _EVAL_1773;
  wire  _EVAL_1774;
  wire  _EVAL_1776;
  wire  _EVAL_1778;
  wire  _EVAL_1781;
  wire  _EVAL_1782;
  wire  _EVAL_1783;
  wire  _EVAL_1784;
  wire  _EVAL_1786;
  wire  _EVAL_1789;
  wire  _EVAL_1792;
  wire  _EVAL_1793;
  wire  _EVAL_1794;
  wire  _EVAL_1795;
  wire  _EVAL_1798;
  wire  _EVAL_1800;
  wire  _EVAL_1801;
  wire  _EVAL_1802;
  wire  _EVAL_1804;
  wire  _EVAL_1807;
  wire  _EVAL_1808;
  wire  _EVAL_1810;
  wire  _EVAL_1811;
  wire  _EVAL_1814;
  wire  _EVAL_1816;
  wire  _EVAL_1818;
  wire  _EVAL_1819;
  wire  _EVAL_1824;
  wire  _EVAL_1830;
  wire  _EVAL_1832;
  wire  _EVAL_1833;
  wire  _EVAL_1835;
  wire  _EVAL_1836;
  wire  _EVAL_1837;
  wire  _EVAL_1838;
  wire  _EVAL_1839;
  wire  _EVAL_1840;
  wire  _EVAL_1841;
  wire  _EVAL_1845;
  wire  _EVAL_1846;
  wire  _EVAL_1847;
  wire  _EVAL_1850;
  wire  _EVAL_1852;
  wire  _EVAL_1853;
  wire  _EVAL_1854;
  wire  _EVAL_1856;
  wire  _EVAL_1858;
  wire  _EVAL_1861;
  wire  _EVAL_1862;
  wire  _EVAL_1865;
  wire  _EVAL_1867;
  wire  _EVAL_1869;
  wire  _EVAL_1870;
  wire  _EVAL_1876;
  wire  _EVAL_1878;
  wire  _EVAL_1879;
  wire  _EVAL_1881;
  wire  _EVAL_1884;
  wire  _EVAL_1887;
  wire  _EVAL_1888;
  wire  _EVAL_1889;
  wire  _EVAL_1893;
  wire  _EVAL_1894;
  wire  _EVAL_1895;
  wire  _EVAL_1896;
  wire  _EVAL_1897;
  wire  _EVAL_1902;
  wire  _EVAL_1905;
  wire  _EVAL_1906;
  wire  _EVAL_1909;
  wire  _EVAL_1910;
  wire  _EVAL_1911;
  wire  _EVAL_1913;
  wire  _EVAL_1915;
  wire  _EVAL_1916;
  wire  _EVAL_1919;
  wire  _EVAL_1920;
  wire  _EVAL_1921;
  wire  _EVAL_1924;
  wire  _EVAL_1926;
  wire  _EVAL_1928;
  wire  _EVAL_1931;
  wire  _EVAL_1932;
  wire  _EVAL_1933;
  wire  _EVAL_1936;
  wire  _EVAL_1938;
  wire  _EVAL_1940;
  wire  _EVAL_1941;
  wire  _EVAL_1944;
  wire  _EVAL_1945;
  wire  _EVAL_1946;
  wire  _EVAL_1947;
  wire  _EVAL_1948;
  wire  _EVAL_1951;
  wire  _EVAL_1954;
  wire  _EVAL_1955;
  wire  _EVAL_1957;
  wire  _EVAL_1958;
  wire  _EVAL_1960;
  wire  _EVAL_1962;
  wire  _EVAL_1965;
  wire  _EVAL_1966;
  wire  _EVAL_1971;
  wire  _EVAL_1972;
  wire  _EVAL_1973;
  wire  _EVAL_1974;
  wire  _EVAL_1975;
  wire  _EVAL_1977;
  wire  _EVAL_1978;
  wire  _EVAL_1980;
  wire  _EVAL_1981;
  wire  _EVAL_1984;
  wire  _EVAL_1985;
  wire  _EVAL_1986;
  wire  _EVAL_1988;
  wire [6:0] _EVAL_1989;
  wire  _EVAL_1991;
  wire  _EVAL_1992;
  wire  _EVAL_1993;
  wire  _EVAL_1994;
  wire  _EVAL_1995;
  wire  _EVAL_1996;
  wire  _EVAL_2000;
  wire  _EVAL_2001;
  wire  _EVAL_2002;
  wire  _EVAL_2005;
  wire  _EVAL_2006;
  wire  _EVAL_2007;
  wire  _EVAL_2008;
  wire  _EVAL_2011;
  wire  _EVAL_2012;
  wire  _EVAL_2014;
  wire  _EVAL_2015;
  wire  _EVAL_2019;
  wire  _EVAL_2021;
  wire  _EVAL_2023;
  wire  _EVAL_2027;
  wire  _EVAL_2028;
  wire  _EVAL_2031;
  wire  _EVAL_2032;
  wire  _EVAL_2033;
  wire  _EVAL_2035;
  wire  _EVAL_2037;
  wire  _EVAL_2038;
  wire  _EVAL_2039;
  wire  _EVAL_2040;
  wire  _EVAL_2041;
  wire  _EVAL_2043;
  wire  _EVAL_2044;
  wire  _EVAL_2045;
  wire  _EVAL_2049;
  wire  _EVAL_2051;
  wire  _EVAL_2059;
  wire  _EVAL_2060;
  wire  _EVAL_2062;
  wire  _EVAL_2064;
  wire  _EVAL_2066;
  wire  _EVAL_2067;
  wire  _EVAL_2068;
  wire  _EVAL_2069;
  wire  _EVAL_2071;
  wire  _EVAL_2072;
  wire  _EVAL_2073;
  wire  _EVAL_2075;
  wire  _EVAL_2076;
  wire  _EVAL_2078;
  wire  _EVAL_2079;
  wire  _EVAL_2082;
  wire  _EVAL_2083;
  wire  _EVAL_2084;
  wire  _EVAL_2087;
  wire  _EVAL_2088;
  wire  _EVAL_2089;
  wire  _EVAL_2093;
  wire  _EVAL_2095;
  wire  _EVAL_2097;
  wire  _EVAL_2100;
  wire  _EVAL_2103;
  wire  _EVAL_2106;
  wire  _EVAL_2107;
  wire  _EVAL_2110;
  wire  _EVAL_2116;
  wire  _EVAL_2117;
  wire  _EVAL_2118;
  wire  _EVAL_2121;
  wire  _EVAL_2123;
  wire  _EVAL_2124;
  wire  _EVAL_2125;
  wire  _EVAL_2126;
  wire  _EVAL_2127;
  wire  _EVAL_2129;
  wire  _EVAL_2131;
  wire  _EVAL_2133;
  wire  _EVAL_2134;
  wire  _EVAL_2135;
  wire  _EVAL_2140;
  wire  _EVAL_2142;
  wire  _EVAL_2144;
  wire  _EVAL_2145;
  wire  _EVAL_2149;
  wire  _EVAL_2150;
  wire  _EVAL_2151;
  wire  _EVAL_2153;
  wire  _EVAL_2163;
  wire  _EVAL_2165;
  wire  _EVAL_2167;
  wire  _EVAL_2169;
  wire  _EVAL_2170;
  wire  _EVAL_2171;
  wire  _EVAL_2172;
  wire  _EVAL_2174;
  wire  _EVAL_2175;
  wire  _EVAL_2179;
  wire  _EVAL_2181;
  wire  _EVAL_2184;
  wire  _EVAL_2187;
  wire  _EVAL_2191;
  wire  _EVAL_2192;
  wire  _EVAL_2193;
  wire  _EVAL_2194;
  wire  _EVAL_2195;
  wire  _EVAL_2200;
  wire  _EVAL_2204;
  wire  _EVAL_2205;
  wire  _EVAL_2207;
  wire  _EVAL_2208;
  wire  _EVAL_2209;
  wire  _EVAL_2210;
  wire  _EVAL_2213;
  wire  _EVAL_2214;
  wire  _EVAL_2217;
  wire  _EVAL_2219;
  wire  _EVAL_2220;
  wire  _EVAL_2221;
  wire  _EVAL_2222;
  wire  _EVAL_2223;
  wire  _EVAL_2224;
  wire  _EVAL_2230;
  wire  _EVAL_2232;
  wire  _EVAL_2235;
  wire [3:0] _EVAL_2236;
  wire  _EVAL_2238;
  wire  _EVAL_2241;
  wire  _EVAL_2242;
  wire  _EVAL_2243;
  wire  _EVAL_2245;
  wire  _EVAL_2246;
  wire  _EVAL_2250;
  wire  _EVAL_2251;
  wire  _EVAL_2252;
  wire  _EVAL_2253;
  wire  _EVAL_2254;
  wire  _EVAL_2255;
  wire  _EVAL_2256;
  wire  _EVAL_2258;
  wire  _EVAL_2260;
  wire  _EVAL_2262;
  wire  _EVAL_2266;
  wire  _EVAL_2268;
  wire  _EVAL_2269;
  wire  _EVAL_2270;
  wire  _EVAL_2271;
  wire  _EVAL_2272;
  wire  _EVAL_2273;
  wire  _EVAL_2274;
  wire  _EVAL_2275;
  wire  _EVAL_2278;
  wire  _EVAL_2280;
  wire  _EVAL_2284;
  wire  _EVAL_2285;
  wire  _EVAL_2288;
  wire  _EVAL_2290;
  wire  _EVAL_2292;
  wire  _EVAL_2294;
  wire  _EVAL_2295;
  wire  _EVAL_2296;
  wire  _EVAL_2297;
  wire  _EVAL_2298;
  wire  _EVAL_2299;
  wire  _EVAL_2302;
  wire  _EVAL_2304;
  wire  _EVAL_2305;
  wire  _EVAL_2306;
  wire  _EVAL_2310;
  wire  _EVAL_2313;
  wire  _EVAL_2314;
  wire  _EVAL_2317;
  wire  _EVAL_2318;
  wire  _EVAL_2320;
  wire  _EVAL_2321;
  wire  _EVAL_2323;
  wire  _EVAL_2325;
  wire  _EVAL_2326;
  wire  _EVAL_2327;
  wire  _EVAL_2328;
  wire  _EVAL_2329;
  wire  _EVAL_2333;
  wire  _EVAL_2334;
  wire  _EVAL_2335;
  wire  _EVAL_2338;
  wire  _EVAL_2340;
  wire  _EVAL_2344;
  wire  _EVAL_2345;
  wire  _EVAL_2347;
  wire  _EVAL_2349;
  wire  _EVAL_2354;
  wire  _EVAL_2355;
  wire  _EVAL_2356;
  wire  _EVAL_2358;
  wire  _EVAL_2361;
  wire  _EVAL_2362;
  wire  _EVAL_2363;
  wire  _EVAL_2364;
  wire  _EVAL_2367;
  wire  _EVAL_2368;
  wire  _EVAL_2370;
  wire  _EVAL_2371;
  wire  _EVAL_2373;
  wire  _EVAL_2375;
  wire  _EVAL_2376;
  wire  _EVAL_2378;
  wire  _EVAL_2379;
  wire  _EVAL_2382;
  wire  _EVAL_2383;
  wire  _EVAL_2384;
  wire  _EVAL_2386;
  wire  _EVAL_2387;
  wire  _EVAL_2388;
  wire  _EVAL_2390;
  wire  _EVAL_2395;
  wire  _EVAL_2397;
  wire  _EVAL_2399;
  wire  _EVAL_2401;
  wire  _EVAL_2402;
  wire  _EVAL_2403;
  wire  _EVAL_2404;
  wire  _EVAL_2405;
  wire  _EVAL_2409;
  wire  _EVAL_2411;
  wire  _EVAL_2412;
  wire  _EVAL_2414;
  wire  _EVAL_2416;
  wire  _EVAL_2419;
  wire  _EVAL_2420;
  wire  _EVAL_2423;
  wire  _EVAL_2424;
  wire  _EVAL_2425;
  wire  _EVAL_2426;
  wire  _EVAL_2427;
  wire  _EVAL_2430;
  wire  _EVAL_2431;
  wire  _EVAL_2432;
  wire  _EVAL_2433;
  wire  _EVAL_2436;
  wire  _EVAL_2437;
  wire  _EVAL_2438;
  wire  _EVAL_2440;
  wire  _EVAL_2441;
  wire  _EVAL_2442;
  wire  _EVAL_2443;
  wire  _EVAL_2445;
  wire  _EVAL_2449;
  wire  _EVAL_2451;
  wire  _EVAL_2452;
  wire  _EVAL_2453;
  wire  _EVAL_2454;
  wire  _EVAL_2455;
  wire  _EVAL_2456;
  wire  _EVAL_2458;
  wire  _EVAL_2459;
  wire  _EVAL_2460;
  wire  _EVAL_2464;
  wire  _EVAL_2465;
  wire  _EVAL_2466;
  wire  _EVAL_2468;
  wire  _EVAL_2469;
  wire  _EVAL_2471;
  wire  _EVAL_2472;
  wire  _EVAL_2475;
  wire  _EVAL_2476;
  wire  _EVAL_2478;
  wire  _EVAL_2479;
  wire  _EVAL_2480;
  wire  _EVAL_2482;
  wire  _EVAL_2483;
  wire  _EVAL_2485;
  wire  _EVAL_2494;
  wire  _EVAL_2496;
  wire  _EVAL_2497;
  wire  _EVAL_2498;
  wire  _EVAL_2500;
  wire  _EVAL_2502;
  wire  _EVAL_2504;
  wire  _EVAL_2505;
  wire  _EVAL_2506;
  wire  _EVAL_2507;
  wire  _EVAL_2509;
  wire  _EVAL_2511;
  wire  _EVAL_2513;
  wire  _EVAL_2514;
  wire  _EVAL_2517;
  wire  _EVAL_2518;
  wire  _EVAL_2524;
  wire  _EVAL_2525;
  wire  _EVAL_2526;
  wire  _EVAL_2529;
  wire  _EVAL_2531;
  wire  _EVAL_2533;
  wire  _EVAL_2536;
  wire  _EVAL_2538;
  wire  _EVAL_2539;
  wire  _EVAL_2540;
  wire  _EVAL_2542;
  wire  _EVAL_2545;
  wire  _EVAL_2548;
  wire  _EVAL_2550;
  wire  _EVAL_2551;
  wire  _EVAL_2552;
  wire  _EVAL_2553;
  wire  _EVAL_2554;
  wire  _EVAL_2555;
  wire  _EVAL_2556;
  wire  _EVAL_2558;
  wire  _EVAL_2560;
  wire  _EVAL_2562;
  wire  _EVAL_2564;
  wire  _EVAL_2565;
  wire  _EVAL_2567;
  wire  _EVAL_2569;
  wire  _EVAL_2570;
  wire  _EVAL_2571;
  wire  _EVAL_2572;
  wire  _EVAL_2573;
  wire  _EVAL_2574;
  wire  _EVAL_2576;
  wire  _EVAL_2581;
  wire  _EVAL_2582;
  wire  _EVAL_2584;
  wire  _EVAL_2585;
  wire  _EVAL_2588;
  wire  _EVAL_2592;
  wire  _EVAL_2593;
  wire  _EVAL_2594;
  wire  _EVAL_2597;
  wire  _EVAL_2599;
  wire  _EVAL_2601;
  wire  _EVAL_2602;
  wire  _EVAL_2604;
  wire  _EVAL_2606;
  wire  _EVAL_2607;
  wire  _EVAL_2608;
  wire  _EVAL_2609;
  wire  _EVAL_2612;
  wire  _EVAL_2613;
  wire  _EVAL_2614;
  wire  _EVAL_2615;
  wire  _EVAL_2617;
  wire  _EVAL_2619;
  wire  _EVAL_2620;
  wire  _EVAL_2624;
  wire  _EVAL_2625;
  wire  _EVAL_2627;
  wire  _EVAL_2628;
  wire  _EVAL_2631;
  wire  _EVAL_2632;
  wire  _EVAL_2634;
  wire  _EVAL_2640;
  wire  _EVAL_2643;
  wire  _EVAL_2644;
  wire  _EVAL_2645;
  wire  _EVAL_2646;
  wire  _EVAL_2647;
  wire  _EVAL_2649;
  wire  _EVAL_2650;
  wire  _EVAL_2651;
  wire  _EVAL_2652;
  wire  _EVAL_2653;
  wire  _EVAL_2655;
  wire  _EVAL_2656;
  wire  _EVAL_2657;
  wire  _EVAL_2658;
  wire  _EVAL_2659;
  wire  _EVAL_2662;
  wire  _EVAL_2663;
  wire  _EVAL_2665;
  wire  _EVAL_2670;
  wire  _EVAL_2672;
  wire  _EVAL_2673;
  wire  _EVAL_2675;
  wire  _EVAL_2676;
  wire  _EVAL_2677;
  wire  _EVAL_2678;
  wire  _EVAL_2679;
  wire  _EVAL_2680;
  wire  _EVAL_2682;
  wire  _EVAL_2684;
  wire  _EVAL_2685;
  wire  _EVAL_2686;
  wire  _EVAL_2687;
  wire [3:0] _EVAL_2688;
  wire  _EVAL_2689;
  wire  _EVAL_2695;
  wire  _EVAL_2698;
  wire  _EVAL_2699;
  wire  _EVAL_2700;
  wire  _EVAL_2702;
  wire  _EVAL_2704;
  wire  _EVAL_2705;
  wire  _EVAL_2708;
  wire  _EVAL_2710;
  wire  _EVAL_2712;
  wire  _EVAL_2713;
  wire  _EVAL_2715;
  wire  _EVAL_2718;
  wire  _EVAL_2720;
  wire  _EVAL_2721;
  wire  _EVAL_2723;
  wire  _EVAL_2724;
  wire  _EVAL_2725;
  wire  _EVAL_2726;
  wire  _EVAL_2729;
  wire  _EVAL_2730;
  wire  _EVAL_2731;
  wire  _EVAL_2732;
  wire  _EVAL_2733;
  wire  _EVAL_2734;
  wire  _EVAL_2735;
  wire  _EVAL_2736;
  wire  _EVAL_2738;
  wire  _EVAL_2742;
  wire  _EVAL_2744;
  wire  _EVAL_2745;
  wire  _EVAL_2746;
  wire  _EVAL_2748;
  wire  _EVAL_2750;
  wire [21:0] _EVAL_2753;
  wire  _EVAL_2754;
  wire  _EVAL_2759;
  wire  _EVAL_2762;
  wire  _EVAL_2763;
  wire  _EVAL_2768;
  wire  _EVAL_2769;
  wire  _EVAL_2770;
  wire  _EVAL_2771;
  wire  _EVAL_2772;
  wire  _EVAL_2773;
  wire  _EVAL_2775;
  wire  _EVAL_2783;
  wire  _EVAL_2785;
  wire  _EVAL_2789;
  wire  _EVAL_2790;
  wire  _EVAL_2791;
  wire  _EVAL_2792;
  wire  _EVAL_2793;
  wire  _EVAL_2795;
  wire  _EVAL_2796;
  wire [3:0] _EVAL_2798;
  wire  _EVAL_2799;
  wire  _EVAL_2803;
  wire  _EVAL_2807;
  wire  _EVAL_2808;
  wire  _EVAL_2809;
  wire  _EVAL_2810;
  wire  _EVAL_2814;
  wire  _EVAL_2816;
  wire  _EVAL_2817;
  wire  _EVAL_2818;
  wire  _EVAL_2821;
  wire  _EVAL_2822;
  wire  _EVAL_2830;
  wire  _EVAL_2831;
  wire  _EVAL_2833;
  wire  _EVAL_2834;
  wire  _EVAL_2835;
  wire  _EVAL_2836;
  wire  _EVAL_2839;
  wire  _EVAL_2842;
  wire  _EVAL_2844;
  wire  _EVAL_2846;
  wire  _EVAL_2849;
  wire  _EVAL_2850;
  wire  _EVAL_2858;
  wire  _EVAL_2859;
  wire  _EVAL_2860;
  wire  _EVAL_2863;
  wire  _EVAL_2868;
  wire  _EVAL_2870;
  wire  _EVAL_2871;
  wire  _EVAL_2872;
  wire  _EVAL_2873;
  wire  _EVAL_2875;
  wire  _EVAL_2877;
  wire  _EVAL_2879;
  wire  _EVAL_2881;
  wire  _EVAL_2885;
  wire  _EVAL_2886;
  wire  _EVAL_2888;
  wire  _EVAL_2890;
  wire  _EVAL_2891;
  wire  _EVAL_2892;
  wire  _EVAL_2893;
  wire  _EVAL_2897;
  wire  _EVAL_2899;
  wire  _EVAL_2900;
  wire  _EVAL_2902;
  wire  _EVAL_2903;
  wire  _EVAL_2904;
  wire  _EVAL_2906;
  wire  _EVAL_2907;
  wire  _EVAL_2908;
  wire  _EVAL_2909;
  wire  _EVAL_2911;
  wire  _EVAL_2913;
  wire  _EVAL_2916;
  wire  _EVAL_2917;
  wire  _EVAL_2919;
  wire  _EVAL_2921;
  wire  _EVAL_2923;
  wire  _EVAL_2924;
  wire  _EVAL_2925;
  wire  _EVAL_2926;
  wire  _EVAL_2927;
  wire  _EVAL_2930;
  wire  _EVAL_2931;
  wire  _EVAL_2934;
  wire  _EVAL_2937;
  wire  _EVAL_2939;
  wire  _EVAL_2941;
  wire  _EVAL_2942;
  wire [6:0] _EVAL_2945;
  wire  _EVAL_2946;
  wire  _EVAL_2947;
  wire  _EVAL_2950;
  wire  _EVAL_2953;
  wire  _EVAL_2955;
  wire  _EVAL_2956;
  wire  _EVAL_2957;
  wire  _EVAL_2960;
  wire  _EVAL_2962;
  wire  _EVAL_2963;
  wire  _EVAL_2965;
  wire  _EVAL_2966;
  wire  _EVAL_2969;
  wire  _EVAL_2972;
  wire  _EVAL_2973;
  wire  _EVAL_2974;
  wire  _EVAL_2975;
  wire  _EVAL_2976;
  wire  _EVAL_2977;
  wire  _EVAL_2982;
  wire  _EVAL_2983;
  wire  _EVAL_2985;
  wire  _EVAL_2986;
  wire  _EVAL_2987;
  wire  _EVAL_2990;
  wire  _EVAL_2991;
  wire  _EVAL_2992;
  wire  _EVAL_2998;
  wire  _EVAL_2999;
  wire  _EVAL_3000;
  wire  _EVAL_3002;
  wire  _EVAL_3004;
  wire  _EVAL_3006;
  wire  _EVAL_3007;
  wire  _EVAL_3008;
  wire  _EVAL_3009;
  wire  _EVAL_3010;
  wire  _EVAL_3013;
  wire  _EVAL_3014;
  wire  _EVAL_3015;
  wire  _EVAL_3021;
  wire  _EVAL_3025;
  wire  _EVAL_3026;
  wire  _EVAL_3028;
  wire  _EVAL_3029;
  wire  _EVAL_3032;
  wire  _EVAL_3033;
  wire  _EVAL_3034;
  wire  _EVAL_3038;
  wire  _EVAL_3041;
  wire  _EVAL_3049;
  wire  _EVAL_3050;
  wire  _EVAL_3052;
  wire  _EVAL_3054;
  wire [3:0] _EVAL_3055;
  wire  _EVAL_3057;
  wire  _EVAL_3060;
  wire  _EVAL_3061;
  wire  _EVAL_3063;
  wire  _EVAL_3065;
  wire  _EVAL_3066;
  wire  _EVAL_3068;
  wire  _EVAL_3069;
  wire  _EVAL_3070;
  wire  _EVAL_3071;
  wire  _EVAL_3072;
  wire  _EVAL_3073;
  wire  _EVAL_3074;
  wire  _EVAL_3075;
  wire  _EVAL_3076;
  wire  _EVAL_3077;
  wire  _EVAL_3078;
  wire  _EVAL_3079;
  wire  _EVAL_3081;
  wire  _EVAL_3082;
  wire  _EVAL_3084;
  wire  _EVAL_3085;
  wire  _EVAL_3089;
  wire  _EVAL_3091;
  wire  _EVAL_3095;
  wire  _EVAL_3097;
  wire  _EVAL_3101;
  wire  _EVAL_3103;
  wire  _EVAL_3106;
  wire  _EVAL_3107;
  wire  _EVAL_3109;
  wire  _EVAL_3112;
  wire  _EVAL_3113;
  wire  _EVAL_3116;
  wire  _EVAL_3117;
  wire  _EVAL_3118;
  wire  _EVAL_3121;
  wire  _EVAL_3122;
  wire  _EVAL_3124;
  wire  _EVAL_3130;
  wire  _EVAL_3132;
  wire  _EVAL_3134;
  wire  _EVAL_3135;
  wire [7:0] _EVAL_3136;
  wire  _EVAL_3137;
  wire  _EVAL_3138;
  wire  _EVAL_3139;
  wire  _EVAL_3142;
  wire  _EVAL_3143;
  wire  _EVAL_3147;
  wire  _EVAL_3151;
  wire  _EVAL_3153;
  wire  _EVAL_3155;
  wire  _EVAL_3156;
  wire  _EVAL_3157;
  wire  _EVAL_3159;
  wire  _EVAL_3160;
  wire  _EVAL_3161;
  wire  _EVAL_3162;
  wire  _EVAL_3163;
  wire  _EVAL_3166;
  wire  _EVAL_3167;
  wire  _EVAL_3170;
  wire  _EVAL_3174;
  wire  _EVAL_3175;
  wire  _EVAL_3176;
  wire  _EVAL_3177;
  wire  _EVAL_3178;
  wire  _EVAL_3179;
  wire  _EVAL_3180;
  wire  _EVAL_3182;
  wire  _EVAL_3183;
  wire  _EVAL_3184;
  wire  _EVAL_3185;
  wire  _EVAL_3186;
  wire  _EVAL_3187;
  wire  _EVAL_3188;
  wire  _EVAL_3192;
  wire  _EVAL_3195;
  wire  _EVAL_3198;
  wire  _EVAL_3199;
  wire  _EVAL_3201;
  wire  _EVAL_3202;
  wire  _EVAL_3206;
  wire  _EVAL_3208;
  wire  _EVAL_3209;
  wire  _EVAL_3210;
  wire  _EVAL_3214;
  wire  _EVAL_3216;
  wire  _EVAL_3218;
  wire  _EVAL_3220;
  wire  _EVAL_3221;
  wire  _EVAL_3223;
  wire  _EVAL_3224;
  wire  _EVAL_3226;
  wire  _EVAL_3227;
  wire  _EVAL_3228;
  wire  _EVAL_3231;
  wire  _EVAL_3232;
  wire  _EVAL_3235;
  wire [3:0] _EVAL_3236;
  wire  _EVAL_3237;
  wire  _EVAL_3238;
  wire  _EVAL_3239;
  wire  _EVAL_3240;
  wire  _EVAL_3241;
  wire  _EVAL_3242;
  wire  _EVAL_3243;
  wire  _EVAL_3244;
  wire  _EVAL_3245;
  wire  _EVAL_3246;
  wire  _EVAL_3247;
  wire  _EVAL_3248;
  wire  _EVAL_3249;
  wire  _EVAL_3250;
  wire  _EVAL_3251;
  wire  _EVAL_3252;
  wire  _EVAL_3257;
  wire  _EVAL_3258;
  wire  _EVAL_3260;
  wire  _EVAL_3261;
  wire  _EVAL_3262;
  wire  _EVAL_3263;
  wire [21:0] _EVAL_3264;
  wire  _EVAL_3265;
  wire  _EVAL_3267;
  wire  _EVAL_3269;
  wire  _EVAL_3276;
  wire  _EVAL_3279;
  wire  _EVAL_3281;
  wire  _EVAL_3282;
  wire  _EVAL_3284;
  wire  _EVAL_3287;
  wire  _EVAL_3288;
  wire  _EVAL_3292;
  wire  _EVAL_3295;
  wire  _EVAL_3296;
  wire  _EVAL_3300;
  wire  _EVAL_3301;
  wire  _EVAL_3302;
  wire  _EVAL_3303;
  wire  _EVAL_3305;
  wire  _EVAL_3306;
  wire  _EVAL_3307;
  wire  _EVAL_3312;
  wire  _EVAL_3313;
  wire  _EVAL_3314;
  wire  _EVAL_3315;
  wire  _EVAL_3316;
  wire [6:0] _EVAL_3321;
  wire  _EVAL_3322;
  wire  _EVAL_3323;
  wire  _EVAL_3326;
  wire  _EVAL_3328;
  wire  _EVAL_3329;
  wire  _EVAL_3331;
  wire  _EVAL_3333;
  wire  _EVAL_3337;
  wire  _EVAL_3338;
  wire  _EVAL_3340;
  wire  _EVAL_3342;
  wire  _EVAL_3346;
  wire  _EVAL_3347;
  wire  _EVAL_3348;
  wire  _EVAL_3349;
  wire [30:0] _EVAL_3350;
  wire  _EVAL_3352;
  wire  _EVAL_3354;
  wire  _EVAL_3360;
  wire  _EVAL_3361;
  wire  _EVAL_3362;
  wire  _EVAL_3364;
  wire  _EVAL_3366;
  wire  _EVAL_3367;
  wire  _EVAL_3369;
  wire  _EVAL_3370;
  wire  _EVAL_3371;
  wire  _EVAL_3373;
  wire  _EVAL_3375;
  wire  _EVAL_3376;
  wire  _EVAL_3377;
  wire  _EVAL_3379;
  wire  _EVAL_3381;
  wire  _EVAL_3382;
  wire  _EVAL_3386;
  wire  _EVAL_3387;
  wire  _EVAL_3388;
  wire  _EVAL_3394;
  wire  _EVAL_3396;
  wire  _EVAL_3398;
  wire  _EVAL_3399;
  wire  _EVAL_3400;
  wire  _EVAL_3401;
  wire  _EVAL_3402;
  wire  _EVAL_3403;
  wire  _EVAL_3406;
  wire  _EVAL_3407;
  wire  _EVAL_3409;
  wire  _EVAL_3412;
  wire  _EVAL_3413;
  wire  _EVAL_3414;
  wire  _EVAL_3417;
  wire  _EVAL_3418;
  wire [7:0] _EVAL_3420;
  wire  _EVAL_3421;
  wire  _EVAL_3424;
  wire  _EVAL_3425;
  wire  _EVAL_3432;
  wire  _EVAL_3433;
  wire  _EVAL_3436;
  wire  _EVAL_3437;
  wire  _EVAL_3440;
  wire  _EVAL_3445;
  wire  _EVAL_3447;
  wire  _EVAL_3448;
  wire  _EVAL_3451;
  wire  _EVAL_3453;
  wire  _EVAL_3455;
  wire  _EVAL_3457;
  wire  _EVAL_3458;
  wire  _EVAL_3459;
  wire  _EVAL_3461;
  wire  _EVAL_3462;
  wire  _EVAL_3468;
  wire  _EVAL_3470;
  wire  _EVAL_3471;
  wire  _EVAL_3473;
  wire  _EVAL_3474;
  wire  _EVAL_3476;
  wire  _EVAL_3478;
  wire  _EVAL_3480;
  wire  _EVAL_3481;
  wire  _EVAL_3484;
  wire [9:0] _EVAL_3485;
  wire  _EVAL_3486;
  wire  _EVAL_3488;
  wire  _EVAL_3489;
  wire  _EVAL_3490;
  wire  _EVAL_3491;
  wire  _EVAL_3492;
  wire  _EVAL_3495;
  wire  _EVAL_3497;
  wire  _EVAL_3500;
  wire  _EVAL_3503;
  wire  _EVAL_3505;
  wire  _EVAL_3506;
  wire  _EVAL_3508;
  wire  _EVAL_3509;
  wire  _EVAL_3510;
  wire  _EVAL_3511;
  wire  _EVAL_3512;
  wire  _EVAL_3514;
  wire  _EVAL_3515;
  wire  _EVAL_3519;
  wire  _EVAL_3520;
  wire  _EVAL_3522;
  wire  _EVAL_3523;
  wire  _EVAL_3524;
  wire  _EVAL_3525;
  wire  _EVAL_3528;
  wire  _EVAL_3529;
  wire  _EVAL_3531;
  wire  _EVAL_3536;
  wire  _EVAL_3539;
  wire  _EVAL_3540;
  wire  _EVAL_3543;
  wire  _EVAL_3545;
  wire  _EVAL_3547;
  wire  _EVAL_3548;
  wire  _EVAL_3551;
  wire  _EVAL_3552;
  wire  _EVAL_3553;
  wire  _EVAL_3556;
  wire  _EVAL_3557;
  wire  _EVAL_3558;
  wire  _EVAL_3562;
  wire  _EVAL_3565;
  wire  _EVAL_3566;
  wire  _EVAL_3568;
  wire  _EVAL_3569;
  wire  _EVAL_3571;
  wire  _EVAL_3572;
  wire  _EVAL_3574;
  wire  _EVAL_3575;
  wire  _EVAL_3577;
  wire  _EVAL_3579;
  wire  _EVAL_3581;
  wire  _EVAL_3582;
  wire  _EVAL_3583;
  wire [3:0] _EVAL_3586;
  wire  _EVAL_3588;
  wire  _EVAL_3592;
  wire  _EVAL_3593;
  wire  _EVAL_3595;
  wire  _EVAL_3596;
  wire  _EVAL_3598;
  wire  _EVAL_3600;
  wire  _EVAL_3601;
  wire  _EVAL_3602;
  wire  _EVAL_3608;
  wire  _EVAL_3610;
  wire  _EVAL_3611;
  wire  _EVAL_3616;
  wire  _EVAL_3617;
  wire  _EVAL_3622;
  wire  _EVAL_3624;
  wire  _EVAL_3626;
  wire  _EVAL_3628;
  wire  _EVAL_3630;
  wire  _EVAL_3631;
  wire  _EVAL_3632;
  wire  _EVAL_3638;
  wire  _EVAL_3640;
  wire  _EVAL_3647;
  wire  _EVAL_3648;
  wire  _EVAL_3649;
  wire  _EVAL_3650;
  wire  _EVAL_3651;
  wire  _EVAL_3655;
  wire  _EVAL_3657;
  wire  _EVAL_3658;
  wire  _EVAL_3659;
  wire  _EVAL_3660;
  wire  _EVAL_3663;
  wire  _EVAL_3664;
  wire  _EVAL_3669;
  wire  _EVAL_3672;
  wire  _EVAL_3677;
  wire  _EVAL_3678;
  wire  _EVAL_3679;
  wire  _EVAL_3680;
  wire  _EVAL_3684;
  wire  _EVAL_3687;
  wire  _EVAL_3688;
  wire  _EVAL_3689;
  wire  _EVAL_3690;
  wire  _EVAL_3691;
  wire  _EVAL_3694;
  wire  _EVAL_3695;
  wire  _EVAL_3698;
  wire  _EVAL_3699;
  wire  _EVAL_3700;
  wire  _EVAL_3701;
  wire  _EVAL_3702;
  wire  _EVAL_3704;
  wire  _EVAL_3706;
  wire  _EVAL_3707;
  wire  _EVAL_3708;
  wire  _EVAL_3710;
  wire  _EVAL_3712;
  wire  _EVAL_3714;
  wire  _EVAL_3718;
  wire  _EVAL_3719;
  wire  _EVAL_3720;
  wire  _EVAL_3721;
  wire  _EVAL_3723;
  wire  _EVAL_3725;
  wire  _EVAL_3727;
  wire  _EVAL_3728;
  wire  _EVAL_3730;
  wire  _EVAL_3734;
  wire  _EVAL_3736;
  wire  _EVAL_3738;
  wire  _EVAL_3740;
  wire  _EVAL_3744;
  wire  _EVAL_3746;
  wire  _EVAL_3747;
  wire  _EVAL_3749;
  wire  _EVAL_3754;
  wire  _EVAL_3755;
  wire  _EVAL_3759;
  wire  _EVAL_3760;
  wire  _EVAL_3761;
  wire  _EVAL_3764;
  wire  _EVAL_3766;
  wire  _EVAL_3768;
  wire  _EVAL_3769;
  wire  _EVAL_3770;
  wire  _EVAL_3773;
  wire  _EVAL_3774;
  wire  _EVAL_3776;
  wire  _EVAL_3777;
  wire  _EVAL_3778;
  wire  _EVAL_3780;
  wire  _EVAL_3781;
  wire  _EVAL_3782;
  wire  _EVAL_3784;
  wire  _EVAL_3785;
  wire  _EVAL_3787;
  wire  _EVAL_3792;
  wire  _EVAL_3794;
  wire  _EVAL_3801;
  wire  _EVAL_3802;
  wire  _EVAL_3803;
  wire  _EVAL_3804;
  wire  _EVAL_3807;
  wire  _EVAL_3809;
  wire  _EVAL_3811;
  wire  _EVAL_3812;
  wire  _EVAL_3813;
  wire  _EVAL_3815;
  wire  _EVAL_3816;
  wire  _EVAL_3817;
  wire  _EVAL_3818;
  wire [6:0] _EVAL_3820;
  wire  _EVAL_3821;
  wire  _EVAL_3822;
  wire  _EVAL_3825;
  wire  _EVAL_3826;
  wire  _EVAL_3828;
  wire  _EVAL_3829;
  wire  _EVAL_3830;
  wire  _EVAL_3833;
  wire  _EVAL_3835;
  wire  _EVAL_3837;
  wire  _EVAL_3840;
  wire  _EVAL_3841;
  wire  _EVAL_3842;
  wire  _EVAL_3844;
  wire  _EVAL_3845;
  wire  _EVAL_3849;
  wire  _EVAL_3850;
  wire  _EVAL_3852;
  wire  _EVAL_3853;
  wire  _EVAL_3856;
  wire  _EVAL_3858;
  wire  _EVAL_3859;
  wire  _EVAL_3860;
  wire  _EVAL_3863;
  wire  _EVAL_3867;
  wire  _EVAL_3868;
  wire  _EVAL_3869;
  wire [2:0] TLMonitor__EVAL;
  wire [1:0] TLMonitor__EVAL_0;
  wire  TLMonitor__EVAL_1;
  wire  TLMonitor__EVAL_2;
  wire [3:0] TLMonitor__EVAL_3;
  wire [2:0] TLMonitor__EVAL_4;
  wire [25:0] TLMonitor__EVAL_5;
  wire [1:0] TLMonitor__EVAL_6;
  wire  TLMonitor__EVAL_7;
  wire [2:0] TLMonitor__EVAL_8;
  wire  TLMonitor__EVAL_9;
  wire  TLMonitor__EVAL_10;
  wire  TLMonitor__EVAL_11;
  wire [2:0] TLMonitor__EVAL_12;
  wire [2:0] TLMonitor__EVAL_13;
  wire  TLMonitor__EVAL_14;
  wire  _EVAL_3873;
  wire  _EVAL_3874;
  wire  _EVAL_3875;
  wire  _EVAL_3878;
  wire  _EVAL_3880;
  wire  _EVAL_3881;
  wire [3:0] _EVAL_3882;
  wire  _EVAL_3884;
  wire  _EVAL_3886;
  wire  _EVAL_3888;
  wire  _EVAL_3889;
  wire  _EVAL_3894;
  wire  _EVAL_3896;
  wire  _EVAL_3897;
  wire  _EVAL_3898;
  wire  _EVAL_3901;
  wire  _EVAL_3902;
  wire  _EVAL_3904;
  wire  _EVAL_3908;
  wire  _EVAL_3909;
  wire  _EVAL_3910;
  wire  _EVAL_3917;
  wire  _EVAL_3919;
  wire  _EVAL_3920;
  wire  _EVAL_3923;
  wire  _EVAL_3924;
  wire  _EVAL_3926;
  wire  _EVAL_3928;
  wire  _EVAL_3931;
  wire  _EVAL_3932;
  wire  _EVAL_3933;
  wire  _EVAL_3935;
  wire  _EVAL_3942;
  wire  _EVAL_3943;
  wire  _EVAL_3948;
  wire  _EVAL_3949;
  wire  _EVAL_3951;
  wire  _EVAL_3952;
  wire  _EVAL_3953;
  wire  _EVAL_3954;
  wire  _EVAL_3955;
  wire  _EVAL_3956;
  wire  _EVAL_3957;
  wire  _EVAL_3959;
  wire  _EVAL_3961;
  wire  _EVAL_3964;
  wire  _EVAL_3966;
  wire  _EVAL_3968;
  wire  _EVAL_3969;
  wire  _EVAL_3972;
  wire  _EVAL_3973;
  wire  _EVAL_3974;
  wire  _EVAL_3976;
  wire  _EVAL_3978;
  wire  _EVAL_3981;
  wire  _EVAL_3982;
  wire  _EVAL_3984;
  wire  _EVAL_3988;
  wire  _EVAL_3990;
  wire  _EVAL_3991;
  wire  _EVAL_3992;
  wire  _EVAL_3993;
  wire  _EVAL_3994;
  wire  _EVAL_3995;
  wire  _EVAL_3996;
  wire  _EVAL_3998;
  wire  _EVAL_4001;
  wire  _EVAL_4002;
  wire  _EVAL_4006;
  wire  _EVAL_4011;
  wire  _EVAL_4016;
  wire  _EVAL_4017;
  wire  _EVAL_4018;
  wire  _EVAL_4020;
  wire  _EVAL_4022;
  wire  _EVAL_4023;
  wire  _EVAL_4024;
  wire  _EVAL_4027;
  wire  _EVAL_4028;
  wire  _EVAL_4029;
  wire  _EVAL_4031;
  wire  _EVAL_4033;
  wire  _EVAL_4034;
  wire  _EVAL_4035;
  wire  _EVAL_4038;
  wire  _EVAL_4039;
  wire  _EVAL_4042;
  wire  _EVAL_4043;
  wire  _EVAL_4044;
  wire  _EVAL_4047;
  wire  _EVAL_4048;
  wire  _EVAL_4049;
  wire  _EVAL_4052;
  wire  _EVAL_4054;
  wire  _EVAL_4057;
  wire  _EVAL_4059;
  wire  _EVAL_4060;
  wire  _EVAL_4061;
  wire  _EVAL_4062;
  wire  _EVAL_4063;
  wire  _EVAL_4066;
  wire  _EVAL_4069;
  wire  _EVAL_4071;
  wire  _EVAL_4072;
  wire  _EVAL_4073;
  wire  _EVAL_4075;
  wire  _EVAL_4077;
  wire  _EVAL_4078;
  wire  _EVAL_4079;
  wire  _EVAL_4082;
  wire  _EVAL_4083;
  wire  _EVAL_4084;
  wire  _EVAL_4086;
  wire  _EVAL_4091;
  wire  _EVAL_4092;
  wire  _EVAL_4093;
  wire  _EVAL_4094;
  wire  _EVAL_4095;
  wire  _EVAL_4097;
  wire  _EVAL_4099;
  wire  _EVAL_4100;
  wire  _EVAL_4101;
  wire  _EVAL_4102;
  wire  _EVAL_4104;
  wire  _EVAL_4106;
  wire  _EVAL_4108;
  wire  _EVAL_4109;
  wire  _EVAL_4110;
  wire  _EVAL_4111;
  wire  _EVAL_4112;
  wire  _EVAL_4113;
  wire  _EVAL_4114;
  wire  _EVAL_4118;
  wire  _EVAL_4120;
  wire  _EVAL_4121;
  wire  _EVAL_4125;
  wire  _EVAL_4126;
  wire  _EVAL_4129;
  wire  _EVAL_4130;
  wire  _EVAL_4132;
  wire  _EVAL_4133;
  wire  _EVAL_4134;
  wire  _EVAL_4135;
  wire  _EVAL_4137;
  wire  _EVAL_4138;
  wire  _EVAL_4139;
  wire  _EVAL_4140;
  wire  _EVAL_4141;
  wire  _EVAL_4144;
  wire  _EVAL_4145;
  wire  _EVAL_4146;
  wire  _EVAL_4149;
  wire  _EVAL_4150;
  wire  _EVAL_4151;
  wire  _EVAL_4152;
  wire  _EVAL_4154;
  wire  _EVAL_4155;
  wire  _EVAL_4157;
  wire  _EVAL_4158;
  wire  _EVAL_4160;
  wire  _EVAL_4163;
  wire  _EVAL_4166;
  wire  _EVAL_4171;
  wire  _EVAL_4175;
  wire  _EVAL_4180;
  wire  _EVAL_4183;
  wire  _EVAL_4185;
  wire  _EVAL_4186;
  wire  _EVAL_4187;
  wire  _EVAL_4188;
  wire  _EVAL_4189;
  wire  _EVAL_4190;
  wire  _EVAL_4191;
  wire  _EVAL_4192;
  wire  _EVAL_4193;
  wire  _EVAL_4194;
  wire  _EVAL_4196;
  wire  _EVAL_4200;
  wire  _EVAL_4201;
  wire  _EVAL_4202;
  wire  _EVAL_4203;
  wire  _EVAL_4205;
  wire  _EVAL_4206;
  wire  _EVAL_4207;
  wire  _EVAL_4208;
  wire  _EVAL_4209;
  wire  _EVAL_4210;
  wire  _EVAL_4211;
  wire  _EVAL_4212;
  wire  _EVAL_4214;
  wire  _EVAL_4216;
  wire  _EVAL_4218;
  wire  _EVAL_4219;
  wire  _EVAL_4220;
  wire  _EVAL_4222;
  wire  _EVAL_4223;
  wire  _EVAL_4224;
  wire  _EVAL_4225;
  wire  _EVAL_4227;
  wire  _EVAL_4228;
  wire  _EVAL_4230;
  wire  _EVAL_4231;
  wire  _EVAL_4232;
  wire  _EVAL_4235;
  wire  _EVAL_4239;
  wire  _EVAL_4240;
  wire  _EVAL_4241;
  wire  _EVAL_4243;
  wire  _EVAL_4245;
  wire  _EVAL_4248;
  wire  _EVAL_4253;
  wire  _EVAL_4254;
  wire  _EVAL_4257;
  wire  _EVAL_4258;
  wire  _EVAL_4259;
  wire  _EVAL_4261;
  wire  _EVAL_4263;
  wire  _EVAL_4265;
  wire  _EVAL_4269;
  wire  _EVAL_4270;
  wire  _EVAL_4273;
  wire  _EVAL_4276;
  wire  _EVAL_4277;
  wire  _EVAL_4278;
  wire  _EVAL_4279;
  wire  _EVAL_4280;
  wire  _EVAL_4281;
  wire  _EVAL_4283;
  wire  _EVAL_4287;
  wire  _EVAL_4288;
  wire  _EVAL_4289;
  wire  _EVAL_4293;
  wire  _EVAL_4294;
  wire  _EVAL_4295;
  wire  _EVAL_4299;
  wire  _EVAL_4300;
  wire  _EVAL_4302;
  wire  _EVAL_4305;
  wire  _EVAL_4306;
  wire  _EVAL_4309;
  wire  _EVAL_4310;
  wire  _EVAL_4311;
  wire  _EVAL_4312;
  wire  _EVAL_4314;
  wire  _EVAL_4315;
  wire  _EVAL_4316;
  wire  _EVAL_4317;
  wire  _EVAL_4319;
  wire  _EVAL_4320;
  wire  _EVAL_4322;
  wire  _EVAL_4323;
  wire  _EVAL_4324;
  wire  _EVAL_4325;
  wire  _EVAL_4326;
  wire  _EVAL_4327;
  wire  _EVAL_4329;
  wire  _EVAL_4330;
  wire  _EVAL_4332;
  wire  _EVAL_4333;
  wire  _EVAL_4334;
  wire  _EVAL_4335;
  wire  _EVAL_4341;
  wire  _EVAL_4342;
  wire  _EVAL_4343;
  wire  _EVAL_4346;
  wire  _EVAL_4350;
  wire  _EVAL_4351;
  wire  _EVAL_4353;
  wire  _EVAL_4357;
  wire  _EVAL_4359;
  wire  _EVAL_4361;
  wire  _EVAL_4362;
  wire  _EVAL_4363;
  wire  _EVAL_4364;
  wire  _EVAL_4365;
  wire  _EVAL_4366;
  wire  _EVAL_4369;
  wire  _EVAL_4371;
  wire  _EVAL_4372;
  wire  _EVAL_4373;
  wire  _EVAL_4375;
  wire  _EVAL_4378;
  wire  _EVAL_4379;
  wire  _EVAL_4380;
  wire  _EVAL_4381;
  wire  _EVAL_4383;
  wire  _EVAL_4385;
  wire  _EVAL_4389;
  wire  _EVAL_4391;
  wire  _EVAL_4392;
  wire  _EVAL_4393;
  wire  _EVAL_4394;
  wire  _EVAL_4395;
  wire  _EVAL_4399;
  wire  _EVAL_4405;
  wire  _EVAL_4407;
  wire  _EVAL_4408;
  wire  _EVAL_4409;
  wire  _EVAL_4411;
  wire  _EVAL_4413;
  wire  _EVAL_4419;
  wire  _EVAL_4420;
  wire  _EVAL_4422;
  wire  _EVAL_4423;
  wire  _EVAL_4424;
  wire  _EVAL_4427;
  wire  _EVAL_4428;
  wire  _EVAL_4429;
  wire  _EVAL_4430;
  wire  _EVAL_4431;
  wire  _EVAL_4432;
  wire  _EVAL_4433;
  wire  _EVAL_4434;
  wire  _EVAL_4435;
  wire  _EVAL_4436;
  wire  _EVAL_4439;
  wire  _EVAL_4442;
  wire  _EVAL_4444;
  wire  _EVAL_4447;
  wire  _EVAL_4450;
  wire  _EVAL_4451;
  wire  _EVAL_4453;
  wire  _EVAL_4454;
  wire  _EVAL_4455;
  wire  _EVAL_4457;
  wire  _EVAL_4459;
  wire  _EVAL_4460;
  wire  _EVAL_4461;
  wire  _EVAL_4462;
  wire  _EVAL_4463;
  wire  _EVAL_4464;
  wire  _EVAL_4468;
  wire  _EVAL_4470;
  wire  _EVAL_4471;
  wire  _EVAL_4472;
  wire  _EVAL_4473;
  wire  _EVAL_4475;
  wire  _EVAL_4481;
  wire  _EVAL_4485;
  wire  _EVAL_4487;
  wire  _EVAL_4488;
  wire  _EVAL_4491;
  wire  _EVAL_4492;
  wire  _EVAL_4494;
  wire [6:0] _EVAL_4495;
  wire  _EVAL_4498;
  wire  _EVAL_4499;
  wire  _EVAL_4501;
  wire  _EVAL_4502;
  wire  _EVAL_4503;
  wire  _EVAL_4504;
  wire  _EVAL_4506;
  wire  _EVAL_4507;
  wire  _EVAL_4512;
  wire  _EVAL_4513;
  wire  _EVAL_4514;
  wire  _EVAL_4516;
  wire  _EVAL_4519;
  wire  _EVAL_4521;
  wire  _EVAL_4522;
  wire  _EVAL_4524;
  wire  _EVAL_4525;
  wire  _EVAL_4527;
  wire  _EVAL_4529;
  wire  _EVAL_4531;
  wire  _EVAL_4533;
  wire  _EVAL_4535;
  wire  _EVAL_4536;
  wire  _EVAL_4537;
  wire  _EVAL_4543;
  wire  _EVAL_4544;
  wire  _EVAL_4545;
  wire  _EVAL_4550;
  wire [7:0] _EVAL_4551;
  wire [7:0] _EVAL_4552;
  wire  _EVAL_4555;
  wire  _EVAL_4557;
  wire  _EVAL_4558;
  wire  _EVAL_4559;
  wire  _EVAL_4560;
  wire  _EVAL_4561;
  wire  _EVAL_4563;
  wire  _EVAL_4564;
  wire  _EVAL_4565;
  wire  _EVAL_4567;
  wire  _EVAL_4568;
  wire  _EVAL_4570;
  wire  _EVAL_4573;
  wire  _EVAL_4575;
  wire  _EVAL_4576;
  wire  _EVAL_4577;
  wire  _EVAL_4579;
  wire  _EVAL_4581;
  wire  _EVAL_4585;
  wire  _EVAL_4586;
  wire  _EVAL_4587;
  wire  _EVAL_4589;
  wire  _EVAL_4591;
  wire  _EVAL_4592;
  wire  _EVAL_4593;
  wire  _EVAL_4594;
  wire  _EVAL_4596;
  wire  _EVAL_4597;
  wire  _EVAL_4598;
  wire  _EVAL_4601;
  wire  _EVAL_4604;
  wire  _EVAL_4605;
  wire  _EVAL_4607;
  wire  _EVAL_4608;
  wire  _EVAL_4609;
  wire  _EVAL_4613;
  wire  _EVAL_4616;
  wire  _EVAL_4617;
  wire  _EVAL_4618;
  wire  _EVAL_4619;
  wire  _EVAL_4623;
  wire  _EVAL_4625;
  wire  _EVAL_4627;
  wire  _EVAL_4628;
  wire  _EVAL_4629;
  wire  _EVAL_4630;
  wire  _EVAL_4635;
  wire  _EVAL_4639;
  wire  _EVAL_4641;
  wire  _EVAL_4643;
  wire  _EVAL_4644;
  wire  _EVAL_4645;
  wire  _EVAL_4647;
  wire  _EVAL_4648;
  wire  _EVAL_4649;
  wire  _EVAL_4651;
  wire  _EVAL_4652;
  wire  _EVAL_4654;
  wire  _EVAL_4655;
  wire  _EVAL_4656;
  wire  _EVAL_4661;
  wire  _EVAL_4664;
  wire  _EVAL_4666;
  wire  _EVAL_4667;
  wire  _EVAL_4668;
  wire  _EVAL_4669;
  wire  _EVAL_4670;
  wire [3:0] _EVAL_4671;
  wire  _EVAL_4673;
  wire  _EVAL_4674;
  wire  _EVAL_4675;
  wire  _EVAL_4678;
  wire  _EVAL_4680;
  wire  _EVAL_4681;
  wire  _EVAL_4682;
  wire  _EVAL_4686;
  wire  _EVAL_4688;
  wire  _EVAL_4689;
  wire  _EVAL_4690;
  wire  _EVAL_4691;
  wire  _EVAL_4692;
  wire  _EVAL_4693;
  wire  _EVAL_4694;
  wire  _EVAL_4695;
  wire  _EVAL_4697;
  wire  _EVAL_4698;
  wire  _EVAL_4701;
  wire  _EVAL_4702;
  wire  _EVAL_4703;
  wire  _EVAL_4706;
  wire  _EVAL_4707;
  wire  _EVAL_4710;
  wire  _EVAL_4712;
  wire  _EVAL_4713;
  wire  _EVAL_4714;
  wire  _EVAL_4715;
  wire  _EVAL_4720;
  wire  _EVAL_4722;
  wire  _EVAL_4723;
  wire  _EVAL_4724;
  wire  _EVAL_4726;
  wire  _EVAL_4727;
  wire  _EVAL_4729;
  wire  _EVAL_4730;
  wire  _EVAL_4731;
  wire  _EVAL_4733;
  wire  _EVAL_4736;
  wire  _EVAL_4737;
  wire  _EVAL_4739;
  wire  _EVAL_4743;
  wire  _EVAL_4744;
  wire  _EVAL_4745;
  wire  _EVAL_4748;
  wire  _EVAL_4750;
  wire  _EVAL_4751;
  wire  _EVAL_4755;
  wire  _EVAL_4756;
  wire  _EVAL_4757;
  wire  _EVAL_4759;
  wire  _EVAL_4760;
  wire  _EVAL_4761;
  wire  _EVAL_4762;
  wire  _EVAL_4764;
  wire  _EVAL_4765;
  wire  _EVAL_4766;
  wire  _EVAL_4767;
  wire  _EVAL_4768;
  wire  _EVAL_4773;
  wire  _EVAL_4775;
  wire  _EVAL_4777;
  wire  _EVAL_4780;
  wire  _EVAL_4781;
  wire  _EVAL_4782;
  wire  _EVAL_4783;
  wire  _EVAL_4784;
  wire  _EVAL_4787;
  wire  _EVAL_4788;
  wire  _EVAL_4790;
  wire  _EVAL_4792;
  wire  _EVAL_4793;
  wire  _EVAL_4794;
  wire  _EVAL_4795;
  wire  _EVAL_4796;
  wire  _EVAL_4798;
  wire  _EVAL_4800;
  wire  _EVAL_4801;
  wire  _EVAL_4802;
  wire  _EVAL_4803;
  wire  _EVAL_4804;
  wire  _EVAL_4806;
  wire  _EVAL_4811;
  wire  _EVAL_4812;
  wire  _EVAL_4813;
  wire  _EVAL_4814;
  wire  _EVAL_4817;
  wire  _EVAL_4821;
  wire  _EVAL_4825;
  wire  _EVAL_4830;
  wire  _EVAL_4831;
  wire [3:0] _EVAL_4832;
  wire  _EVAL_4833;
  wire  _EVAL_4834;
  wire  _EVAL_4836;
  wire  _EVAL_4838;
  wire  _EVAL_4841;
  wire  _EVAL_4842;
  wire  _EVAL_4844;
  wire  _EVAL_4845;
  wire  _EVAL_4847;
  wire [7:0] _EVAL_4850;
  wire  _EVAL_4851;
  wire  _EVAL_4854;
  wire  _EVAL_4855;
  wire  _EVAL_4856;
  wire  _EVAL_4857;
  wire  _EVAL_4859;
  wire  _EVAL_4861;
  wire  _EVAL_4862;
  wire  _EVAL_4866;
  wire  _EVAL_4867;
  wire  _EVAL_4868;
  wire  _EVAL_4870;
  wire  _EVAL_4871;
  wire  _EVAL_4872;
  wire  _EVAL_4873;
  wire  _EVAL_4874;
  wire  _EVAL_4877;
  wire  _EVAL_4879;
  wire  _EVAL_4881;
  wire  _EVAL_4886;
  wire  _EVAL_4887;
  wire  _EVAL_4888;
  wire  _EVAL_4890;
  wire  _EVAL_4891;
  wire  _EVAL_4892;
  wire  _EVAL_4896;
  wire  _EVAL_4898;
  wire  _EVAL_4900;
  wire  _EVAL_4904;
  wire  _EVAL_4907;
  wire  _EVAL_4909;
  wire  _EVAL_4910;
  wire  _EVAL_4912;
  wire  _EVAL_4914;
  wire  _EVAL_4915;
  wire  _EVAL_4916;
  wire  _EVAL_4917;
  wire  _EVAL_4918;
  wire  _EVAL_4920;
  wire  _EVAL_4923;
  wire  _EVAL_4925;
  wire  _EVAL_4926;
  wire  _EVAL_4928;
  wire  _EVAL_4930;
  wire  _EVAL_4931;
  wire  _EVAL_4934;
  wire  _EVAL_4936;
  wire  _EVAL_4938;
  wire  _EVAL_4939;
  wire  _EVAL_4946;
  wire  _EVAL_4947;
  wire  _EVAL_4949;
  wire  _EVAL_4950;
  wire  _EVAL_4951;
  wire  _EVAL_4952;
  wire  _EVAL_4957;
  wire  _EVAL_4960;
  wire  _EVAL_4961;
  wire  _EVAL_4962;
  wire  _EVAL_4963;
  wire  _EVAL_4964;
  wire  _EVAL_4966;
  wire  _EVAL_4967;
  wire  _EVAL_4971;
  wire  _EVAL_4974;
  wire  _EVAL_4975;
  wire  _EVAL_4976;
  wire  _EVAL_4979;
  wire  _EVAL_4981;
  wire  _EVAL_4983;
  wire  _EVAL_4984;
  wire  _EVAL_4985;
  wire  _EVAL_4987;
  wire  _EVAL_4988;
  wire  _EVAL_4989;
  wire  _EVAL_4991;
  wire  _EVAL_4993;
  wire  _EVAL_4996;
  wire  _EVAL_4999;
  wire  _EVAL_5003;
  wire  _EVAL_5005;
  wire  _EVAL_5006;
  wire  _EVAL_5015;
  wire  _EVAL_5016;
  wire  _EVAL_5017;
  wire  _EVAL_5018;
  wire  _EVAL_5020;
  wire  _EVAL_5021;
  wire  _EVAL_5023;
  wire  _EVAL_5025;
  wire  _EVAL_5027;
  wire  _EVAL_5028;
  wire  _EVAL_5032;
  wire  _EVAL_5033;
  wire  _EVAL_5035;
  wire  _EVAL_5036;
  wire  _EVAL_5037;
  wire  _EVAL_5040;
  wire  _EVAL_5042;
  wire  _EVAL_5043;
  wire  _EVAL_5050;
  wire  _EVAL_5051;
  wire  _EVAL_5053;
  wire  _EVAL_5054;
  wire  _EVAL_5055;
  wire  _EVAL_5056;
  wire  _EVAL_5057;
  wire  _EVAL_5059;
  wire  _EVAL_5060;
  wire  _EVAL_5063;
  wire  _EVAL_5066;
  wire  _EVAL_5067;
  wire  _EVAL_5069;
  wire  _EVAL_5071;
  wire  _EVAL_5072;
  wire  _EVAL_5074;
  wire  _EVAL_5075;
  wire  _EVAL_5076;
  wire  _EVAL_5077;
  wire  _EVAL_5078;
  wire  _EVAL_5079;
  wire  _EVAL_5081;
  wire  _EVAL_5082;
  wire  _EVAL_5083;
  wire  _EVAL_5084;
  wire  _EVAL_5085;
  wire  _EVAL_5087;
  wire  _EVAL_5088;
  wire  _EVAL_5090;
  wire  _EVAL_5091;
  wire  _EVAL_5092;
  wire  _EVAL_5094;
  wire  _EVAL_5099;
  wire  _EVAL_5100;
  wire  _EVAL_5102;
  wire  _EVAL_5103;
  wire  _EVAL_5105;
  wire  _EVAL_5110;
  wire  _EVAL_5114;
  wire  _EVAL_5116;
  wire  _EVAL_5118;
  wire  _EVAL_5119;
  wire  _EVAL_5121;
  wire  _EVAL_5122;
  wire  _EVAL_5123;
  wire  _EVAL_5124;
  wire  _EVAL_5127;
  wire  _EVAL_5128;
  wire  _EVAL_5129;
  wire  _EVAL_5130;
  wire  _EVAL_5132;
  wire  _EVAL_5133;
  wire  _EVAL_5134;
  wire  _EVAL_5135;
  wire  _EVAL_5136;
  wire  _EVAL_5138;
  wire  _EVAL_5141;
  wire  _EVAL_5144;
  wire  _EVAL_5148;
  wire  _EVAL_5149;
  wire  _EVAL_5152;
  wire  _EVAL_5153;
  wire  _EVAL_5155;
  wire  _EVAL_5157;
  wire  _EVAL_5158;
  wire  _EVAL_5159;
  wire  _EVAL_5160;
  wire  _EVAL_5161;
  wire  _EVAL_5162;
  wire  _EVAL_5167;
  wire  _EVAL_5170;
  wire  _EVAL_5173;
  wire  _EVAL_5175;
  wire  _EVAL_5177;
  wire  _EVAL_5178;
  wire  _EVAL_5179;
  wire  _EVAL_5182;
  wire  _EVAL_5184;
  wire  _EVAL_5187;
  wire  _EVAL_5189;
  wire  _EVAL_5192;
  wire  _EVAL_5193;
  wire  _EVAL_5194;
  wire  _EVAL_5196;
  wire  _EVAL_5199;
  wire  _EVAL_5200;
  wire  _EVAL_5201;
  wire  _EVAL_5205;
  wire  _EVAL_5206;
  wire  _EVAL_5207;
  wire  _EVAL_5208;
  wire  _EVAL_5209;
  wire  _EVAL_5210;
  wire  _EVAL_5211;
  wire  _EVAL_5212;
  wire  _EVAL_5213;
  wire  _EVAL_5214;
  wire  _EVAL_5215;
  wire  _EVAL_5216;
  wire  _EVAL_5217;
  wire  _EVAL_5218;
  wire  _EVAL_5219;
  wire  _EVAL_5223;
  wire  _EVAL_5226;
  wire  _EVAL_5228;
  wire  _EVAL_5229;
  wire  _EVAL_5230;
  wire  _EVAL_5233;
  wire  _EVAL_5234;
  wire  _EVAL_5235;
  wire  _EVAL_5236;
  wire  _EVAL_5238;
  wire  _EVAL_5239;
  wire  _EVAL_5240;
  wire  _EVAL_5241;
  wire  _EVAL_5242;
  wire  _EVAL_5243;
  wire  _EVAL_5245;
  wire  _EVAL_5246;
  wire  _EVAL_5250;
  wire  _EVAL_5251;
  wire  _EVAL_5252;
  wire  _EVAL_5259;
  wire  _EVAL_5260;
  wire  _EVAL_5261;
  wire  _EVAL_5264;
  wire  _EVAL_5268;
  wire  _EVAL_5271;
  wire  _EVAL_5272;
  wire  _EVAL_5273;
  wire  _EVAL_5274;
  wire  _EVAL_5276;
  wire  _EVAL_5277;
  wire  _EVAL_5280;
  wire  _EVAL_5281;
  wire  _EVAL_5282;
  wire  _EVAL_5283;
  wire  _EVAL_5284;
  wire  _EVAL_5285;
  wire  _EVAL_5286;
  wire  _EVAL_5289;
  wire  _EVAL_5291;
  wire  _EVAL_5292;
  wire  _EVAL_5296;
  wire  _EVAL_5298;
  wire  _EVAL_5299;
  wire  _EVAL_5302;
  wire  _EVAL_5303;
  wire  _EVAL_5304;
  wire  _EVAL_5305;
  wire  _EVAL_5306;
  wire  _EVAL_5308;
  wire  _EVAL_5310;
  wire  _EVAL_5313;
  wire  _EVAL_5316;
  wire  _EVAL_5317;
  wire  _EVAL_5319;
  wire  _EVAL_5320;
  wire  _EVAL_5327;
  wire  _EVAL_5328;
  wire  _EVAL_5329;
  wire  _EVAL_5336;
  wire  _EVAL_5338;
  wire  _EVAL_5341;
  wire  _EVAL_5342;
  wire  _EVAL_5343;
  wire  _EVAL_5344;
  wire  _EVAL_5347;
  wire  _EVAL_5349;
  wire  _EVAL_5351;
  wire  _EVAL_5352;
  wire  _EVAL_5353;
  wire  _EVAL_5354;
  wire  _EVAL_5355;
  wire  _EVAL_5356;
  wire  _EVAL_5357;
  wire  _EVAL_5360;
  wire  _EVAL_5361;
  wire  _EVAL_5362;
  wire  _EVAL_5365;
  wire  _EVAL_5367;
  wire  _EVAL_5368;
  wire  _EVAL_5370;
  wire  _EVAL_5371;
  wire  _EVAL_5372;
  wire  _EVAL_5376;
  wire  _EVAL_5379;
  wire  _EVAL_5380;
  wire  _EVAL_5381;
  wire  _EVAL_5383;
  wire  _EVAL_5385;
  wire  _EVAL_5387;
  wire  _EVAL_5395;
  wire  _EVAL_5398;
  wire  _EVAL_5400;
  wire  _EVAL_5401;
  wire  _EVAL_5402;
  wire  _EVAL_5404;
  wire  _EVAL_5408;
  wire  _EVAL_5412;
  wire  _EVAL_5414;
  wire  _EVAL_5416;
  wire  _EVAL_5417;
  wire  _EVAL_5418;
  wire  _EVAL_5419;
  wire  _EVAL_5420;
  wire  _EVAL_5422;
  wire  _EVAL_5423;
  wire  _EVAL_5424;
  wire  _EVAL_5425;
  wire  _EVAL_5427;
  wire  _EVAL_5428;
  wire  _EVAL_5430;
  wire  _EVAL_5431;
  wire  _EVAL_5433;
  wire  _EVAL_5434;
  wire  _EVAL_5437;
  wire  _EVAL_5438;
  wire  _EVAL_5439;
  wire  _EVAL_5440;
  wire  _EVAL_5443;
  wire  _EVAL_5444;
  wire  _EVAL_5445;
  wire  _EVAL_5446;
  wire  _EVAL_5447;
  wire  _EVAL_5449;
  wire  _EVAL_5450;
  wire  _EVAL_5451;
  wire  _EVAL_5452;
  wire  _EVAL_5454;
  wire  _EVAL_5455;
  wire  _EVAL_5456;
  wire  _EVAL_5457;
  wire  _EVAL_5458;
  wire  _EVAL_5461;
  wire  _EVAL_5464;
  wire  _EVAL_5465;
  wire  _EVAL_5466;
  wire  _EVAL_5470;
  wire  _EVAL_5471;
  wire  _EVAL_5473;
  wire  _EVAL_5474;
  wire  _EVAL_5476;
  wire  _EVAL_5477;
  wire  _EVAL_5478;
  wire  _EVAL_5482;
  wire  _EVAL_5483;
  wire  _EVAL_5486;
  wire  _EVAL_5488;
  wire  _EVAL_5489;
  wire  _EVAL_5490;
  wire  _EVAL_5492;
  wire  _EVAL_5493;
  wire  _EVAL_5496;
  wire  _EVAL_5497;
  wire  _EVAL_5498;
  wire  _EVAL_5500;
  wire  _EVAL_5502;
  wire  _EVAL_5507;
  wire  _EVAL_5508;
  wire  _EVAL_5509;
  wire  _EVAL_5510;
  wire  _EVAL_5512;
  wire  _EVAL_5514;
  wire  _EVAL_5517;
  wire  _EVAL_5524;
  wire  _EVAL_5525;
  wire  _EVAL_5527;
  wire  _EVAL_5528;
  wire  _EVAL_5529;
  wire  _EVAL_5530;
  wire  _EVAL_5531;
  wire  _EVAL_5532;
  wire  _EVAL_5534;
  wire  _EVAL_5538;
  wire  _EVAL_5541;
  wire  _EVAL_5542;
  wire  _EVAL_5543;
  wire  _EVAL_5544;
  wire  _EVAL_5549;
  wire  _EVAL_5559;
  wire  _EVAL_5560;
  wire  _EVAL_5561;
  wire  _EVAL_5564;
  wire  _EVAL_5565;
  wire  _EVAL_5566;
  wire  _EVAL_5568;
  wire  _EVAL_5569;
  wire  _EVAL_5570;
  wire  _EVAL_5573;
  wire  _EVAL_5574;
  wire  _EVAL_5575;
  wire  _EVAL_5576;
  wire  _EVAL_5578;
  wire  _EVAL_5583;
  wire  _EVAL_5586;
  wire  _EVAL_5587;
  wire  _EVAL_5588;
  wire  _EVAL_5589;
  wire  _EVAL_5590;
  wire  _EVAL_5592;
  wire  _EVAL_5593;
  wire  _EVAL_5594;
  wire  _EVAL_5596;
  wire  _EVAL_5598;
  wire  _EVAL_5599;
  wire  _EVAL_5601;
  wire  _EVAL_5602;
  wire  _EVAL_5604;
  wire  _EVAL_5607;
  wire  _EVAL_5610;
  wire  _EVAL_5613;
  wire  _EVAL_5616;
  wire  _EVAL_5618;
  wire  _EVAL_5620;
  wire  _EVAL_5622;
  wire  _EVAL_5625;
  wire  _EVAL_5630;
  wire  _EVAL_5631;
  wire  _EVAL_5632;
  wire  _EVAL_5633;
  wire  _EVAL_5634;
  wire  _EVAL_5639;
  wire  _EVAL_5640;
  wire  _EVAL_5641;
  wire  _EVAL_5642;
  wire  _EVAL_5643;
  wire  _EVAL_5647;
  wire  _EVAL_5648;
  wire  _EVAL_5649;
  wire  _EVAL_5650;
  wire  _EVAL_5651;
  wire  _EVAL_5652;
  wire  _EVAL_5654;
  wire  _EVAL_5656;
  wire  _EVAL_5659;
  wire  _EVAL_5662;
  wire  _EVAL_5663;
  wire  _EVAL_5664;
  wire  _EVAL_5666;
  wire  _EVAL_5668;
  wire  _EVAL_5671;
  wire  _EVAL_5672;
  wire  _EVAL_5673;
  wire  _EVAL_5676;
  wire  _EVAL_5678;
  wire  _EVAL_5679;
  wire  _EVAL_5680;
  wire  _EVAL_5685;
  wire  _EVAL_5686;
  wire  _EVAL_5688;
  wire  _EVAL_5692;
  wire  _EVAL_5693;
  wire  _EVAL_5695;
  wire  _EVAL_5700;
  wire  _EVAL_5702;
  wire  _EVAL_5703;
  wire  _EVAL_5704;
  wire  _EVAL_5705;
  wire  _EVAL_5707;
  wire  _EVAL_5708;
  wire  _EVAL_5720;
  wire  _EVAL_5721;
  wire  _EVAL_5722;
  wire  _EVAL_5723;
  wire  _EVAL_5724;
  wire  _EVAL_5726;
  wire  _EVAL_5729;
  wire  _EVAL_5733;
  wire  _EVAL_5734;
  wire  _EVAL_5736;
  wire  _EVAL_5737;
  wire  _EVAL_5739;
  wire  _EVAL_5740;
  wire  _EVAL_5744;
  wire  _EVAL_5747;
  wire  _EVAL_5750;
  wire  _EVAL_5752;
  wire  _EVAL_5753;
  wire  _EVAL_5754;
  wire  _EVAL_5755;
  wire  _EVAL_5756;
  wire  _EVAL_5760;
  wire  _EVAL_5761;
  wire  _EVAL_5764;
  wire  _EVAL_5766;
  wire  _EVAL_5772;
  wire  _EVAL_5773;
  wire  _EVAL_5774;
  wire  _EVAL_5775;
  wire  _EVAL_5776;
  wire  _EVAL_5778;
  wire  _EVAL_5779;
  wire  _EVAL_5784;
  wire  _EVAL_5786;
  wire  _EVAL_5788;
  wire  _EVAL_5789;
  wire  _EVAL_5790;
  wire  _EVAL_5795;
  wire  _EVAL_5796;
  wire  _EVAL_5797;
  wire  _EVAL_5798;
  wire  _EVAL_5809;
  wire  _EVAL_5810;
  wire  _EVAL_5811;
  wire  _EVAL_5812;
  wire  _EVAL_5814;
  wire  _EVAL_5816;
  wire  _EVAL_5819;
  wire  _EVAL_5822;
  wire  _EVAL_5823;
  wire  _EVAL_5825;
  wire  _EVAL_5826;
  wire  _EVAL_5827;
  wire  _EVAL_5831;
  wire  _EVAL_5832;
  wire  _EVAL_5834;
  wire  _EVAL_5837;
  wire  _EVAL_5838;
  wire  _EVAL_5839;
  wire  _EVAL_5840;
  wire  _EVAL_5842;
  wire  _EVAL_5843;
  wire  _EVAL_5845;
  wire  _EVAL_5848;
  wire  _EVAL_5850;
  wire  _EVAL_5853;
  wire  _EVAL_5854;
  wire  _EVAL_5855;
  wire  _EVAL_5856;
  wire  _EVAL_5857;
  wire  _EVAL_5858;
  wire  _EVAL_5866;
  wire  _EVAL_5867;
  wire  _EVAL_5868;
  wire  _EVAL_5869;
  wire  _EVAL_5874;
  wire  _EVAL_5877;
  wire  _EVAL_5879;
  wire  _EVAL_5880;
  wire  _EVAL_5882;
  wire  _EVAL_5886;
  wire  _EVAL_5887;
  wire  _EVAL_5888;
  wire  _EVAL_5889;
  wire  _EVAL_5892;
  wire  _EVAL_5893;
  wire  _EVAL_5895;
  wire  _EVAL_5896;
  wire  _EVAL_5897;
  wire  _EVAL_5900;
  wire  _EVAL_5902;
  wire  _EVAL_5904;
  wire  _EVAL_5911;
  wire  _EVAL_5912;
  wire  _EVAL_5914;
  wire  _EVAL_5917;
  wire  _EVAL_5919;
  wire  _EVAL_5920;
  wire  _EVAL_5921;
  wire [3:0] _EVAL_5922;
  wire  _EVAL_5927;
  wire  _EVAL_5930;
  wire  _EVAL_5932;
  wire  _EVAL_5936;
  wire  _EVAL_5937;
  wire  _EVAL_5938;
  wire  _EVAL_5941;
  wire  _EVAL_5943;
  wire  _EVAL_5945;
  wire  _EVAL_5946;
  wire  _EVAL_5947;
  wire  _EVAL_5948;
  wire  _EVAL_5950;
  wire  _EVAL_5953;
  wire  _EVAL_5954;
  wire  _EVAL_5955;
  wire  _EVAL_5956;
  wire  _EVAL_5959;
  wire  _EVAL_5964;
  wire  _EVAL_5968;
  wire  _EVAL_5970;
  wire  _EVAL_5971;
  wire  _EVAL_5973;
  wire  _EVAL_5974;
  wire  _EVAL_5975;
  wire  _EVAL_5976;
  wire  _EVAL_5977;
  wire  _EVAL_5978;
  wire  _EVAL_5979;
  wire  _EVAL_5980;
  wire  _EVAL_5982;
  wire  _EVAL_5986;
  wire  _EVAL_5987;
  wire  _EVAL_5988;
  wire  _EVAL_5990;
  wire  _EVAL_5991;
  wire  _EVAL_5992;
  wire  _EVAL_5994;
  wire  _EVAL_5998;
  wire  _EVAL_5999;
  wire  _EVAL_6001;
  wire  _EVAL_6002;
  wire  _EVAL_6003;
  wire  _EVAL_6005;
  wire  _EVAL_6007;
  wire  _EVAL_6008;
  wire  _EVAL_6010;
  wire  _EVAL_6011;
  wire  _EVAL_6015;
  wire  _EVAL_6017;
  wire  _EVAL_6022;
  wire  _EVAL_6024;
  wire  _EVAL_6026;
  wire  _EVAL_6029;
  wire  _EVAL_6032;
  wire  _EVAL_6033;
  wire  _EVAL_6036;
  wire  _EVAL_6037;
  wire  _EVAL_6038;
  wire  _EVAL_6039;
  wire  _EVAL_6045;
  wire  _EVAL_6047;
  wire  _EVAL_6048;
  wire  _EVAL_6050;
  wire  _EVAL_6051;
  wire  _EVAL_6054;
  wire  _EVAL_6055;
  wire  _EVAL_6057;
  wire  _EVAL_6059;
  wire  _EVAL_6062;
  wire  _EVAL_6065;
  wire  _EVAL_6068;
  wire  _EVAL_6069;
  wire  _EVAL_6070;
  wire  _EVAL_6075;
  wire  _EVAL_6076;
  wire  _EVAL_6077;
  wire  _EVAL_6080;
  wire  _EVAL_6083;
  wire  _EVAL_6084;
  wire  _EVAL_6085;
  wire  _EVAL_6086;
  wire  _EVAL_6087;
  wire [30:0] _EVAL_6088;
  wire  _EVAL_6089;
  wire  _EVAL_6090;
  wire  _EVAL_6093;
  wire  _EVAL_6094;
  wire  _EVAL_6095;
  wire  _EVAL_6096;
  wire  _EVAL_6097;
  wire  _EVAL_6099;
  wire  _EVAL_6102;
  _EVAL_114_assert TLMonitor (
    ._EVAL(TLMonitor__EVAL),
    ._EVAL_0(TLMonitor__EVAL_0),
    ._EVAL_1(TLMonitor__EVAL_1),
    ._EVAL_2(TLMonitor__EVAL_2),
    ._EVAL_3(TLMonitor__EVAL_3),
    ._EVAL_4(TLMonitor__EVAL_4),
    ._EVAL_5(TLMonitor__EVAL_5),
    ._EVAL_6(TLMonitor__EVAL_6),
    ._EVAL_7(TLMonitor__EVAL_7),
    ._EVAL_8(TLMonitor__EVAL_8),
    ._EVAL_9(TLMonitor__EVAL_9),
    ._EVAL_10(TLMonitor__EVAL_10),
    ._EVAL_11(TLMonitor__EVAL_11),
    ._EVAL_12(TLMonitor__EVAL_12),
    ._EVAL_13(TLMonitor__EVAL_13),
    ._EVAL_14(TLMonitor__EVAL_14)
  );
  assign _EVAL_2258 = ~_EVAL_4738;
  assign _EVAL_1449 = _EVAL_3639 & _EVAL_5211;
  assign _EVAL_596 = _EVAL_3524 & _EVAL_5543;
  assign _EVAL_5994 = _EVAL_4134 & _EVAL_673;
  assign _EVAL_1299 = _EVAL_1145[582];
  assign _EVAL_4129 = _EVAL_5478 & _EVAL_3398;
  assign _EVAL_3101 = _EVAL_4843 & _EVAL_2921;
  assign _EVAL_1568 = _EVAL_1242 & _EVAL_3418;
  assign _EVAL_3143 = _EVAL_5132 & _EVAL_847;
  assign _EVAL_242 = _EVAL_5816 & _EVAL_3508;
  assign _EVAL_5943 = _EVAL_4707 & _EVAL_3766;
  assign _EVAL_479 = _EVAL_3801 & _EVAL_3379;
  assign _EVAL_247 = _EVAL_961 & _EVAL_5543;
  assign _EVAL_3531 = _EVAL_2471 & _EVAL_3154;
  assign _EVAL_5032 = _EVAL_4372 & _EVAL_3702;
  assign _EVAL_2977 = _EVAL_5998 & _EVAL_3170;
  assign _EVAL_4208 = _EVAL_386 & _EVAL_2748;
  assign _EVAL_2424 = _EVAL_3321 != 7'h0;
  assign _EVAL_5118 = _EVAL_3859 & _EVAL_1198;
  assign _EVAL_208 = ~_EVAL_3594;
  assign _EVAL_3038 = _EVAL_1145[670];
  assign _EVAL_3013 = _EVAL_1675 & _EVAL_369;
  assign _EVAL_1051 = _EVAL_4627 & _EVAL_4564;
  assign _EVAL_6068 = _EVAL_1158 & _EVAL_882;
  assign _EVAL_3981 = _EVAL_4831 & _EVAL_673;
  assign _EVAL_2095 = _EVAL_2454 & _EVAL_3170;
  assign _EVAL_3314 = _EVAL_4627 & _EVAL_5937;
  assign _EVAL_1185 = ~_EVAL_1245;
  assign _EVAL_909 = _EVAL_4567 & _EVAL_882;
  assign _EVAL_5632 = _EVAL_1553 & _EVAL_1009;
  assign _EVAL_5695 = _EVAL_3845 & _EVAL_1198;
  assign _EVAL_3628 = _EVAL_5353 & _EVAL_2424;
  assign _EVAL_2412 = _EVAL_5063 & _EVAL_3261;
  assign _EVAL_5721 = _EVAL_2170 & _EVAL_6084;
  assign _EVAL_2441 = _EVAL_4374 & _EVAL_208;
  assign _EVAL_1651 = _EVAL_3156 & _EVAL_2748;
  assign _EVAL_5138 = _EVAL_6075 & _EVAL_3418;
  assign _EVAL_5622 = _EVAL_4525 & _EVAL_1735;
  assign _EVAL_4288 = _EVAL_4987 & _EVAL_1198;
  assign _EVAL_5361 = _EVAL_1242 & _EVAL_882;
  assign _EVAL_3807 = _EVAL_1145[675];
  assign _EVAL_931 = _EVAL_1145[641];
  assign _EVAL_1294 = _EVAL_984 & _EVAL_2956;
  assign _EVAL_6095 = _EVAL_3082 & _EVAL_369;
  assign _EVAL_5489 = _EVAL_4093 & _EVAL_882;
  assign _EVAL_5496 = ~_EVAL_2993;
  assign _EVAL_5371 = _EVAL_3920 & _EVAL_587;
  assign _EVAL_4928 = _EVAL_5994 & _EVAL_3398;
  assign _EVAL_482 = _EVAL_2868 & _EVAL_3398;
  assign _EVAL_2327 = _EVAL_5074 & _EVAL_2975;
  assign _EVAL_4341 = _EVAL_1145[595];
  assign _EVAL_3991 = _EVAL_774 & _EVAL_3702;
  assign _EVAL_1819 = _EVAL_3993 & _EVAL_3418;
  assign _EVAL_1405 = _EVAL_3710 & _EVAL_2969;
  assign _EVAL_223 = _EVAL_5450 & _EVAL_3170;
  assign _EVAL_217 = _EVAL_1542 & _EVAL_3261;
  assign _EVAL_875 = _EVAL_5662 & _EVAL_847;
  assign _EVAL_721 = _EVAL_4200 & _EVAL_3261;
  assign _EVAL_3548 = ~_EVAL_1942;
  assign _EVAL_3249 = _EVAL_1211 & _EVAL_256;
  assign _EVAL_4144 = _EVAL_2569 & _EVAL_3379;
  assign _EVAL_5158 = ~_EVAL_3001;
  assign _EVAL_4462 = _EVAL_6089 & _EVAL_673;
  assign _EVAL_3401 = _EVAL_4916 & _EVAL_5850;
  assign _EVAL_4201 = _EVAL_4200 & _EVAL_3398;
  assign _EVAL_358 = _EVAL_5344 & _EVAL_2382;
  assign _EVAL_2358 = _EVAL_538 & _EVAL_3702;
  assign _EVAL_2539 = _EVAL_4550 & _EVAL_5543;
  assign _EVAL_3183 = _EVAL_2419 & _EVAL_3379;
  assign _EVAL_3780 = _EVAL_4916 & _EVAL_1735;
  assign _EVAL_4084 = _EVAL_4627 & _EVAL_2609;
  assign _EVAL_2038 = _EVAL_5074 & _EVAL_4154;
  assign _EVAL_3969 = _EVAL_3815 & _EVAL_2382;
  assign _EVAL_3473 = _EVAL_3710 & _EVAL_2424;
  assign _EVAL_3734 = _EVAL_3689 & _EVAL_5543;
  assign _EVAL_4385 = _EVAL_504 & _EVAL_2956;
  assign _EVAL_2909 = _EVAL_3216 & _EVAL_3261;
  assign _EVAL_6050 = _EVAL_6059 & _EVAL_3154;
  assign _EVAL_3842 = _EVAL_4488 & _EVAL_847;
  assign _EVAL_1365 = _EVAL_263 & _EVAL_2956;
  assign _EVAL_3631 = _EVAL_905 & _EVAL_847;
  assign _EVAL_1702 = _EVAL_407 & _EVAL_3702;
  assign _EVAL_2624 = _EVAL_529 & _EVAL_5299;
  assign _EVAL_2772 = _EVAL_5074 & _EVAL_2609;
  assign _EVAL_6062 = _EVAL_3845 & _EVAL_3284;
  assign _EVAL_5450 = _EVAL_2676 & _EVAL_3379;
  assign _EVAL_869 = _EVAL_4627 & _EVAL_4408;
  assign _EVAL_2028 = _EVAL_5246 & _EVAL_3398;
  assign _EVAL_4591 = _EVAL_284 & _EVAL_6084;
  assign _EVAL_5560 = _EVAL_751 & _EVAL_1488;
  assign _EVAL_6045 = _EVAL_2907 & _EVAL_2424;
  assign _EVAL_442 = _EVAL_5028 & _EVAL_1735;
  assign _EVAL_365 = _EVAL_1370 & _EVAL_882;
  assign _EVAL_4481 = _EVAL_504 & _EVAL_3284;
  assign _EVAL_5920 = _EVAL_5676 & _EVAL_3398;
  assign _EVAL_2384 = _EVAL_2907 & _EVAL_2748;
  assign _EVAL_4536 = ~_EVAL_1929;
  assign _EVAL_1485 = _EVAL_751 & _EVAL_2748;
  assign _EVAL_5457 = _EVAL_2907 & _EVAL_2969;
  assign _EVAL_2320 = _EVAL_4551 != 8'h0;
  assign _EVAL_885 = _EVAL_1145[602];
  assign _EVAL_1694 = _EVAL_5705 & _EVAL_369;
  assign _EVAL_4950 = _EVAL_3689 & _EVAL_2969;
  assign _EVAL_2807 = _EVAL_3651 & _EVAL_2748;
  assign _EVAL_1039 = _EVAL_1099 & _EVAL_673;
  assign _EVAL_1038 = _EVAL_1745 & _EVAL_5464;
  assign _EVAL_5182 = _EVAL_5427 & _EVAL_3154;
  assign _EVAL_1197 = _EVAL_4689 & _EVAL_3170;
  assign _EVAL_2382 = _EVAL_3586 != 4'h0;
  assign _EVAL_3232 = _EVAL_5561 & _EVAL_5173;
  assign _EVAL_4381 = _EVAL_4311 & _EVAL_4775;
  assign _EVAL_4727 = _EVAL_5561 & _EVAL_2817;
  assign _EVAL_4886 = _EVAL_4783 & _EVAL_2969;
  assign _EVAL_2564 = _EVAL_5074 & _EVAL_5837;
  assign _EVAL_1242 = _EVAL_1063 & _EVAL_673;
  assign _EVAL_5867 = _EVAL_1145[0];
  assign _EVAL_1291 = _EVAL_961 & _EVAL_2424;
  assign _EVAL_4535 = _EVAL_1731 != 2'h0;
  assign _EVAL_1043 = _EVAL_1125 & _EVAL_882;
  assign _EVAL_955 = _EVAL_5398 & _EVAL_2969;
  assign _EVAL_4034 = _EVAL_407 & _EVAL_6084;
  assign _EVAL_5207 = _EVAL_1500 & _EVAL_3487;
  assign _EVAL_797 = _EVAL_5370 & _EVAL_3702;
  assign _EVAL_900 = _EVAL_4093 & _EVAL_847;
  assign _EVAL_2849 = _EVAL_1158 & _EVAL_3418;
  assign _EVAL_4309 = _EVAL_386 & _EVAL_1488;
  assign _EVAL_4457 = _EVAL_3052 & _EVAL_847;
  assign _EVAL_2051 = _EVAL_4661 & _EVAL_1009;
  assign _EVAL_2270 = _EVAL_1876 & _EVAL_3154;
  assign _EVAL_3583 = ~_EVAL_5101;
  assign _EVAL_5649 = _EVAL_4755 & _EVAL_1735;
  assign _EVAL_2494 = _EVAL_1854 & _EVAL_3261;
  assign _EVAL_3188 = _EVAL_4120 & _EVAL_673;
  assign _EVAL_254 = _EVAL_3996 & _EVAL_587;
  assign _EVAL_3352 = _EVAL_1145[530];
  assign _EVAL_904 = ~_EVAL_2580;
  assign _EVAL_532 = _EVAL_5561 & _EVAL_5115;
  assign _EVAL_5704 = _EVAL_5074 & _EVAL_3701;
  assign _EVAL_3136 = _EVAL_949 ? 8'hff : 8'h0;
  assign _EVAL_1010 = _EVAL_6032 & _EVAL_2969;
  assign _EVAL_1418 = _EVAL_5074 & _EVAL_2465;
  assign _EVAL_935 = _EVAL_5157 & _EVAL_3379;
  assign _EVAL_5212 = _EVAL_1649 & _EVAL_1488;
  assign _EVAL_4618 = _EVAL_1729 & _EVAL_673;
  assign _EVAL_2419 = _EVAL_5074 & _EVAL_5236;
  assign _EVAL_4694 = _EVAL_3981 & _EVAL_3418;
  assign _EVAL_2505 = _EVAL_5074 & _EVAL_3761;
  assign _EVAL_3313 = _EVAL_3058 != 8'h0;
  assign _EVAL_3942 = _EVAL_2338 & _EVAL_3702;
  assign _EVAL_2574 = _EVAL_5193 & _EVAL_2748;
  assign _EVAL_2121 = _EVAL_1254 & _EVAL_673;
  assign _EVAL_870 = _EVAL_4175 & _EVAL_3418;
  assign _EVAL_1616 = _EVAL_2550 & _EVAL_3766;
  assign _EVAL_2241 = _EVAL_4269 & _EVAL_3379;
  assign _EVAL_4936 = _EVAL_4627 & _EVAL_5936;
  assign _EVAL_5272 = _EVAL_751 & _EVAL_6084;
  assign _EVAL_2458 = _EVAL_5994 & _EVAL_882;
  assign _EVAL_914 = _EVAL_4222 & _EVAL_3398;
  assign _EVAL_354 = ~_EVAL_4398;
  assign _EVAL_2601 = _EVAL_1145[579];
  assign _EVAL_5425 = _EVAL_4525 & _EVAL_3170;
  assign _EVAL_920 = _EVAL_3935 & _EVAL_2424;
  assign _EVAL_2431 = _EVAL_2793 & _EVAL_3261;
  assign _EVAL_4668 = _EVAL_5561 & _EVAL_5405;
  assign _EVAL_4487 = _EVAL_5148 & _EVAL_6084;
  assign _EVAL_1277 = ~_EVAL_4732;
  assign _EVAL_2404 = _EVAL_3216 & _EVAL_3418;
  assign _EVAL_5282 = _EVAL_5676 & _EVAL_3154;
  assign _EVAL_4760 = _EVAL_4604 & _EVAL_1009;
  assign _EVAL_441 = _EVAL_4322 & _EVAL_369;
  assign _EVAL_2672 = _EVAL_4567 & _EVAL_3261;
  assign _EVAL_5094 = _EVAL_6080 & _EVAL_3170;
  assign _EVAL_1896 = _EVAL_4745 & _EVAL_3261;
  assign _EVAL_5242 = _EVAL_4627 & _EVAL_1299;
  assign _EVAL_4269 = _EVAL_4627 & _EVAL_4097;
  assign _EVAL_1989 = _EVAL_1316[7:1];
  assign _EVAL_3509 = _EVAL_1145[599];
  assign _EVAL_1173 = _EVAL_5068[543];
  assign _EVAL_2957 = _EVAL_3202 & _EVAL_2748;
  assign _EVAL_3162 = _EVAL_6075 & _EVAL_3154;
  assign _EVAL_4923 = _EVAL_1865 & _EVAL_3154;
  assign _EVAL_5428 = _EVAL_3183 & _EVAL_369;
  assign _EVAL_4430 = _EVAL_5561 & _EVAL_2952;
  assign _EVAL_1846 = _EVAL_4627 & _EVAL_5236;
  assign _EVAL_5703 = _EVAL_5193 & _EVAL_3702;
  assign _EVAL_2335 = _EVAL_3242 & _EVAL_3379;
  assign _EVAL_5178 = _EVAL_4224 & _EVAL_2382;
  assign _EVAL_5473 = _EVAL_284 & _EVAL_3702;
  assign _EVAL_6037 = _EVAL_3070 & _EVAL_1198;
  assign _EVAL_328 = ~_EVAL_1602;
  assign _EVAL_5177 = ~_EVAL_507;
  assign _EVAL_1555 = ~_EVAL_2162;
  assign _EVAL_4804 = _EVAL_735 & _EVAL_5464;
  assign _EVAL_2689 = _EVAL_2251 & _EVAL_2424;
  assign _EVAL_1001 = _EVAL_2616 & _EVAL_1029;
  assign _EVAL_4273 = _EVAL_6075 & _EVAL_4477;
  assign _EVAL_5349 = _EVAL_2877 & _EVAL_6084;
  assign _EVAL_2097 = _EVAL_5642 & _EVAL_3702;
  assign _EVAL_1978 = _EVAL_4311 & _EVAL_4664;
  assign _EVAL_1591 = _EVAL_1242 & _EVAL_3261;
  assign _EVAL_4939 = _EVAL_5074 & _EVAL_4564;
  assign _EVAL_4183 = _EVAL_1149 & _EVAL_2748;
  assign _EVAL_470 = _EVAL_5662 & _EVAL_882;
  assign _EVAL_3982 = _EVAL_5561 & _EVAL_4441;
  assign _EVAL_5978 = _EVAL_5618 & _EVAL_2748;
  assign _EVAL_3495 = _EVAL_3220 & _EVAL_6084;
  assign _EVAL_6033 = _EVAL_1389 & _EVAL_673;
  assign _EVAL_2704 = _EVAL_5930 & _EVAL_2969;
  assign _EVAL_4155 = _EVAL_4974 & _EVAL_1735;
  assign _EVAL_1920 = _EVAL_3596 & _EVAL_673;
  assign _EVAL_3760 = _EVAL_1536 & _EVAL_2969;
  assign _EVAL_714 = ~_EVAL_3133;
  assign _EVAL_1223 = _EVAL_5704 & _EVAL_3379;
  assign _EVAL_5427 = _EVAL_3982 & _EVAL_673;
  assign _EVAL_3014 = _EVAL_2631 & _EVAL_3418;
  assign _EVAL_5932 = _EVAL_1145[609];
  assign _EVAL_5076 = _EVAL_897 & _EVAL_1198;
  assign _EVAL_6102 = _EVAL_2100 & _EVAL_847;
  assign _EVAL_583 = _EVAL_5192 & _EVAL_2748;
  assign _EVAL_4463 = _EVAL_2100 & _EVAL_3398;
  assign _EVAL_3943 = _EVAL_4692 & _EVAL_882;
  assign _EVAL_1004 = _EVAL_5795 & _EVAL_3766;
  assign _EVAL_3769 = _EVAL_1149 & _EVAL_3702;
  assign _EVAL_800 = ~_EVAL_5985;
  assign _EVAL_2793 = _EVAL_2570 & _EVAL_673;
  assign _EVAL_3690 = _EVAL_1314 & _EVAL_5177;
  assign _EVAL_3714 = _EVAL_1149 & _EVAL_6084;
  assign _EVAL_5451 = _EVAL_2631 & _EVAL_3261;
  assign _EVAL_4575 = _EVAL_897 & _EVAL_3284;
  assign _EVAL_5464 = _EVAL_2688 != 4'h0;
  assign _EVAL_4185 = _EVAL_4224 & _EVAL_4108;
  assign _EVAL_3457 = _EVAL_921 & _EVAL_3418;
  assign _EVAL_3572 = _EVAL_446 & _EVAL_5299;
  assign _EVAL_1015 = _EVAL_1344 & _EVAL_3487;
  assign _EVAL_5671 = _EVAL_263 & _EVAL_3284;
  assign _EVAL_2652 = _EVAL_4856 & _EVAL_1488;
  assign _EVAL_2135 = _EVAL_4627 & _EVAL_1824;
  assign _EVAL_2859 = _EVAL_5561 & _EVAL_1155;
  assign _EVAL_5379 = _EVAL_4093 & _EVAL_3418;
  assign _EVAL_4095 = _EVAL_2702 & _EVAL_1653;
  assign _EVAL_1696 = _EVAL_5561 & _EVAL_4992;
  assign _EVAL_5219 = _EVAL_5074 & _EVAL_739;
  assign _EVAL_2558 = _EVAL_6059 & _EVAL_882;
  assign _EVAL_1501 = _EVAL_774 & _EVAL_5543;
  assign _EVAL_1954 = _EVAL_5549 & _EVAL_5299;
  assign _EVAL_2763 = _EVAL_2592 & _EVAL_1488;
  assign _EVAL_2562 = _EVAL_4627 & _EVAL_845;
  assign _EVAL_326 = _EVAL_4755 & _EVAL_4751;
  assign _EVAL_5205 = _EVAL_1145[594];
  assign _EVAL_5149 = _EVAL_2631 & _EVAL_4477;
  assign _EVAL_3174 = _EVAL_4627 & _EVAL_5438;
  assign _EVAL_573 = _EVAL_5074 & _EVAL_4259;
  assign _EVAL_3515 = _EVAL_3945 == 4'h0;
  assign _EVAL_2556 = _EVAL_3414 & _EVAL_6084;
  assign _EVAL_4695 = _EVAL_727 & _EVAL_714;
  assign _EVAL_3622 = _EVAL_2675 & _EVAL_1488;
  assign _EVAL_1692 = _EVAL_1689 & _EVAL_369;
  assign _EVAL_4447 = _EVAL_1675 & _EVAL_2748;
  assign _EVAL_4984 = _EVAL_1082 & _EVAL_5543;
  assign _EVAL_1928 = _EVAL_5478 & _EVAL_847;
  assign _EVAL_5874 = _EVAL_5184 & _EVAL_587;
  assign _EVAL_1068 = _EVAL_5074 & _EVAL_931;
  assign _EVAL_4739 = _EVAL_5816 & _EVAL_4993;
  assign _EVAL_3990 = _EVAL_5662 & _EVAL_3487;
  assign _EVAL_5308 = _EVAL_5068[539];
  assign _EVAL_1329 = _EVAL_905 & _EVAL_3154;
  assign _EVAL_2089 = _EVAL_3632 & _EVAL_3170;
  assign _EVAL_5187 = _EVAL_688 & _EVAL_3154;
  assign _EVAL_3163 = _EVAL_4044 & _EVAL_3418;
  assign _EVAL_3417 = _EVAL_2106 & _EVAL_2748;
  assign _EVAL_5153 = _EVAL_4043 & _EVAL_2892;
  assign _EVAL_1126 = _EVAL_2998 & _EVAL_3487;
  assign _EVAL_4550 = _EVAL_4558 & _EVAL_3379;
  assign _EVAL_1940 = _EVAL_434 & _EVAL_3154;
  assign _EVAL_6065 = _EVAL_5077 & _EVAL_882;
  assign _EVAL_2153 = _EVAL_2753[21];
  assign _EVAL_1463 = _EVAL_4202 & _EVAL_4160;
  assign _EVAL_2775 = _EVAL_4596 & _EVAL_3766;
  assign _EVAL_5215 = _EVAL_5353 & _EVAL_369;
  assign _EVAL_1210 = _EVAL_1361 & _EVAL_3487;
  assign _EVAL_3187 = _EVAL_1393 & _EVAL_369;
  assign _EVAL_319 = _EVAL_921 & _EVAL_882;
  assign _EVAL_5161 = _EVAL_6033 & _EVAL_1009;
  assign _EVAL_4442 = _EVAL_1677 & _EVAL_847;
  assign _EVAL_2700 = _EVAL_774 & _EVAL_2424;
  assign _EVAL_2582 = _EVAL_4627 & _EVAL_374;
  assign _EVAL_2569 = _EVAL_5074 & _EVAL_5936;
  assign _EVAL_5209 = _EVAL_3220 & _EVAL_2424;
  assign _EVAL_537 = _EVAL_4054 & _EVAL_1333;
  assign _EVAL_660 = _EVAL_4235 & _EVAL_2424;
  assign _EVAL_5299 = _EVAL_2236 == 4'hf;
  assign _EVAL_843 = _EVAL_475 & _EVAL_2956;
  assign _EVAL_4372 = _EVAL_974 & _EVAL_3379;
  assign _EVAL_2754 = _EVAL_4856 & _EVAL_6084;
  assign _EVAL_4648 = _EVAL_3082 & _EVAL_5543;
  assign _EVAL_554 = _EVAL_2100 & _EVAL_3418;
  assign _EVAL_826 = _EVAL_5662 & _EVAL_3418;
  assign _EVAL_5285 = _EVAL_1986 & _EVAL_3379;
  assign _EVAL_3897 = _EVAL_3961 & _EVAL_3702;
  assign _EVAL_6005 = _EVAL_4200 & _EVAL_847;
  assign _EVAL_451 = _EVAL_4900 & _EVAL_673;
  assign _EVAL_4560 = _EVAL_1675 & _EVAL_6084;
  assign _EVAL_4171 = _EVAL_594 & _EVAL_1290;
  assign _EVAL_4395 = _EVAL_5023 & _EVAL_3487;
  assign _EVAL_3853 = _EVAL_2972 & _EVAL_1290;
  assign _EVAL_652 = ~_EVAL_4135;
  assign _EVAL_734 = _EVAL_534 & _EVAL_2382;
  assign _EVAL_3510 = _EVAL_4291 & _EVAL_4434;
  assign _EVAL_5477 = _EVAL_5063 & _EVAL_3487;
  assign _EVAL_5134 = _EVAL_3847 & _EVAL_410;
  assign _EVAL_5886 = _EVAL_5493 & _EVAL_5299;
  assign _EVAL_2643 = _EVAL_537 & _EVAL_3313;
  assign _EVAL_940 = _EVAL_4499 & _EVAL_4108;
  assign _EVAL_3068 = _EVAL_3082 & _EVAL_2748;
  assign _EVAL_5129 = _EVAL_3704 & _EVAL_1735;
  assign _EVAL_2255 = _EVAL_5074 & _EVAL_398;
  assign _EVAL_4914 = _EVAL_5132 & _EVAL_3418;
  assign _EVAL_4459 = _EVAL_828 & _EVAL_4108;
  assign _EVAL_5999 = _EVAL_617 & _EVAL_6084;
  assign _EVAL_5631 = _EVAL_4144 & _EVAL_1198;
  assign _EVAL_1542 = _EVAL_2235 & _EVAL_673;
  assign _EVAL_1274 = _EVAL_4627 & _EVAL_2514;
  assign _EVAL_458 = _EVAL_538 & _EVAL_2748;
  assign _EVAL_1852 = _EVAL_4137 & _EVAL_3418;
  assign _EVAL_3723 = _EVAL_4783 & _EVAL_2424;
  assign _EVAL_4224 = _EVAL_5779 & _EVAL_3379;
  assign _EVAL_265 = _EVAL_2454 & _EVAL_5464;
  assign _EVAL_1697 = _EVAL_1446 & _EVAL_2424;
  assign _EVAL_2584 = _EVAL_1945 & _EVAL_1290;
  assign _EVAL_3638 = _EVAL_2842 & _EVAL_1198;
  assign _EVAL_4558 = _EVAL_5074 & _EVAL_5932;
  assign _EVAL_1070 = _EVAL_4563 & _EVAL_6084;
  assign _EVAL_2907 = _EVAL_5144 & _EVAL_3379;
  assign _EVAL_4343 = _EVAL_5609 & _EVAL_2071;
  assign _EVAL_1189 = _EVAL_5741 & _EVAL_997;
  assign _EVAL_5604 = _EVAL_3826 & _EVAL_1198;
  assign _EVAL_3366 = _EVAL_1542 & _EVAL_3398;
  assign _EVAL_6051 = _EVAL_1490 & _EVAL_3379;
  assign _EVAL_2472 = _EVAL_5153 & _EVAL_3508;
  assign _EVAL_5170 = _EVAL_4563 & _EVAL_369;
  assign _EVAL_249 = _EVAL_5561 & _EVAL_2726;
  assign _EVAL_2349 = _EVAL_4596 & _EVAL_1290;
  assign _EVAL_4567 = _EVAL_5430 & _EVAL_673;
  assign _EVAL_4513 = _EVAL_2252 & _EVAL_4477;
  assign _EVAL_4047 = _EVAL_3706 & _EVAL_1488;
  assign _EVAL_3718 = _EVAL_3188 & _EVAL_5289;
  assign _EVAL_2140 = _EVAL_6087 & _EVAL_369;
  assign _EVAL_3418 = _EVAL_4495 != 7'h0;
  assign _EVAL_600 = _EVAL_4627 & _EVAL_3807;
  assign _EVAL_1701 = _EVAL_5561 & _EVAL_202;
  assign _EVAL_1731 = _EVAL_1159[6:5];
  assign _EVAL_865 = _EVAL_3928 & _EVAL_3418;
  assign _EVAL_3103 = _EVAL_4618 & _EVAL_3766;
  assign _EVAL_4428 = _EVAL_1145[537];
  assign _EVAL_5832 = _EVAL_1655 & _EVAL_847;
  assign _EVAL_5439 = _EVAL_4257 & _EVAL_3702;
  assign _EVAL_3659 = _EVAL_3346 & _EVAL_3261;
  assign _EVAL_253 = _EVAL_4044 & _EVAL_847;
  assign _EVAL_5385 = _EVAL_1158 & _EVAL_3487;
  assign _EVAL_3263 = _EVAL_1542 & _EVAL_3154;
  assign _EVAL_2916 = ~_EVAL_560;
  assign _EVAL_4001 = _EVAL_1145[547];
  assign _EVAL_1596 = _EVAL_1145[255];
  assign _EVAL_1012 = _EVAL_1500 & _EVAL_882;
  assign _EVAL_1003 = _EVAL_1920 & _EVAL_3261;
  assign _EVAL_204 = _EVAL_4779 & _EVAL_4891;
  assign _EVAL_873 = _EVAL_5684 & _EVAL_3571;
  assign _EVAL_1658 = _EVAL_5561 & _EVAL_3805;
  assign _EVAL_5525 = _EVAL_4627 & _EVAL_1562;
  assign _EVAL_4762 = _EVAL_2986 & _EVAL_5850;
  assign _EVAL_4502 = _EVAL_5074 & _EVAL_3210;
  assign _EVAL_4018 = _EVAL_5766 & _EVAL_4775;
  assign _EVAL_1058 = _EVAL_5561 & _EVAL_1089;
  assign _EVAL_1599 = _EVAL_362 & _EVAL_1290;
  assign _EVAL_3868 = _EVAL_2550 & _EVAL_4664;
  assign _EVAL_599 = _EVAL_5629 & _EVAL_1277;
  assign _EVAL_3519 = ~_EVAL_1641;
  assign _EVAL_2628 = _EVAL_594 & _EVAL_3766;
  assign _EVAL_807 = _EVAL_4904 & _EVAL_673;
  assign _EVAL_1557 = _EVAL_5074 & _EVAL_374;
  assign _EVAL_2465 = _EVAL_1145[591];
  assign _EVAL_1452 = _EVAL_5598 & _EVAL_847;
  assign _EVAL_656 = _EVAL_5132 & _EVAL_882;
  assign _EVAL_4192 = _EVAL_1977 & _EVAL_3379;
  assign _EVAL_4784 = _EVAL_5427 & _EVAL_3398;
  assign _EVAL_2870 = _EVAL_5795 & _EVAL_4664;
  assign _EVAL_5159 = _EVAL_1536 & _EVAL_369;
  assign _EVAL_1559 = _EVAL_4888 & _EVAL_3702;
  assign _EVAL_5672 = _EVAL_4596 & _EVAL_5753;
  assign _EVAL_4723 = _EVAL_3815 & _EVAL_5850;
  assign _EVAL_1034 = _EVAL_3066 & _EVAL_3379;
  assign _EVAL_1695 = _EVAL_5068[516];
  assign _EVAL_4433 = _EVAL_4627 & _EVAL_1175;
  assign _EVAL_1511 = _EVAL_1971 & _EVAL_2969;
  assign _EVAL_4872 = ~_EVAL_4808;
  assign _EVAL_4305 = _EVAL_6051 & _EVAL_4751;
  assign _EVAL_5583 = _EVAL_2454 & _EVAL_2382;
  assign _EVAL_1679 = _EVAL_3993 & _EVAL_847;
  assign _EVAL_523 = _EVAL_1316[7:0];
  assign _EVAL_5056 = _EVAL_5869 & _EVAL_3487;
  assign _EVAL_323 = _EVAL_1316[19:16];
  assign _EVAL_5037 = _EVAL_2192 & _EVAL_3702;
  assign _EVAL_4724 = _EVAL_284 & _EVAL_1488;
  assign _EVAL_2913 = _EVAL_5561 & _EVAL_5217;
  assign _EVAL_4892 = _EVAL_5869 & _EVAL_847;
  assign _EVAL_974 = _EVAL_5074 & _EVAL_4225;
  assign _EVAL_2831 = _EVAL_1446 & _EVAL_5543;
  assign _EVAL_726 = ~_EVAL_1187;
  assign _EVAL_3577 = _EVAL_2646 & _EVAL_1924;
  assign _EVAL_3281 = _EVAL_4627 & _EVAL_5593;
  assign _EVAL_5105 = _EVAL_1677 & _EVAL_3154;
  assign _EVAL_1733 = _EVAL_1854 & _EVAL_3398;
  assign _EVAL_1419 = _EVAL_3402 & _EVAL_3379;
  assign _EVAL_5408 = _EVAL_6075 & _EVAL_3398;
  assign _EVAL_5319 = _EVAL_1242 & _EVAL_3154;
  assign _EVAL_882 = _EVAL_408 != 7'h0;
  assign _EVAL_3130 = _EVAL_2545 & _EVAL_3379;
  assign _EVAL_2713 = _EVAL_5162 & _EVAL_369;
  assign _EVAL_239 = _EVAL_3787 & _EVAL_1009;
  assign _EVAL_4755 = _EVAL_4565 & _EVAL_3379;
  assign _EVAL_1647 = _EVAL_5153 & _EVAL_4993;
  assign _EVAL_4993 = _EVAL_334 != 8'h0;
  assign _EVAL_4359 = _EVAL_4235 & _EVAL_2748;
  assign _EVAL_878 = _EVAL_6087 & _EVAL_1488;
  assign _EVAL_2250 = _EVAL_5193 & _EVAL_1488;
  assign _EVAL_1582 = _EVAL_1145[517];
  assign _EVAL_6032 = _EVAL_2963 & _EVAL_3379;
  assign _EVAL_461 = _EVAL_528 & _EVAL_3170;
  assign _EVAL_3265 = _EVAL_4338 & _EVAL_926;
  assign _EVAL_1434 = _EVAL_1344 & _EVAL_3154;
  assign _EVAL_3199 = _EVAL_5353 & _EVAL_2748;
  assign _EVAL_2049 = _EVAL_4745 & _EVAL_3418;
  assign _EVAL_4075 = _EVAL_3183 & _EVAL_2748;
  assign _EVAL_1773 = _EVAL_3524 & _EVAL_3702;
  assign _EVAL_5692 = _EVAL_3364 & _EVAL_882;
  assign _EVAL_1754 = _EVAL_4106 & _EVAL_4664;
  assign _EVAL_1373 = _EVAL_1312 & _EVAL_6084;
  assign _EVAL_2427 = _EVAL_1312 & _EVAL_2969;
  assign _EVAL_4607 = _EVAL_6087 & _EVAL_5543;
  assign _EVAL_5774 = _EVAL_3032 & _EVAL_587;
  assign _EVAL_243 = _EVAL_4745 & _EVAL_3398;
  assign _EVAL_1310 = _EVAL_4588 & _EVAL_539;
  assign _EVAL_1300 = _EVAL_5068[522];
  assign _EVAL_1319 = _EVAL_4870 & _EVAL_3284;
  assign _EVAL_5896 = _EVAL_2585 & _EVAL_3487;
  assign _EVAL_2294 = _EVAL_6022 & _EVAL_2424;
  assign _EVAL_1266 = _EVAL_1039 & _EVAL_3418;
  assign _EVAL_4324 = _EVAL_2005 & _EVAL_6084;
  assign _EVAL_709 = _EVAL_1316[23:17];
  assign _EVAL_4393 = _EVAL_5561 & _EVAL_5266;
  assign _EVAL_2275 = _EVAL_3710 & _EVAL_369;
  assign _EVAL_1584 = ~_EVAL_2360;
  assign _EVAL_2872 = _EVAL_5869 & _EVAL_3154;
  assign _EVAL_2338 = _EVAL_2038 & _EVAL_3379;
  assign _EVAL_2445 = _EVAL_528 & _EVAL_5850;
  assign _EVAL_989 = _EVAL_402 & _EVAL_3284;
  assign _EVAL_1312 = _EVAL_2232 & _EVAL_3379;
  assign _EVAL_4209 = ~_EVAL_2357;
  assign _EVAL_3849 = _EVAL_3436 & _EVAL_3313;
  assign _EVAL_4254 = _EVAL_1392 & _EVAL_673;
  assign _EVAL_2759 = _EVAL_2100 & _EVAL_882;
  assign _EVAL_509 = _EVAL_4755 & _EVAL_5850;
  assign _EVAL_3243 = _EVAL_5542 & _EVAL_4751;
  assign _EVAL_528 = _EVAL_4750 & _EVAL_3379;
  assign _EVAL_4915 = _EVAL_1920 & _EVAL_4477;
  assign _EVAL_4471 = _EVAL_3689 & _EVAL_6084;
  assign _EVAL_1677 = _EVAL_1151 & _EVAL_673;
  assign _EVAL_216 = _EVAL_1393 & _EVAL_3702;
  assign _EVAL_1254 = _EVAL_5561 & _EVAL_3757;
  assign _EVAL_4287 = ~_EVAL_3294;
  assign _EVAL_5601 = _EVAL_3220 & _EVAL_1488;
  assign _EVAL_1067 = _EVAL_941 & _EVAL_673;
  assign _EVAL_4544 = _EVAL_4604 & _EVAL_4664;
  assign _EVAL_486 = _EVAL_222 & _EVAL_3379;
  assign _EVAL_588 = _EVAL_2233 & _EVAL_5573;
  assign _EVAL_1203 = _EVAL_1962 & _EVAL_3284;
  assign _EVAL_5530 = _EVAL_5074 & _EVAL_3329;
  assign _EVAL_2926 = _EVAL_688 & _EVAL_882;
  assign _EVAL_581 = _EVAL_2564 & _EVAL_3379;
  assign _EVAL_1523 = _EVAL_5561 & _EVAL_5984;
  assign _EVAL_586 = _EVAL_623 & _EVAL_3702;
  assign _EVAL_3331 = _EVAL_1158 & _EVAL_3398;
  assign _EVAL_2213 = _EVAL_1675 & _EVAL_5543;
  assign _EVAL_3147 = _EVAL_4567 & _EVAL_4477;
  assign _EVAL_2602 = _EVAL_1361 & _EVAL_3154;
  assign _EVAL_1539 = _EVAL_4661 & _EVAL_4775;
  assign _EVAL_1781 = _EVAL_1536 & _EVAL_6084;
  assign _EVAL_3993 = _EVAL_3006 & _EVAL_673;
  assign _EVAL_4126 = _EVAL_1731 == 2'h3;
  assign _EVAL_2966 = _EVAL_5478 & _EVAL_882;
  assign _EVAL_770 = _EVAL_6087 & _EVAL_6084;
  assign _EVAL_1711 = _EVAL_2550 & _EVAL_5289;
  assign _EVAL_3600 = _EVAL_3346 & _EVAL_3418;
  assign _EVAL_3262 = _EVAL_446 & _EVAL_2956;
  assign _EVAL_5071 = _EVAL_932 & _EVAL_1198;
  assign _EVAL_2607 = _EVAL_1343 & _EVAL_3379;
  assign _EVAL_4261 = _EVAL_1034 & _EVAL_3284;
  assign _EVAL_5121 = _EVAL_617 & _EVAL_2969;
  assign _EVAL_2942 = _EVAL_5023 & _EVAL_847;
  assign _EVAL_5490 = _EVAL_5549 & _EVAL_3284;
  assign _EVAL_5199 = _EVAL_479 & _EVAL_2969;
  assign _EVAL_4768 = _EVAL_3032 & _EVAL_5289;
  assign _EVAL_2345 = _EVAL_935 & _EVAL_369;
  assign _EVAL_2919 = _EVAL_5246 & _EVAL_3261;
  assign _EVAL_2609 = _EVAL_1145[646];
  assign _EVAL_5354 = _EVAL_4836 & _EVAL_3412;
  assign _EVAL_3867 = _EVAL_4627 & _EVAL_464;
  assign _EVAL_917 = _EVAL_4224 & _EVAL_5464;
  assign _EVAL_3055 = _EVAL_1316[4:1];
  assign _EVAL_5514 = _EVAL_5162 & _EVAL_1488;
  assign _EVAL_5680 = _EVAL_3787 & _EVAL_587;
  assign _EVAL_4561 = _EVAL_2585 & _EVAL_3398;
  assign _EVAL_510 = _EVAL_606 & _EVAL_4126;
  assign _EVAL_3007 = _EVAL_4257 & _EVAL_5543;
  assign _EVAL_1125 = _EVAL_390 & _EVAL_673;
  assign _EVAL_3364 = _EVAL_3804 & _EVAL_673;
  assign _EVAL_373 = _EVAL_407 & _EVAL_2748;
  assign _EVAL_775 = _EVAL_3581 & _EVAL_5445;
  assign _EVAL_5128 = _EVAL_6087 & _EVAL_3702;
  assign _EVAL_2379 = _EVAL_6080 & _EVAL_4109;
  assign _EVAL_3777 = _EVAL_5450 & _EVAL_4108;
  assign _EVAL_4316 = _EVAL_5478 & _EVAL_3418;
  assign _EVAL_2210 = _EVAL_4627 & _EVAL_885;
  assign _EVAL_4453 = _EVAL_2471 & _EVAL_3418;
  assign _EVAL_2253 = _EVAL_4488 & _EVAL_3487;
  assign _EVAL_5724 = _EVAL_5561 & _EVAL_4386;
  assign _EVAL_2423 = _EVAL_5561 & _EVAL_1528;
  assign _EVAL_3218 = _EVAL_1145[540];
  assign _EVAL_5512 = _EVAL_2631 & _EVAL_3154;
  assign _EVAL_157 = _EVAL_2005 & _EVAL_1488;
  assign _EVAL_5493 = _EVAL_1068 & _EVAL_3379;
  assign _EVAL_1878 = _EVAL_4627 & _EVAL_2425;
  assign _EVAL_3371 = _EVAL_735 & _EVAL_2382;
  assign _EVAL_3445 = _EVAL_5074 & _EVAL_4341;
  assign _EVAL_3988 = _EVAL_5344 & _EVAL_3170;
  assign _EVAL_5723 = _EVAL_5249 & _EVAL_2783;
  assign _EVAL_1921 = _EVAL_1945 & _EVAL_587;
  assign _EVAL_4499 = _EVAL_3113 & _EVAL_3379;
  assign _EVAL_2529 = _EVAL_2902 & _EVAL_3702;
  assign _EVAL_1450 = _EVAL_2454 & _EVAL_4109;
  assign _EVAL_4838 = _EVAL_4254 & _EVAL_4664;
  assign _EVAL_3974 = _EVAL_3787 & _EVAL_4664;
  assign _EVAL_4413 = _EVAL_5162 & _EVAL_2424;
  assign _EVAL_5936 = _EVAL_1145[666];
  assign _EVAL_159 = _EVAL_594 & _EVAL_4775;
  assign _EVAL_5042 = _EVAL_5028 & _EVAL_5464;
  assign _EVAL_5292 = _EVAL_538 & _EVAL_2969;
  assign _EVAL_1580 = _EVAL_451 & _EVAL_4788;
  assign _EVAL_5238 = _EVAL_5930 & _EVAL_369;
  assign _EVAL_3350 = _EVAL_1159[31:1];
  assign _EVAL_4429 = _EVAL_1361 & _EVAL_3261;
  assign _EVAL_4320 = _EVAL_3815 & _EVAL_4108;
  assign _EVAL_971 = _EVAL_4627 & _EVAL_3218;
  assign _EVAL_2223 = _EVAL_2454 & _EVAL_1735;
  assign _EVAL_2171 = _EVAL_3706 & _EVAL_3702;
  assign _EVAL_2908 = _EVAL_3651 & _EVAL_369;
  assign _EVAL_3702 = _EVAL_1316[24];
  assign _EVAL_2742 = _EVAL_3961 & _EVAL_1488;
  assign _EVAL_5998 = _EVAL_3077 & _EVAL_3379;
  assign _EVAL_3388 = _EVAL_383 != 2'h0;
  assign _EVAL_1894 = _EVAL_589 & _EVAL_5464;
  assign _EVAL_3569 = _EVAL_4707 & _EVAL_1009;
  assign _EVAL_2194 = _EVAL_6022 & _EVAL_6084;
  assign _EVAL_4644 = _EVAL_4563 & _EVAL_3702;
  assign _EVAL_3792 = _EVAL_5344 & _EVAL_4108;
  assign _EVAL_1505 = _EVAL_1393 & _EVAL_1488;
  assign _EVAL_4134 = _EVAL_5561 & _EVAL_4651;
  assign _EVAL_1491 = _EVAL_5561 & _EVAL_2884;
  assign _EVAL_2354 = _EVAL_2338 & _EVAL_5543;
  assign _EVAL_3034 = _EVAL_783 & _EVAL_4522;
  assign _EVAL_4424 = _EVAL_4627 & _EVAL_5760;
  assign _EVAL_2390 = _EVAL_4627 & _EVAL_3761;
  assign _EVAL_4604 = _EVAL_3740 & _EVAL_673;
  assign _EVAL_5175 = _EVAL_4841 & _EVAL_3154;
  assign _EVAL_4593 = _EVAL_3451 & _EVAL_3487;
  assign _EVAL_3952 = _EVAL_4550 & _EVAL_369;
  assign _EVAL_5639 = _EVAL_5598 & _EVAL_3154;
  assign _EVAL_3124 = _EVAL_1971 & _EVAL_2748;
  assign _EVAL_1088 = _EVAL_5676 & _EVAL_847;
  assign _EVAL_4961 = ~_EVAL_1671;
  assign _EVAL_3137 = _EVAL_2877 & _EVAL_3702;
  assign _EVAL_2592 = _EVAL_5380 & _EVAL_3379;
  assign _EVAL_5162 = _EVAL_1841 & _EVAL_3379;
  assign _EVAL_4870 = _EVAL_3825 & _EVAL_3379;
  assign _EVAL_4946 = _EVAL_2646 & _EVAL_5281;
  assign _EVAL_4190 = _EVAL_4627 & _EVAL_4154;
  assign _EVAL_4537 = _EVAL_528 & _EVAL_4751;
  assign _EVAL_5947 = _EVAL_3082 & _EVAL_3702;
  assign _EVAL_5654 = _EVAL_2868 & _EVAL_4477;
  assign _EVAL_1370 = _EVAL_183 & _EVAL_673;
  assign _EVAL_209 = _EVAL_2877 & _EVAL_2748;
  assign _EVAL_2067 = _EVAL_5344 & _EVAL_5850;
  assign _EVAL_2640 = _EVAL_1971 & _EVAL_5543;
  assign _EVAL_5072 = _EVAL_479 & _EVAL_6084;
  assign _EVAL_4335 = _EVAL_4577 & _EVAL_1009;
  assign _EVAL_973 = _EVAL_4692 & _EVAL_3261;
  assign _EVAL_4952 = _EVAL_3632 & _EVAL_4109;
  assign _EVAL_4617 = _EVAL_6032 & _EVAL_1488;
  assign _EVAL_3424 = _EVAL_5766 & _EVAL_5289;
  assign _EVAL_2597 = _EVAL_5561 & _EVAL_1706;
  assign _EVAL_536 = _EVAL_1536 & _EVAL_2748;
  assign _EVAL_4847 = _EVAL_1962 & _EVAL_5299;
  assign _EVAL_4551 = _EVAL_1316[23:16];
  assign _EVAL_5809 = _EVAL_251 & _EVAL_2748;
  assign _EVAL_1256 = _EVAL_5074 & _EVAL_5937;
  assign _EVAL_4907 = _EVAL_2242 & _EVAL_5543;
  assign _EVAL_3459 = _EVAL_1945 & _EVAL_1009;
  assign _EVAL_1622 = _EVAL_5084 & _EVAL_673;
  assign _EVAL_1960 = _EVAL_5274 & _EVAL_673;
  assign _EVAL_818 = _EVAL_4627 & _EVAL_4225;
  assign _EVAL_1285 = _EVAL_2793 & _EVAL_3154;
  assign _EVAL_3247 = _EVAL_1622 & _EVAL_1290;
  assign _EVAL_5193 = _EVAL_818 & _EVAL_3379;
  assign _EVAL_2877 = _EVAL_2288 & _EVAL_3379;
  assign _EVAL_5756 = _EVAL_4604 & _EVAL_4775;
  assign _EVAL_5063 = _EVAL_1627 & _EVAL_673;
  assign _EVAL_2604 = _EVAL_5788 & _EVAL_4108;
  assign _EVAL_346 = _EVAL_4367 & _EVAL_2615;
  assign _EVAL_5613 = _EVAL_5766 & _EVAL_4664;
  assign _EVAL_1144 = _EVAL_5068[537];
  assign _EVAL_5043 = _EVAL_4627 & _EVAL_1582;
  assign _EVAL_1014 = _EVAL_298 & _EVAL_2320;
  assign _EVAL_3373 = ~_EVAL_3580;
  assign _EVAL_1895 = _EVAL_5788 & _EVAL_1735;
  assign _EVAL_2676 = _EVAL_4627 & _EVAL_3461;
  assign _EVAL_2314 = _EVAL_2205 & _EVAL_4109;
  assign _EVAL_2214 = _EVAL_4080 & _EVAL_3184;
  assign _EVAL_413 = _EVAL_1145[592];
  assign _EVAL_3664 = _EVAL_3070 & _EVAL_2956;
  assign _EVAL_817 = _EVAL_5077 & _EVAL_3487;
  assign _EVAL_2440 = _EVAL_4689 & _EVAL_2382;
  assign _EVAL_3362 = _EVAL_3346 & _EVAL_3398;
  assign _EVAL_2373 = _EVAL_1677 & _EVAL_3487;
  assign _EVAL_2131 = _EVAL_5561 & _EVAL_1762;
  assign _EVAL_4793 = _EVAL_5561 & _EVAL_2864;
  assign _EVAL_4066 = _EVAL_4757 & _EVAL_847;
  assign _EVAL_434 = _EVAL_5006 & _EVAL_673;
  assign _EVAL_668 = _EVAL_971 & _EVAL_3379;
  assign _EVAL_5005 = _EVAL_3350 != 31'h0;
  assign _EVAL_5970 = _EVAL_4627 & _EVAL_177;
  assign _EVAL_3097 = _EVAL_1125 & _EVAL_4477;
  assign _EVAL_3182 = _EVAL_965 & _EVAL_4788;
  assign _EVAL_3601 = _EVAL_3706 & _EVAL_369;
  assign _EVAL_3000 = _EVAL_3704 & _EVAL_4109;
  assign _EVAL_4059 = _EVAL_2646 & _EVAL_1653;
  assign _EVAL_1955 = _EVAL_3107 & _EVAL_2748;
  assign _EVAL_2803 = _EVAL_2675 & _EVAL_5543;
  assign _EVAL_3557 = _EVAL_1876 & _EVAL_882;
  assign _EVAL_4525 = _EVAL_4084 & _EVAL_3379;
  assign _EVAL_4062 = _EVAL_2205 & _EVAL_3170;
  assign _EVAL_3840 = _EVAL_2873 & _EVAL_1198;
  assign _EVAL_4464 = _EVAL_620 & _EVAL_4108;
  assign _EVAL_722 = ~_EVAL_3946;
  assign _EVAL_4516 = _EVAL_4841 & _EVAL_3418;
  assign _EVAL_2507 = _EVAL_1145[513];
  assign _EVAL_3073 = _EVAL_4974 & _EVAL_5850;
  assign _EVAL_3821 = ~_EVAL_2837;
  assign _EVAL_2785 = _EVAL_4372 & _EVAL_5543;
  assign _EVAL_2062 = _EVAL_1533 & _EVAL_4109;
  assign _EVAL_4473 = _EVAL_880 & _EVAL_193;
  assign _EVAL_773 = _EVAL_1655 & _EVAL_3418;
  assign _EVAL_251 = _EVAL_4947 & _EVAL_3379;
  assign _EVAL_3539 = _EVAL_905 & _EVAL_882;
  assign _EVAL_3242 = _EVAL_5074 & _EVAL_2425;
  assign _EVAL_3919 = _EVAL_4856 & _EVAL_2748;
  assign _EVAL_1750 = _EVAL_5206 & _EVAL_5299;
  assign _EVAL_2986 = _EVAL_5446 & _EVAL_3379;
  assign TLMonitor__EVAL_5 = _EVAL_131;
  assign _EVAL_5950 = _EVAL_2096 & _EVAL_364;
  assign _EVAL_2576 = _EVAL_3710 & _EVAL_2748;
  assign _EVAL_5508 = _EVAL_4014 & _EVAL_746;
  assign _EVAL_4722 = _EVAL_6022 & _EVAL_1488;
  assign _EVAL_3678 = _EVAL_1067 & _EVAL_5753;
  assign _EVAL_2663 = _EVAL_4604 & _EVAL_587;
  assign _EVAL_2531 = _EVAL_407 & _EVAL_2424;
  assign _EVAL_3061 = _EVAL_3346 & _EVAL_847;
  assign _EVAL_5383 = _EVAL_4325 & _EVAL_3379;
  assign _EVAL_897 = _EVAL_5992 & _EVAL_3379;
  assign _EVAL_1412 = _EVAL_3993 & _EVAL_3487;
  assign _EVAL_4782 = _EVAL_4627 & _EVAL_5656;
  assign _EVAL_3650 = _EVAL_4627 & _EVAL_3701;
  assign _EVAL_290 = _EVAL_2241 & _EVAL_1488;
  assign _EVAL_1909 = _EVAL_3704 & _EVAL_4108;
  assign _EVAL_2606 = _EVAL_5054 & _EVAL_3418;
  assign _EVAL_5904 = _EVAL_5561 & _EVAL_2898;
  assign _EVAL_5218 = _EVAL_2205 & _EVAL_5464;
  assign _EVAL_4656 = _EVAL_1145[581];
  assign _EVAL_2792 = _EVAL_5549 & _EVAL_2956;
  assign _EVAL_2313 = _EVAL_1136 & _EVAL_3261;
  assign _EVAL_735 = _EVAL_1878 & _EVAL_3379;
  assign _EVAL_512 = _EVAL_3421 & _EVAL_4477;
  assign _EVAL_769 = _EVAL_4697 & _EVAL_673;
  assign _EVAL_2644 = _EVAL_6033 & _EVAL_4664;
  assign _EVAL_4519 = _EVAL_4916 & _EVAL_4108;
  assign _EVAL_932 = _EVAL_6024 & _EVAL_3379;
  assign _EVAL_2678 = _EVAL_4909 & _EVAL_4993;
  assign _EVAL_5705 = _EVAL_4455 & _EVAL_3379;
  assign _EVAL_3889 = _EVAL_5561 & _EVAL_3613;
  assign _EVAL_258 = _EVAL_1745 & _EVAL_4108;
  assign _EVAL_2631 = _EVAL_5313 & _EVAL_673;
  assign _EVAL_2551 = _EVAL_1202 & _EVAL_882;
  assign _EVAL_4675 = _EVAL_1664 & _EVAL_321;
  assign _EVAL_3829 = _EVAL_1542 & _EVAL_4477;
  assign _EVAL_4054 = _EVAL_5561 & _EVAL_5800;
  assign _EVAL_2318 = _EVAL_3704 & _EVAL_5850;
  assign _EVAL_5252 = _EVAL_5561 & _EVAL_1087;
  assign _EVAL_2076 = _EVAL_5561 & _EVAL_550;
  assign _EVAL_4874 = _EVAL_2005 & _EVAL_2424;
  assign _EVAL_2687 = _EVAL_1622 & _EVAL_587;
  assign _EVAL_5189 = _EVAL_5676 & _EVAL_3261;
  assign _EVAL_3451 = _EVAL_2913 & _EVAL_673;
  assign _EVAL_2513 = _EVAL_4888 & _EVAL_369;
  assign _EVAL_767 = _EVAL_4419 & _EVAL_882;
  assign _EVAL_635 = _EVAL_4627 & _EVAL_2601;
  assign _EVAL_2677 = _EVAL_3935 & _EVAL_5543;
  assign _EVAL_5964 = _EVAL_932 & _EVAL_5299;
  assign _EVAL_5298 = _EVAL_5246 & _EVAL_847;
  assign _EVAL_2103 = _EVAL_6033 & _EVAL_4775;
  assign _EVAL_5160 = _EVAL_3451 & _EVAL_4477;
  assign _EVAL_2347 = _EVAL_2037 & _EVAL_5543;
  assign _EVAL_3296 = _EVAL_2972 & _EVAL_5753;
  assign _EVAL_4364 = _EVAL_905 & _EVAL_3418;
  assign _EVAL_5235 = _EVAL_6033 & _EVAL_1290;
  assign _EVAL_1053 = _EVAL_3032 & _EVAL_4664;
  assign _EVAL_395 = _EVAL_1145[601];
  assign _EVAL_5700 = _EVAL_5074 & _EVAL_395;
  assign _EVAL_6083 = _EVAL_3421 & _EVAL_847;
  assign _EVAL_2619 = _EVAL_4149 & _EVAL_1488;
  assign _EVAL_4756 = _EVAL_4106 & _EVAL_5753;
  assign _EVAL_3596 = _EVAL_5561 & _EVAL_2632;
  assign _EVAL_330 = _EVAL_3961 & _EVAL_369;
  assign _EVAL_2151 = _EVAL_5074 & _EVAL_2480;
  assign _EVAL_5868 = _EVAL_3216 & _EVAL_3154;
  assign _EVAL_2974 = _EVAL_4974 & _EVAL_5464;
  assign _EVAL_4729 = _EVAL_2471 & _EVAL_882;
  assign _EVAL_1328 = _EVAL_1364 & _EVAL_3284;
  assign _EVAL_4930 = _EVAL_3935 & _EVAL_3702;
  assign _EVAL_3153 = _EVAL_668 & _EVAL_2424;
  assign _EVAL_746 = ~_EVAL_4932;
  assign _EVAL_4743 = _EVAL_3961 & _EVAL_5543;
  assign _EVAL_3118 = _EVAL_4175 & _EVAL_3261;
  assign _EVAL_1640 = _EVAL_2471 & _EVAL_3261;
  assign _EVAL_5327 = _EVAL_4955 & _EVAL_2999;
  assign _EVAL_4375 = _EVAL_5068[532];
  assign _EVAL_1194 = _EVAL_4627 & _EVAL_395;
  assign _EVAL_1932 = _EVAL_1145[606];
  assign _EVAL_252 = _EVAL_1689 & _EVAL_5543;
  assign _EVAL_1612 = _EVAL_2998 & _EVAL_3261;
  assign _EVAL_4667 = _EVAL_4627 & _EVAL_227;
  assign TLMonitor__EVAL_12 = {{2'd0}, _EVAL_4791};
  assign _EVAL_1655 = _EVAL_2145 & _EVAL_673;
  assign _EVAL_387 = _EVAL_4856 & _EVAL_5543;
  assign _EVAL_2219 = _EVAL_4581 & _EVAL_3284;
  assign _EVAL_1104 = _EVAL_3226 & _EVAL_4751;
  assign _EVAL_4113 = _EVAL_1633 & _EVAL_6084;
  assign _EVAL_474 = _EVAL_778 & _EVAL_5289;
  assign _EVAL_4100 = ~_EVAL_5484;
  assign _EVAL_5826 = _EVAL_5561 & _EVAL_676;
  assign _EVAL_1546 = _EVAL_1393 & _EVAL_2424;
  assign _EVAL_3773 = _EVAL_1553 & _EVAL_587;
  assign _EVAL_3079 = _EVAL_2986 & _EVAL_4108;
  assign _EVAL_2729 = _EVAL_4254 & _EVAL_5753;
  assign _EVAL_2386 = _EVAL_5132 & _EVAL_4477;
  assign _EVAL_5776 = ~_EVAL_1820;
  assign _EVAL_4751 = _EVAL_2236 != 4'h0;
  assign _EVAL_3901 = _EVAL_3844 & _EVAL_369;
  assign _EVAL_5296 = _EVAL_5342 & _EVAL_3284;
  assign _EVAL_5992 = _EVAL_5074 & _EVAL_1069;
  assign _EVAL_3556 = _EVAL_5023 & _EVAL_3154;
  assign _EVAL_1317 = _EVAL_1121 & _EVAL_5977;
  assign _EVAL_3260 = _EVAL_5542 & _EVAL_4109;
  assign _EVAL_2839 = _EVAL_828 & _EVAL_4751;
  assign _EVAL_4867 = _EVAL_4627 & _EVAL_925;
  assign _EVAL_4531 = _EVAL_5344 & _EVAL_5464;
  assign _EVAL_2368 = _EVAL_807 & _EVAL_3766;
  assign _EVAL_1778 = _EVAL_2907 & _EVAL_1488;
  assign _EVAL_2256 = _EVAL_3301 & _EVAL_5299;
  assign _EVAL_4783 = _EVAL_335 & _EVAL_3379;
  assign _EVAL_4713 = _EVAL_5561 & _EVAL_4293;
  assign _EVAL_1099 = _EVAL_5561 & _EVAL_5556;
  assign _EVAL_4322 = _EVAL_2538 & _EVAL_3379;
  assign _EVAL_3026 = _EVAL_6059 & _EVAL_4477;
  assign _EVAL_4311 = _EVAL_3347 & _EVAL_673;
  assign _EVAL_1835 = _EVAL_4604 & _EVAL_5753;
  assign _EVAL_4757 = _EVAL_449 & _EVAL_673;
  assign _EVAL_3028 = _EVAL_3451 & _EVAL_847;
  assign _EVAL_4166 = _EVAL_1854 & _EVAL_4477;
  assign _EVAL_4407 = ~_EVAL_6030;
  assign _EVAL_453 = _EVAL_362 & _EVAL_5289;
  assign _EVAL_2438 = ~_EVAL_3607;
  assign _EVAL_5422 = _EVAL_4581 & _EVAL_1198;
  assign _EVAL_3060 = _EVAL_5074 & _EVAL_5739;
  assign _EVAL_1007 = _EVAL_5398 & _EVAL_1488;
  assign _EVAL_4351 = _EVAL_4024 & _EVAL_3379;
  assign _EVAL_2795 = _EVAL_3188 & _EVAL_3766;
  assign _EVAL_1479 = _EVAL_4202 & _EVAL_3313;
  assign _EVAL_4017 = _EVAL_3961 & _EVAL_6084;
  assign _EVAL_2509 = _EVAL_3188 & _EVAL_1009;
  assign _EVAL_5273 = _EVAL_1854 & _EVAL_847;
  assign _EVAL_4231 = _EVAL_551 & _EVAL_5299;
  assign _EVAL_2685 = _EVAL_4219 & _EVAL_1488;
  assign _EVAL_4925 = _EVAL_668 & _EVAL_3702;
  assign _EVAL_5283 = _EVAL_3710 & _EVAL_5543;
  assign _EVAL_5367 = _EVAL_3981 & _EVAL_4477;
  assign _EVAL_521 = _EVAL_5528 & _EVAL_1009;
  assign _EVAL_3953 = _EVAL_5068[542];
  assign _EVAL_2808 = _EVAL_1034 & _EVAL_2956;
  assign _EVAL_1906 = _EVAL_5028 & _EVAL_4751;
  assign _EVAL_1853 = _EVAL_4224 & _EVAL_3170;
  assign _EVAL_1703 = _EVAL_2251 & _EVAL_3702;
  assign _EVAL_2172 = _EVAL_5074 & _EVAL_530;
  assign _EVAL_2087 = _EVAL_302 & _EVAL_2748;
  assign _EVAL_821 = _EVAL_857 & _EVAL_6084;
  assign _EVAL_3759 = _EVAL_2753[4];
  assign _EVAL_3503 = _EVAL_4707 & _EVAL_4664;
  assign _EVAL_2221 = _EVAL_1312 & _EVAL_2748;
  assign _EVAL_2620 = _EVAL_383 == 2'h3;
  assign _EVAL_3333 = _EVAL_617 & _EVAL_5543;
  assign _EVAL_4317 = _EVAL_3706 & _EVAL_2748;
  assign _EVAL_1151 = _EVAL_5561 & _EVAL_1173;
  assign _EVAL_538 = _EVAL_2562 & _EVAL_3379;
  assign _EVAL_754 = _EVAL_3981 & _EVAL_3154;
  assign _EVAL_3935 = _EVAL_3323 & _EVAL_3379;
  assign _EVAL_310 = _EVAL_4596 & _EVAL_1009;
  assign _EVAL_5305 = _EVAL_5784 & _EVAL_3379;
  assign _EVAL_3909 = _EVAL_5561 & _EVAL_543;
  assign _EVAL_3315 = _EVAL_2753[2];
  assign _EVAL_2084 = _EVAL_2675 & _EVAL_369;
  assign _EVAL_5531 = _EVAL_4623 & _EVAL_5543;
  assign _EVAL_4031 = _EVAL_5450 & _EVAL_5464;
  assign _EVAL_679 = _EVAL_3712 & _EVAL_3379;
  assign TLMonitor__EVAL_6 = _EVAL_26;
  assign _EVAL_4102 = _EVAL_3082 & _EVAL_2969;
  assign _EVAL_836 = _EVAL_2005 & _EVAL_2748;
  assign _EVAL_4327 = _EVAL_3202 & _EVAL_1488;
  assign _EVAL_3917 = _EVAL_4755 & _EVAL_4109;
  assign _EVAL_3860 = _EVAL_3581 & _EVAL_1924;
  assign _EVAL_1652 = _EVAL_5705 & _EVAL_2748;
  assign _EVAL_2594 = _EVAL_1125 & _EVAL_3154;
  assign _EVAL_5816 = _EVAL_4867 & _EVAL_3379;
  assign _EVAL_3348 = _EVAL_4707 & _EVAL_4775;
  assign _EVAL_2715 = _EVAL_1622 & _EVAL_4664;
  assign _EVAL_694 = _EVAL_5662 & _EVAL_3261;
  assign _EVAL_1945 = _EVAL_5826 & _EVAL_673;
  assign _EVAL_3491 = _EVAL_3414 & _EVAL_5543;
  assign _EVAL_535 = _EVAL_4175 & _EVAL_3398;
  assign _EVAL_1512 = _EVAL_3451 & _EVAL_3154;
  assign _EVAL_4011 = _EVAL_5427 & _EVAL_4477;
  assign _EVAL_5953 = _EVAL_3624 & _EVAL_3702;
  assign _EVAL_1387 = _EVAL_1718 & _EVAL_5569;
  assign _EVAL_1008 = _EVAL_5561 & _EVAL_4246;
  assign _EVAL_3303 = _EVAL_5766 & _EVAL_1290;
  assign _EVAL_6047 = _EVAL_2907 & _EVAL_5543;
  assign _EVAL_623 = _EVAL_4433 & _EVAL_3379;
  assign _EVAL_1757 = _EVAL_5930 & _EVAL_2424;
  assign _EVAL_5858 = _EVAL_4525 & _EVAL_5850;
  assign _EVAL_2947 = _EVAL_668 & _EVAL_5543;
  assign _EVAL_1344 = _EVAL_3232 & _EVAL_673;
  assign _EVAL_3468 = _EVAL_5705 & _EVAL_2424;
  assign _EVAL_5775 = _EVAL_4623 & _EVAL_2748;
  assign _EVAL_357 = _EVAL_2229 & _EVAL_1808;
  assign _EVAL_196 = _EVAL_3322 & _EVAL_5299;
  assign _EVAL_1838 = _EVAL_751 & _EVAL_3702;
  assign _EVAL_4263 = _EVAL_5561 & _EVAL_1665;
  assign _EVAL_4597 = _EVAL_5074 & _EVAL_4703;
  assign _EVAL_3543 = _EVAL_4623 & _EVAL_3702;
  assign _EVAL_2093 = _EVAL_1145[543];
  assign _EVAL_1136 = _EVAL_2019 & _EVAL_673;
  assign _EVAL_5438 = _EVAL_1145[605];
  assign _EVAL_5973 = _EVAL_921 & _EVAL_4477;
  assign _EVAL_424 = _EVAL_857 & _EVAL_1488;
  assign _EVAL_4844 = _EVAL_5074 & _EVAL_622;
  assign _EVAL_1529 = _EVAL_2868 & _EVAL_3487;
  assign _EVAL_2454 = _EVAL_713 & _EVAL_3379;
  assign _EVAL_4796 = _EVAL_3414 & _EVAL_2748;
  assign _EVAL_837 = _EVAL_4106 & _EVAL_1009;
  assign _EVAL_2127 = _EVAL_1625 & _EVAL_369;
  assign _EVAL_5157 = _EVAL_5074 & _EVAL_5201;
  assign _EVAL_302 = _EVAL_3650 & _EVAL_3379;
  assign _EVAL_5853 = _EVAL_3993 & _EVAL_882;
  assign _EVAL_6075 = _EVAL_4411 & _EVAL_673;
  assign _EVAL_4748 = _EVAL_594 & _EVAL_4664;
  assign _EVAL_2791 = _EVAL_4462 & _EVAL_1009;
  assign _EVAL_4966 = _EVAL_1136 & _EVAL_3154;
  assign _EVAL_4071 = _EVAL_3107 & _EVAL_6084;
  assign _EVAL_1209 = _EVAL_479 & _EVAL_369;
  assign _EVAL_2956 = _EVAL_4832 == 4'hf;
  assign _EVAL_3959 = _EVAL_1125 & _EVAL_3261;
  assign _EVAL_895 = _EVAL_1620 & _EVAL_1735;
  assign _EVAL_2325 = _EVAL_2100 & _EVAL_3487;
  assign _EVAL_5688 = _EVAL_1655 & _EVAL_3398;
  assign _EVAL_3719 = _EVAL_1145[527];
  assign _EVAL_5592 = _EVAL_3364 & _EVAL_3418;
  assign _EVAL_5245 = _EVAL_594 & _EVAL_1009;
  assign _EVAL_5402 = _EVAL_1446 & _EVAL_1488;
  assign _EVAL_231 = _EVAL_6059 & _EVAL_3418;
  assign _EVAL_5351 = _EVAL_4627 & _EVAL_574;
  assign _EVAL_4641 = _EVAL_1625 & _EVAL_1488;
  assign _EVAL_4186 = _EVAL_5561 & _EVAL_5838;
  assign _EVAL_3257 = _EVAL_4083 & _EVAL_847;
  assign _EVAL_3966 = _EVAL_961 & _EVAL_369;
  assign _EVAL_2069 = _EVAL_1542 & _EVAL_3487;
  assign _EVAL_3553 = _EVAL_2505 & _EVAL_3379;
  assign _EVAL_1938 = _EVAL_3364 & _EVAL_3154;
  assign _EVAL_5729 = _EVAL_4311 & _EVAL_587;
  assign _EVAL_5452 = _EVAL_2241 & _EVAL_369;
  assign _EVAL_1687 = _EVAL_2277 & _EVAL_1584;
  assign _EVAL_221 = _EVAL_4200 & _EVAL_3418;
  assign _EVAL_3132 = _EVAL_2254 & _EVAL_5543;
  assign _EVAL_922 = _EVAL_4627 & _EVAL_3509;
  assign _EVAL_2702 = _EVAL_6086 & _EVAL_2892;
  assign _EVAL_3710 = _EVAL_635 & _EVAL_3379;
  assign _EVAL_415 = _EVAL_3992 & _EVAL_5281;
  assign _EVAL_4512 = _EVAL_1145[597];
  assign _EVAL_3184 = ~_EVAL_5535;
  assign _EVAL_2133 = _EVAL_5598 & _EVAL_3418;
  assign _EVAL_4216 = _EVAL_1067 & _EVAL_3766;
  assign _EVAL_776 = _EVAL_251 & _EVAL_2969;
  assign _EVAL_3813 = _EVAL_4841 & _EVAL_882;
  assign _EVAL_342 = _EVAL_4045 & _EVAL_4077;
  assign _EVAL_5889 = _EVAL_1633 & _EVAL_3702;
  assign _EVAL_1634 = _EVAL_4141 & _EVAL_369;
  assign _EVAL_1620 = _EVAL_1707 & _EVAL_3379;
  assign _EVAL_3349 = _EVAL_5315 & _EVAL_5304;
  assign _EVAL_5006 = _EVAL_5561 & _EVAL_5582;
  assign _EVAL_5210 = _EVAL_4419 & _EVAL_3398;
  assign _EVAL_3924 = _EVAL_3689 & _EVAL_3702;
  assign _EVAL_5823 = _EVAL_1039 & _EVAL_847;
  assign _EVAL_3764 = _EVAL_4916 & _EVAL_5464;
  assign _EVAL_5303 = _EVAL_2241 & _EVAL_6084;
  assign _EVAL_1078 = _EVAL_251 & _EVAL_3702;
  assign _EVAL_4029 = _EVAL_4627 & _EVAL_2397;
  assign _EVAL_2925 = ~_EVAL_4051;
  assign _EVAL_1840 = ~_EVAL_1880;
  assign _EVAL_5938 = _EVAL_4085 & _EVAL_5260;
  assign _EVAL_905 = _EVAL_5087 & _EVAL_673;
  assign _EVAL_1198 = _EVAL_5922 == 4'hf;
  assign _EVAL_5866 = _EVAL_5074 & _EVAL_925;
  assign _EVAL_2673 = _EVAL_4627 & _EVAL_4817;
  assign _EVAL_3617 = _EVAL_4488 & _EVAL_3261;
  assign _EVAL_2317 = _EVAL_2106 & _EVAL_5543;
  assign _EVAL_3367 = _EVAL_6080 & _EVAL_1735;
  assign _EVAL_4792 = _EVAL_1446 & _EVAL_3702;
  assign _EVAL_3236 = _EVAL_1159[19:16];
  assign _EVAL_490 = _EVAL_4550 & _EVAL_2748;
  assign _EVAL_4016 = _EVAL_5206 & _EVAL_2956;
  assign _EVAL_3736 = _EVAL_5100 & _EVAL_4751;
  assign _EVAL_1816 = _EVAL_778 & _EVAL_587;
  assign _EVAL_1327 = _EVAL_5743 & _EVAL_4981;
  assign _EVAL_194 = _EVAL_1158 & _EVAL_3261;
  assign _EVAL_4577 = _EVAL_2433 & _EVAL_673;
  assign _EVAL_3588 = _EVAL_4507 & _EVAL_1198;
  assign _EVAL_248 = _EVAL_2106 & _EVAL_3702;
  assign _EVAL_5446 = _EVAL_4627 & _EVAL_3209;
  assign _EVAL_849 = _EVAL_2252 & _EVAL_3154;
  assign _EVAL_2502 = _EVAL_5054 & _EVAL_3261;
  assign _EVAL_3091 = _EVAL_2037 & _EVAL_2748;
  assign _EVAL_2449 = _EVAL_5370 & _EVAL_2748;
  assign _EVAL_4240 = _EVAL_3107 & _EVAL_369;
  assign _EVAL_5069 = _EVAL_4627 & _EVAL_3352;
  assign _EVAL_5018 = _EVAL_594 & _EVAL_587;
  assign _EVAL_4057 = _EVAL_581 & _EVAL_1198;
  assign _EVAL_1722 = _EVAL_534 & _EVAL_5850;
  assign _EVAL_3250 = _EVAL_2242 & _EVAL_369;
  assign _EVAL_4730 = _EVAL_5561 & _EVAL_3535;
  assign _EVAL_2437 = _EVAL_5819 & _EVAL_1290;
  assign _EVAL_2355 = _EVAL_1146 & _EVAL_3154;
  assign _EVAL_2167 = _EVAL_4783 & _EVAL_369;
  assign _EVAL_2762 = _EVAL_857 & _EVAL_2969;
  assign _EVAL_6055 = _EVAL_5068[535];
  assign _EVAL_5641 = ~_EVAL_3213;
  assign _EVAL_4411 = _EVAL_5561 & _EVAL_1144;
  assign _EVAL_860 = _EVAL_5386 & _EVAL_5075;
  assign _EVAL_638 = _EVAL_4525 & _EVAL_2382;
  assign _EVAL_1984 = _EVAL_1136 & _EVAL_882;
  assign _EVAL_4504 = ~_EVAL_3234;
  assign _EVAL_684 = _EVAL_4137 & _EVAL_3261;
  assign _EVAL_5078 = _EVAL_3945 > 4'h0;
  assign _EVAL_1086 = _EVAL_4093 & _EVAL_3154;
  assign _EVAL_4436 = _EVAL_3704 & _EVAL_2382;
  assign _EVAL_3342 = _EVAL_2192 & _EVAL_369;
  assign _EVAL_4120 = _EVAL_5561 & _EVAL_671;
  assign _EVAL_594 = _EVAL_6077 & _EVAL_673;
  assign _EVAL_4276 = _EVAL_5642 & _EVAL_5543;
  assign _EVAL_3176 = _EVAL_778 & _EVAL_4775;
  assign _EVAL_2296 = _EVAL_4499 & _EVAL_4109;
  assign _EVAL_5027 = _EVAL_831 & _EVAL_3702;
  assign _EVAL_4766 = _EVAL_3945 <= 4'h8;
  assign _EVAL_1833 = _EVAL_5411 & _EVAL_1555;
  assign _EVAL_5726 = _EVAL_4308 & _EVAL_3312;
  assign _EVAL_374 = _EVAL_1145[663];
  assign _EVAL_1179 = _EVAL_3935 & _EVAL_6084;
  assign _EVAL_637 = _EVAL_529 & _EVAL_3284;
  assign _EVAL_4346 = _EVAL_1281 & _EVAL_3313;
  assign _EVAL_1951 = _EVAL_2422 & _EVAL_4407;
  assign _EVAL_1146 = _EVAL_3478 & _EVAL_673;
  assign _EVAL_5902 = _EVAL_1370 & _EVAL_3418;
  assign _EVAL_1118 = _EVAL_5478 & _EVAL_3154;
  assign _EVAL_256 = ~_EVAL_603;
  assign _EVAL_5877 = _EVAL_1675 & _EVAL_3702;
  assign _EVAL_5568 = _EVAL_534 & _EVAL_1735;
  assign _EVAL_5416 = ~_EVAL_1618;
  assign _EVAL_3657 = _EVAL_3581 & _EVAL_1653;
  assign _EVAL_1847 = _EVAL_4567 & _EVAL_3398;
  assign _EVAL_3386 = _EVAL_3986 & _EVAL_1804;
  assign _EVAL_5102 = _EVAL_4192 & _EVAL_2748;
  assign _EVAL_1814 = _EVAL_4499 & _EVAL_2382;
  assign TLMonitor__EVAL_4 = _EVAL_25;
  assign _EVAL_1941 = _EVAL_4627 & _EVAL_1932;
  assign _EVAL_5433 = _EVAL_3226 & _EVAL_2382;
  assign _EVAL_3931 = _EVAL_5028 & _EVAL_5850;
  assign _EVAL_477 = _EVAL_1553 & _EVAL_1290;
  assign _EVAL_4983 = _EVAL_1125 & _EVAL_3398;
  assign _EVAL_5211 = ~_EVAL_2828;
  assign _EVAL_5133 = _EVAL_1361 & _EVAL_3398;
  assign _EVAL_5054 = _EVAL_3889 & _EVAL_673;
  assign _EVAL_3420 = _EVAL_626 ? 8'hff : 8'h0;
  assign _EVAL_1017 = _EVAL_5063 & _EVAL_4477;
  assign _EVAL_1667 = _EVAL_5074 & _EVAL_574;
  assign _EVAL_5693 = _EVAL_6075 & _EVAL_847;
  assign _EVAL_1793 = _EVAL_1876 & _EVAL_4477;
  assign _EVAL_1700 = _EVAL_5063 & _EVAL_3398;
  assign _EVAL_181 = _EVAL_1633 & _EVAL_369;
  assign _EVAL_5895 = _EVAL_1146 & _EVAL_3261;
  assign _EVAL_3691 = _EVAL_4783 & _EVAL_6084;
  assign _EVAL_6022 = _EVAL_4190 & _EVAL_3379;
  assign _EVAL_5090 = _EVAL_4909 & _EVAL_2320;
  assign _EVAL_829 = _EVAL_4745 & _EVAL_3154;
  assign _EVAL_771 = _EVAL_5994 & _EVAL_3154;
  assign _EVAL_1391 = _EVAL_3047 != 4'h0;
  assign _EVAL_515 = _EVAL_5184 & _EVAL_4664;
  assign _EVAL_1567 = _EVAL_984 & _EVAL_3284;
  assign _EVAL_1016 = _EVAL_5478 & _EVAL_3261;
  assign _EVAL_5243 = _EVAL_4627 & _EVAL_731;
  assign _EVAL_5753 = _EVAL_4671 != 4'h0;
  assign _EVAL_3595 = _EVAL_4563 & _EVAL_2424;
  assign _EVAL_2858 = _EVAL_2793 & _EVAL_4477;
  assign _EVAL_5003 = _EVAL_4757 & _EVAL_3154;
  assign _EVAL_4024 = _EVAL_5074 & _EVAL_1299;
  assign _EVAL_3852 = _EVAL_828 & _EVAL_5850;
  assign _EVAL_402 = _EVAL_888 & _EVAL_3379;
  assign _EVAL_779 = _EVAL_623 & _EVAL_369;
  assign _EVAL_2268 = _EVAL_5147 & _EVAL_3821;
  assign _EVAL_275 = _EVAL_4419 & _EVAL_847;
  assign _EVAL_3481 = _EVAL_3202 & _EVAL_6084;
  assign _EVAL_2963 = _EVAL_4627 & _EVAL_2480;
  assign _EVAL_4149 = _EVAL_1846 & _EVAL_3379;
  assign _EVAL_3228 = _EVAL_2251 & _EVAL_2969;
  assign _EVAL_5261 = _EVAL_1242 & _EVAL_3398;
  assign _EVAL_731 = _EVAL_1145[588];
  assign _EVAL_1175 = _EVAL_1145[529];
  assign _EVAL_3804 = _EVAL_5561 & _EVAL_2174;
  assign _EVAL_5110 = _EVAL_5398 & _EVAL_369;
  assign _EVAL_3744 = _EVAL_5148 & _EVAL_2969;
  assign _EVAL_2496 = _EVAL_3364 & _EVAL_4477;
  assign _EVAL_6026 = _EVAL_5074 & _EVAL_2008;
  assign _EVAL_584 = _EVAL_1658 & _EVAL_673;
  assign _EVAL_5347 = _EVAL_1625 & _EVAL_3702;
  assign _EVAL_3025 = _EVAL_2998 & _EVAL_3154;
  assign _EVAL_4692 = _EVAL_3540 & _EVAL_673;
  assign _EVAL_2436 = _EVAL_5618 & _EVAL_2969;
  assign _EVAL_2987 = _EVAL_3961 & _EVAL_2748;
  assign _EVAL_4353 = _EVAL_451 & _EVAL_3766;
  assign _EVAL_4706 = _EVAL_620 & _EVAL_3170;
  assign _EVAL_210 = _EVAL_1145[522];
  assign _EVAL_5208 = _EVAL_1854 & _EVAL_3418;
  assign _EVAL_5788 = _EVAL_2001 & _EVAL_3379;
  assign _EVAL_1214 = _EVAL_5998 & _EVAL_4751;
  assign _EVAL_2888 = ~_EVAL_236;
  assign _EVAL_4187 = _EVAL_460 & _EVAL_673;
  assign _EVAL_478 = ~_EVAL_4233;
  assign _EVAL_4434 = ~_EVAL_1287;
  assign _EVAL_3747 = _EVAL_3935 & _EVAL_369;
  assign _EVAL_4787 = _EVAL_1103 & _EVAL_2748;
  assign _EVAL_580 = _EVAL_905 & _EVAL_3261;
  assign _EVAL_1169 = _EVAL_751 & _EVAL_2424;
  assign _EVAL_1802 = _EVAL_4106 & _EVAL_587;
  assign _EVAL_5812 = _EVAL_4821 & _EVAL_3702;
  assign _EVAL_5912 = _EVAL_5561 & _EVAL_2216;
  assign _EVAL_5085 = _EVAL_3920 & _EVAL_1009;
  assign _EVAL_4803 = _EVAL_5705 & _EVAL_3702;
  assign _EVAL_2035 = _EVAL_5440 & _EVAL_3398;
  assign _EVAL_921 = _EVAL_532 & _EVAL_673;
  assign _EVAL_3264 = _EVAL_2753 & 22'h1fecc0;
  assign _EVAL_2222 = _EVAL_2260 & _EVAL_3418;
  assign _EVAL_1993 = _EVAL_1202 & _EVAL_3154;
  assign _EVAL_235 = _EVAL_2254 & _EVAL_369;
  assign _EVAL_1800 = _EVAL_3843 & _EVAL_1585;
  assign _EVAL_4206 = _EVAL_2868 & _EVAL_3261;
  assign _EVAL_3170 = _EVAL_4832 != 4'h0;
  assign _EVAL_5136 = _EVAL_5068[529];
  assign _EVAL_739 = _EVAL_1145[642];
  assign _EVAL_3896 = _EVAL_3322 & _EVAL_3284;
  assign _EVAL_2306 = _EVAL_1145[515];
  assign _EVAL_2432 = _EVAL_807 & _EVAL_1290;
  assign _EVAL_2846 = _EVAL_1865 & _EVAL_3418;
  assign _EVAL_3874 = ~_EVAL_1383;
  assign _EVAL_1369 = _EVAL_3928 & _EVAL_3261;
  assign _EVAL_1764 = _EVAL_799 & _EVAL_2969;
  assign _EVAL_4698 = _EVAL_4627 & _EVAL_936;
  assign _EVAL_4802 = _EVAL_1533 & _EVAL_3998;
  assign _EVAL_1638 = _EVAL_2242 & _EVAL_2424;
  assign _EVAL_5449 = _EVAL_4870 & _EVAL_5299;
  assign _EVAL_5116 = _EVAL_5561 & _EVAL_2281;
  assign _EVAL_179 = _EVAL_5608 & _EVAL_257;
  assign _EVAL_2553 = _EVAL_2550 & _EVAL_587;
  assign _EVAL_1789 = _EVAL_3220 & _EVAL_2748;
  assign TLMonitor__EVAL_13 = _EVAL_77;
  assign _EVAL_2834 = _EVAL_1675 & _EVAL_2969;
  assign _EVAL_3951 = _EVAL_4224 & _EVAL_4109;
  assign _EVAL_2985 = _EVAL_4462 & _EVAL_5289;
  assign _EVAL_428 = _EVAL_961 & _EVAL_2969;
  assign _EVAL_4951 = _EVAL_4106 & _EVAL_4775;
  assign _EVAL_4325 = _EVAL_5074 & _EVAL_2601;
  assign _EVAL_1724 = _EVAL_5077 & _EVAL_4477;
  assign _EVAL_1924 = _EVAL_523 == 8'hff;
  assign _EVAL_1037 = _EVAL_4053 & _EVAL_3223;
  assign _EVAL_2344 = _EVAL_4149 & _EVAL_2424;
  assign _EVAL_1715 = _EVAL_1960 & _EVAL_5753;
  assign _EVAL_5764 = _EVAL_961 & _EVAL_2748;
  assign _EVAL_3227 = _EVAL_4106 & _EVAL_3766;
  assign _EVAL_4976 = _EVAL_6021 & _EVAL_4931;
  assign TLMonitor__EVAL_9 = _EVAL_112;
  assign _EVAL_2411 = _EVAL_2100 & _EVAL_4477;
  assign _EVAL_4042 = _EVAL_392 & _EVAL_3379;
  assign _EVAL_4999 = _EVAL_5305 & _EVAL_5299;
  assign _EVAL_2718 = _EVAL_4596 & _EVAL_4664;
  assign _EVAL_704 = ~_EVAL_3962;
  assign _EVAL_4427 = _EVAL_1082 & _EVAL_2748;
  assign _EVAL_4563 = _EVAL_5566 & _EVAL_3379;
  assign _EVAL_4248 = _EVAL_4499 & _EVAL_3170;
  assign _EVAL_5573 = ~_EVAL_1342;
  assign _EVAL_3223 = ~_EVAL_1645;
  assign _EVAL_2299 = _EVAL_4965 & _EVAL_5776;
  assign _EVAL_5395 = _EVAL_4689 & _EVAL_4751;
  assign _EVAL_551 = _EVAL_5219 & _EVAL_3379;
  assign _EVAL_175 = _EVAL_5074 & _EVAL_4101;
  assign _EVAL_5708 = _EVAL_5074 & _EVAL_1562;
  assign _EVAL_2721 = _EVAL_2170 & _EVAL_5543;
  assign _EVAL_2960 = _EVAL_2346 & _EVAL_5168;
  assign _EVAL_3492 = _EVAL_4627 & _EVAL_1363;
  assign _EVAL_5542 = _EVAL_1570 & _EVAL_3379;
  assign _EVAL_4813 = _EVAL_2675 & _EVAL_2424;
  assign _EVAL_4245 = _EVAL_4618 & _EVAL_4775;
  assign _EVAL_2118 = _EVAL_5023 & _EVAL_4477;
  assign _EVAL_193 = ~_EVAL_3584;
  assign _EVAL_3694 = _EVAL_5068[520];
  assign _EVAL_5720 = _EVAL_1533 & _EVAL_3508;
  assign _EVAL_5825 = _EVAL_4795 & _EVAL_369;
  assign _EVAL_1628 = _EVAL_1649 & _EVAL_3702;
  assign _EVAL_4257 = _EVAL_5616 & _EVAL_3379;
  assign _EVAL_5941 = _EVAL_5246 & _EVAL_4477;
  assign _EVAL_1543 = _EVAL_5788 & _EVAL_5850;
  assign _EVAL_1213 = _EVAL_2516 & _EVAL_904;
  assign _EVAL_5977 = ~_EVAL_5916;
  assign _EVAL_3157 = ~_EVAL_3221;
  assign _EVAL_4833 = _EVAL_4577 & _EVAL_4775;
  assign _EVAL_5822 = _EVAL_617 & _EVAL_2424;
  assign _EVAL_348 = _EVAL_4974 & _EVAL_4109;
  assign _EVAL_751 = _EVAL_2135 & _EVAL_3379;
  assign _EVAL_5534 = _EVAL_4795 & _EVAL_1488;
  assign _EVAL_2284 = _EVAL_5795 & _EVAL_587;
  assign _EVAL_5784 = _EVAL_5074 & _EVAL_4306;
  assign _EVAL_6080 = _EVAL_4851 & _EVAL_3379;
  assign _EVAL_3575 = _EVAL_2998 & _EVAL_3398;
  assign _EVAL_2517 = _EVAL_1158 & _EVAL_3154;
  assign _EVAL_2387 = _EVAL_4627 & _EVAL_2044;
  assign _EVAL_5887 = _EVAL_4200 & _EVAL_4477;
  assign _EVAL_3052 = _EVAL_4629 & _EVAL_673;
  assign _EVAL_534 = _EVAL_600 & _EVAL_3379;
  assign _EVAL_1443 = ~_EVAL_4087;
  assign _EVAL_269 = _EVAL_2205 & _EVAL_1735;
  assign _EVAL_363 = _EVAL_2793 & _EVAL_882;
  assign _EVAL_5230 = ~_EVAL_546;
  assign _EVAL_3761 = _EVAL_1145[643];
  assign _EVAL_4212 = _EVAL_4836 & _EVAL_369;
  assign _EVAL_4138 = _EVAL_3421 & _EVAL_882;
  assign _EVAL_4651 = _EVAL_5068[533];
  assign _EVAL_508 = _EVAL_589 & _EVAL_3170;
  assign _EVAL_504 = _EVAL_1957 & _EVAL_3379;
  assign _EVAL_3547 = _EVAL_486 & _EVAL_369;
  assign _EVAL_1607 = _EVAL_1136 & _EVAL_3398;
  assign _EVAL_1064 = _EVAL_3202 & _EVAL_369;
  assign _EVAL_5648 = _EVAL_6033 & _EVAL_587;
  assign _EVAL_1675 = _EVAL_5492 & _EVAL_3379;
  assign _EVAL_4092 = _EVAL_1625 & _EVAL_6084;
  assign _EVAL_5544 = _EVAL_4314 & _EVAL_369;
  assign _EVAL_3774 = _EVAL_1067 & _EVAL_4775;
  assign _EVAL_952 = _EVAL_434 & _EVAL_4477;
  assign _EVAL_3610 = _EVAL_2192 & _EVAL_2748;
  assign _EVAL_4342 = _EVAL_3512 & _EVAL_1488;
  assign _EVAL_2163 = _EVAL_5370 & _EVAL_5543;
  assign _EVAL_1606 = _EVAL_2873 & _EVAL_2956;
  assign _EVAL_4974 = _EVAL_1167 & _EVAL_3379;
  assign _EVAL_3721 = _EVAL_1034 & _EVAL_1198;
  assign _EVAL_339 = ~_EVAL_1506;
  assign _EVAL_3651 = _EVAL_3437 & _EVAL_3379;
  assign _EVAL_951 = _EVAL_309 & _EVAL_5464;
  assign _EVAL_1570 = _EVAL_4627 & _EVAL_4259;
  assign _EVAL_4150 = _EVAL_857 & _EVAL_5543;
  assign _EVAL_5357 = _EVAL_5153 & _EVAL_3998;
  assign _EVAL_5400 = _EVAL_3476 & _EVAL_2424;
  assign _EVAL_3399 = _EVAL_538 & _EVAL_1488;
  assign _EVAL_4350 = _EVAL_1446 & _EVAL_2969;
  assign _EVAL_3009 = _EVAL_3651 & _EVAL_5543;
  assign _EVAL_2816 = _EVAL_4987 & _EVAL_3284;
  assign _EVAL_982 = _EVAL_5383 & _EVAL_369;
  assign _EVAL_4078 = _EVAL_869 & _EVAL_3379;
  assign _EVAL_2627 = _EVAL_2366 & _EVAL_2925;
  assign _EVAL_5834 = _EVAL_1149 & _EVAL_5543;
  assign _EVAL_3116 = _EVAL_3581 & _EVAL_5281;
  assign _EVAL_4678 = _EVAL_284 & _EVAL_2748;
  assign _EVAL_792 = _EVAL_5561 & _EVAL_234;
  assign _EVAL_4871 = _EVAL_3996 & _EVAL_1290;
  assign _EVAL_2955 = _EVAL_2251 & _EVAL_1488;
  assign _EVAL_1355 = _EVAL_5074 & _EVAL_3528;
  assign _EVAL_2426 = _EVAL_4627 & _EVAL_3719;
  assign _EVAL_1879 = _EVAL_3815 & _EVAL_4109;
  assign _EVAL_5893 = _EVAL_5708 & _EVAL_3379;
  assign _EVAL_3076 = _EVAL_4916 & _EVAL_3170;
  assign _EVAL_5642 = _EVAL_4597 & _EVAL_3379;
  assign _EVAL_1719 = _EVAL_5100 & _EVAL_4108;
  assign _EVAL_4365 = _EVAL_6051 & _EVAL_4109;
  assign _EVAL_1727 = _EVAL_5561 & _EVAL_2074;
  assign _EVAL_5016 = _EVAL_4627 & _EVAL_206;
  assign _EVAL_4669 = _EVAL_3920 & _EVAL_4775;
  assign _EVAL_1862 = _EVAL_5002 & _EVAL_4492;
  assign _EVAL_2731 = _EVAL_5599 & _EVAL_3379;
  assign _EVAL_5424 = ~_EVAL_5232;
  assign _EVAL_541 = ~_EVAL_3203;
  assign _EVAL_2645 = _EVAL_1281 & _EVAL_4788;
  assign _EVAL_1386 = _EVAL_5074 & _EVAL_2044;
  assign _EVAL_2371 = _EVAL_302 & _EVAL_369;
  assign _EVAL_1535 = _EVAL_5440 & _EVAL_3487;
  assign _EVAL_4831 = _EVAL_5561 & _EVAL_1464;
  assign _EVAL_3882 = _EVAL_1159[27:24];
  assign _EVAL_1533 = _EVAL_2370 & _EVAL_3379;
  assign _EVAL_2738 = _EVAL_6080 & _EVAL_2382;
  assign _EVAL_2821 = _EVAL_6033 & _EVAL_3766;
  assign _EVAL_1861 = _EVAL_3945 == 4'h8;
  assign _EVAL_2655 = _EVAL_5074 & _EVAL_4408;
  assign _EVAL_2930 = _EVAL_6080 & _EVAL_5464;
  assign _EVAL_2565 = ~_EVAL_1166;
  assign _EVAL_2106 = _EVAL_3267 & _EVAL_3379;
  assign _EVAL_2012 = _EVAL_3689 & _EVAL_369;
  assign _EVAL_5843 = _EVAL_2471 & _EVAL_3487;
  assign _EVAL_4967 = _EVAL_1136 & _EVAL_3487;
  assign _EVAL_1281 = _EVAL_3909 & _EVAL_673;
  assign _EVAL_2071 = ~_EVAL_896;
  assign _EVAL_1776 = _EVAL_4974 & _EVAL_4751;
  assign _EVAL_5919 = _EVAL_1649 & _EVAL_2969;
  assign _EVAL_4841 = _EVAL_2131 & _EVAL_673;
  assign _EVAL_1772 = _EVAL_2170 & _EVAL_369;
  assign _EVAL_2187 = _EVAL_5162 & _EVAL_3702;
  assign _EVAL_985 = _EVAL_1103 & _EVAL_369;
  assign _EVAL_4737 = _EVAL_5054 & _EVAL_3154;
  assign _EVAL_2033 = _EVAL_688 & _EVAL_3487;
  assign _EVAL_1905 = _EVAL_1875 & _EVAL_1631;
  assign _EVAL_347 = _EVAL_1145[523];
  assign _EVAL_2224 = _EVAL_1396 & _EVAL_3558;
  assign _EVAL_6090 = _EVAL_2252 & _EVAL_3398;
  assign _EVAL_5594 = _EVAL_1361 & _EVAL_847;
  assign _EVAL_1455 = _EVAL_1971 & _EVAL_6084;
  assign _EVAL_2748 = _EVAL_1316[16];
  assign _EVAL_5431 = _EVAL_3837 & _EVAL_2748;
  assign _EVAL_6038 = _EVAL_4044 & _EVAL_3261;
  assign _EVAL_804 = _EVAL_2471 & _EVAL_3398;
  assign _EVAL_5959 = _EVAL_6059 & _EVAL_847;
  assign _EVAL_345 = _EVAL_3512 & _EVAL_5543;
  assign _EVAL_1804 = ~_EVAL_355;
  assign _EVAL_4027 = _EVAL_4807 & _EVAL_5496;
  assign _EVAL_4405 = _EVAL_1593 & _EVAL_4872;
  assign _EVAL_2193 = _EVAL_4567 & _EVAL_847;
  assign _EVAL_1109 = _EVAL_2005 & _EVAL_3702;
  assign _EVAL_4811 = _EVAL_5193 & _EVAL_2424;
  assign _EVAL_4996 = _EVAL_1960 & _EVAL_4664;
  assign _EVAL_3525 = _EVAL_1158 & _EVAL_4477;
  assign _EVAL_422 = _EVAL_2972 & _EVAL_1009;
  assign _EVAL_2442 = _EVAL_935 & _EVAL_3702;
  assign _EVAL_5561 = _EVAL_970 & Queue__EVAL_2;
  assign _EVAL_5362 = _EVAL_3476 & _EVAL_6084;
  assign _EVAL_1579 = _EVAL_3689 & _EVAL_1488;
  assign _EVAL_1180 = _EVAL_5184 & _EVAL_1290;
  assign _EVAL_460 = _EVAL_5561 & _EVAL_747;
  assign _EVAL_5036 = _EVAL_5561 & _EVAL_5203;
  assign _EVAL_1142 = _EVAL_3887 & _EVAL_2208;
  assign _EVAL_5857 = _EVAL_623 & _EVAL_2424;
  assign _EVAL_2195 = _EVAL_1920 & _EVAL_3418;
  assign _EVAL_370 = _EVAL_3981 & _EVAL_3487;
  assign _EVAL_4693 = _EVAL_4757 & _EVAL_4477;
  assign _EVAL_4207 = _EVAL_984 & _EVAL_1198;
  assign _EVAL_2647 = _EVAL_623 & _EVAL_6084;
  assign _EVAL_884 = _EVAL_1312 & _EVAL_3702;
  assign _EVAL_3432 = _EVAL_309 & _EVAL_2382;
  assign _EVAL_610 = _EVAL_5074 & _EVAL_464;
  assign _EVAL_227 = _EVAL_1145[587];
  assign _EVAL_1839 = _EVAL_4742 & _EVAL_5927;
  assign _EVAL_3306 = _EVAL_4419 & _EVAL_3154;
  assign _EVAL_764 = _EVAL_735 & _EVAL_5850;
  assign _EVAL_3312 = ~_EVAL_1131;
  assign _EVAL_1413 = _EVAL_1234 & _EVAL_369;
  assign _EVAL_1689 = _EVAL_3995 & _EVAL_3379;
  assign _EVAL_2608 = _EVAL_4351 & _EVAL_369;
  assign _EVAL_5173 = _EVAL_5068[547];
  assign _EVAL_4697 = _EVAL_5561 & _EVAL_4566;
  assign _EVAL_2945 = _EVAL_1159[31:25];
  assign _EVAL_481 = _EVAL_4618 & _EVAL_5289;
  assign TLMonitor__EVAL_3 = _EVAL_124;
  assign _EVAL_5790 = _EVAL_3706 & _EVAL_2969;
  assign _EVAL_3142 = _EVAL_5342 & _EVAL_5299;
  assign _EVAL_1406 = _EVAL_362 & _EVAL_4664;
  assign _EVAL_2245 = _EVAL_1500 & _EVAL_4477;
  assign _EVAL_2903 = _EVAL_1370 & _EVAL_3487;
  assign _EVAL_3995 = _EVAL_4627 & _EVAL_2405;
  assign _EVAL_4299 = _EVAL_3346 & _EVAL_882;
  assign _EVAL_362 = _EVAL_5317 & _EVAL_673;
  assign TLMonitor__EVAL_7 = _EVAL_24;
  assign _EVAL_4842 = _EVAL_4661 & _EVAL_587;
  assign _EVAL_3649 = _EVAL_5705 & _EVAL_6084;
  assign _EVAL_4795 = _EVAL_5069 & _EVAL_3379;
  assign _EVAL_1302 = _EVAL_302 & _EVAL_6084;
  assign _EVAL_5355 = _EVAL_857 & _EVAL_2424;
  assign _EVAL_4568 = _EVAL_589 & _EVAL_2382;
  assign _EVAL_2367 = _EVAL_5561 & _EVAL_3365;
  assign _EVAL_4605 = _EVAL_1145[661];
  assign _EVAL_4108 = _EVAL_2798 != 4'h0;
  assign _EVAL_4800 = _EVAL_4755 & _EVAL_5464;
  assign _EVAL_3241 = _EVAL_4507 & _EVAL_5299;
  assign _EVAL_1649 = _EVAL_4720 & _EVAL_3379;
  assign _EVAL_2682 = _EVAL_4577 & _EVAL_1290;
  assign _EVAL_3835 = _EVAL_4224 & _EVAL_5850;
  assign _EVAL_3524 = _EVAL_1256 & _EVAL_3379;
  assign _EVAL_809 = _EVAL_5819 & _EVAL_3766;
  assign _EVAL_4281 = _EVAL_1625 & _EVAL_5543;
  assign _EVAL_778 = _EVAL_2323 & _EVAL_673;
  assign _EVAL_3949 = _EVAL_5100 & _EVAL_2382;
  assign _EVAL_5668 = _EVAL_5427 & _EVAL_3487;
  assign _EVAL_4373 = _EVAL_2177 & _EVAL_3548;
  assign _EVAL_5033 = _EVAL_2778 & _EVAL_3015;
  assign _EVAL_392 = _EVAL_4627 & _EVAL_3329;
  assign _EVAL_4573 = _EVAL_2725 & _EVAL_3398;
  assign _EVAL_3070 = _EVAL_2772 & _EVAL_3379;
  assign _EVAL_3186 = _EVAL_1145[533];
  assign _EVAL_4916 = _EVAL_4698 & _EVAL_3379;
  assign _EVAL_5740 = _EVAL_2292 & _EVAL_5464;
  assign _EVAL_825 = _EVAL_4836 & _EVAL_3388;
  assign _EVAL_2208 = ~_EVAL_1331;
  assign _EVAL_5795 = _EVAL_2597 & _EVAL_673;
  assign _EVAL_3833 = _EVAL_3928 & _EVAL_3154;
  assign _EVAL_1902 = _EVAL_4745 & _EVAL_4477;
  assign _EVAL_2364 = _EVAL_381 & _EVAL_876;
  assign _EVAL_4825 = _EVAL_5068[525];
  assign _EVAL_4294 = _EVAL_1689 & _EVAL_3702;
  assign _EVAL_5842 = _EVAL_5440 & _EVAL_882;
  assign _EVAL_711 = _EVAL_4661 & _EVAL_3766;
  assign _EVAL_2946 = _EVAL_1125 & _EVAL_3487;
  assign _EVAL_787 = _EVAL_5074 & _EVAL_1932;
  assign _EVAL_2833 = _EVAL_4888 & _EVAL_2748;
  assign _EVAL_3084 = _EVAL_6075 & _EVAL_3487;
  assign _EVAL_2720 = _EVAL_4254 & _EVAL_1290;
  assign _EVAL_5213 = _EVAL_2192 & _EVAL_2424;
  assign _EVAL_6017 = _EVAL_4322 & _EVAL_2748;
  assign _EVAL_322 = _EVAL_4596 & _EVAL_5289;
  assign _EVAL_3928 = _EVAL_4186 & _EVAL_673;
  assign _EVAL_2175 = _EVAL_584 & _EVAL_3313;
  assign _EVAL_4330 = _EVAL_3220 & _EVAL_3702;
  assign _EVAL_1639 = _EVAL_6007 & _EVAL_4477;
  assign _EVAL_5470 = _EVAL_4689 & _EVAL_5464;
  assign _EVAL_2082 = _EVAL_1145[611];
  assign _EVAL_2844 = _EVAL_6032 & _EVAL_369;
  assign _EVAL_4794 = _EVAL_1146 & _EVAL_4477;
  assign _EVAL_4110 = _EVAL_620 & _EVAL_4751;
  assign _EVAL_2514 = _EVAL_1145[514];
  assign _EVAL_5848 = _EVAL_3920 & _EVAL_4664;
  assign _EVAL_627 = _EVAL_4661 & _EVAL_4664;
  assign _EVAL_1137 = _EVAL_6007 & _EVAL_3154;
  assign _EVAL_4323 = _EVAL_965 & _EVAL_1290;
  assign _EVAL_3054 = _EVAL_4627 & _EVAL_4001;
  assign _EVAL_1467 = _EVAL_1364 & _EVAL_2956;
  assign _EVAL_5260 = ~_EVAL_3634;
  assign TLMonitor__EVAL_0 = Queue__EVAL_11;
  assign _EVAL_4938 = _EVAL_3364 & _EVAL_3261;
  assign _EVAL_2134 = _EVAL_5370 & _EVAL_2424;
  assign _EVAL_3400 = _EVAL_799 & _EVAL_2424;
  assign _EVAL_3506 = _EVAL_1446 & _EVAL_6084;
  assign _EVAL_2897 = _EVAL_5074 & _EVAL_6008;
  assign _EVAL_3447 = ~_EVAL_2203;
  assign _EVAL_1767 = _EVAL_3629 & _EVAL_4163;
  assign _EVAL_5686 = _EVAL_263 & _EVAL_5299;
  assign _EVAL_2217 = _EVAL_623 & _EVAL_2969;
  assign _EVAL_3069 = _EVAL_1311 & _EVAL_3663;
  assign _EVAL_2073 = _EVAL_2902 & _EVAL_369;
  assign _EVAL_3730 = _EVAL_3837 & _EVAL_6084;
  assign _EVAL_1625 = _EVAL_6069 & _EVAL_3379;
  assign _EVAL_4857 = _EVAL_4488 & _EVAL_3154;
  assign _EVAL_5827 = _EVAL_2753[5];
  assign _EVAL_2990 = _EVAL_1689 & _EVAL_2424;
  assign _EVAL_391 = _EVAL_1960 & _EVAL_3766;
  assign _EVAL_5017 = _EVAL_1370 & _EVAL_847;
  assign _EVAL_4363 = _EVAL_5305 & _EVAL_1198;
  assign _EVAL_954 = ~_EVAL_2381;
  assign _EVAL_755 = _EVAL_4311 & _EVAL_5753;
  assign _EVAL_3845 = _EVAL_6026 & _EVAL_3379;
  assign _EVAL_5291 = _EVAL_3624 & _EVAL_1488;
  assign _EVAL_5234 = _EVAL_277 & _EVAL_5194;
  assign _EVAL_4023 = _EVAL_5998 & _EVAL_4108;
  assign _EVAL_4408 = _EVAL_1145[600];
  assign _EVAL_1684 = _EVAL_3171 & _EVAL_4279;
  assign _EVAL_259 = _EVAL_3965 & _EVAL_4570;
  assign _EVAL_3770 = _EVAL_4078 & _EVAL_1488;
  assign _EVAL_2117 = _EVAL_1145[545];
  assign _EVAL_5559 = _EVAL_3476 & _EVAL_5543;
  assign _EVAL_1913 = _EVAL_4577 & _EVAL_587;
  assign _EVAL_2524 = _EVAL_2907 & _EVAL_6084;
  assign _EVAL_1196 = _EVAL_5193 & _EVAL_6084;
  assign _EVAL_1176 = _EVAL_4627 & _EVAL_931;
  assign _EVAL_6008 = _EVAL_1145[651];
  assign _EVAL_3858 = _EVAL_3981 & _EVAL_3261;
  assign _EVAL_2232 = _EVAL_4627 & _EVAL_4086;
  assign _EVAL_280 = _EVAL_623 & _EVAL_2748;
  assign _EVAL_5946 = _EVAL_6075 & _EVAL_882;
  assign _EVAL_2079 = ~_EVAL_1301;
  assign _EVAL_5368 = _EVAL_5478 & _EVAL_3487;
  assign _EVAL_1305 = _EVAL_2731 & _EVAL_2748;
  assign _EVAL_1341 = _EVAL_1039 & _EVAL_3154;
  assign _EVAL_3201 = _EVAL_774 & _EVAL_6084;
  assign _EVAL_3920 = _EVAL_1523 & _EVAL_673;
  assign _EVAL_4470 = _EVAL_5676 & _EVAL_4477;
  assign _EVAL_6085 = _EVAL_362 & _EVAL_4775;
  assign _EVAL_2550 = _EVAL_908 & _EVAL_673;
  assign _EVAL_3235 = _EVAL_5077 & _EVAL_3261;
  assign _EVAL_1296 = _EVAL_3632 & _EVAL_4108;
  assign TLMonitor__EVAL_8 = Queue__EVAL_0;
  assign _EVAL_4106 = _EVAL_5454 & _EVAL_673;
  assign _EVAL_3113 = _EVAL_4627 & _EVAL_2991;
  assign _EVAL_2459 = _EVAL_4200 & _EVAL_3487;
  assign _EVAL_3138 = _EVAL_2121 & _EVAL_3487;
  assign _EVAL_5445 = _EVAL_1475 == 8'hff;
  assign _EVAL_5023 = _EVAL_4263 & _EVAL_673;
  assign _EVAL_2443 = _EVAL_1745 & _EVAL_4751;
  assign _EVAL_1709 = _EVAL_356 & _EVAL_4961;
  assign _EVAL_1994 = _EVAL_251 & _EVAL_2424;
  assign _EVAL_965 = _EVAL_2076 & _EVAL_673;
  assign _EVAL_5167 = _EVAL_5676 & _EVAL_3418;
  assign _EVAL_1049 = _EVAL_2585 & _EVAL_3418;
  assign _EVAL_4814 = _EVAL_4577 & _EVAL_4664;
  assign _EVAL_617 = _EVAL_5461 & _EVAL_3379;
  assign _EVAL_4759 = _EVAL_4202 & _EVAL_4788;
  assign _EVAL_3261 = _EVAL_2945 != 7'h0;
  assign _EVAL_2378 = _EVAL_2242 & _EVAL_2748;
  assign _EVAL_241 = _EVAL_1145[534];
  assign _EVAL_3078 = _EVAL_2873 & _EVAL_5299;
  assign _EVAL_1910 = _EVAL_4078 & _EVAL_2969;
  assign _EVAL_4020 = _EVAL_4257 & _EVAL_2748;
  assign _EVAL_4671 = _EVAL_1159[3:0];
  assign _EVAL_1158 = _EVAL_4713 & _EVAL_673;
  assign _EVAL_3902 = _EVAL_3815 & _EVAL_3170;
  assign _EVAL_5744 = _EVAL_1745 & _EVAL_2382;
  assign _EVAL_975 = _EVAL_1854 & _EVAL_3154;
  assign _EVAL_2110 = _EVAL_857 & _EVAL_369;
  assign _EVAL_4979 = _EVAL_688 & _EVAL_3418;
  assign _EVAL_2455 = _EVAL_4627 & _EVAL_2008;
  assign _EVAL_1691 = _EVAL_6051 & _EVAL_5464;
  assign _EVAL_2149 = _EVAL_3845 & _EVAL_2956;
  assign _EVAL_1769 = _EVAL_2592 & _EVAL_5543;
  assign _EVAL_4731 = _EVAL_2251 & _EVAL_369;
  assign _EVAL_4585 = _EVAL_5705 & _EVAL_1488;
  assign _EVAL_744 = _EVAL_3574 & _EVAL_3508;
  assign _EVAL_5524 = _EVAL_5854 & _EVAL_2956;
  assign _EVAL_5050 = _EVAL_5068[536];
  assign _EVAL_480 = _EVAL_2292 & _EVAL_4108;
  assign _EVAL_383 = _EVAL_1316[6:5];
  assign _EVAL_4879 = _EVAL_1500 & _EVAL_3154;
  assign _EVAL_3856 = _EVAL_921 & _EVAL_3261;
  assign _EVAL_3387 = _EVAL_1149 & _EVAL_2969;
  assign _EVAL_2401 = _EVAL_3130 & _EVAL_1488;
  assign _EVAL_2688 = _EVAL_1316[7:4];
  assign _EVAL_1660 = _EVAL_4488 & _EVAL_4477;
  assign _EVAL_4866 = _EVAL_1763 > 4'h8;
  assign _EVAL_1516 = ~_EVAL_6098;
  assign _EVAL_5766 = _EVAL_1491 & _EVAL_673;
  assign _EVAL_1297 = _EVAL_6007 & _EVAL_3487;
  assign _EVAL_1065 = _EVAL_4627 & _EVAL_4601;
  assign _EVAL_1633 = _EVAL_5970 & _EVAL_3379;
  assign _EVAL_4654 = _EVAL_3322 & _EVAL_2956;
  assign _EVAL_4564 = _EVAL_1145[608];
  assign _EVAL_5986 = _EVAL_3216 & _EVAL_4477;
  assign _EVAL_1604 = _EVAL_1145[538];
  assign _EVAL_1521 = _EVAL_5528 & _EVAL_5753;
  assign _EVAL_3226 = _EVAL_3867 & _EVAL_3379;
  assign _EVAL_5779 = _EVAL_4627 & _EVAL_1558;
  assign _EVAL_169 = _EVAL_3928 & _EVAL_3487;
  assign _EVAL_5317 = _EVAL_5561 & _EVAL_2693;
  assign _EVAL_670 = _EVAL_538 & _EVAL_6084;
  assign _EVAL_4133 = _EVAL_5353 & _EVAL_2969;
  assign _EVAL_802 = _EVAL_1240 & _EVAL_726;
  assign _EVAL_612 = _EVAL_5100 & _EVAL_5850;
  assign _EVAL_4702 = _EVAL_5028 & _EVAL_4108;
  assign _EVAL_798 = _EVAL_5054 & _EVAL_882;
  assign _EVAL_4854 = ~_EVAL_3194;
  assign _EVAL_1085 = _EVAL_4078 & _EVAL_3702;
  assign _EVAL_1167 = _EVAL_4627 & _EVAL_5837;
  assign _EVAL_3904 = _EVAL_3364 & _EVAL_3487;
  assign _EVAL_1708 = _EVAL_309 & _EVAL_4108;
  assign _EVAL_5035 = _EVAL_4841 & _EVAL_3487;
  assign _EVAL_375 = _EVAL_5074 & _EVAL_5760;
  assign _EVAL_1371 = _EVAL_2877 & _EVAL_2424;
  assign _EVAL_3994 = _EVAL_298 & _EVAL_3508;
  assign _EVAL_1389 = _EVAL_5561 & _EVAL_3466;
  assign _EVAL_4680 = _EVAL_1393 & _EVAL_5543;
  assign _EVAL_1723 = _EVAL_799 & _EVAL_5543;
  assign _EVAL_3680 = _EVAL_2260 & _EVAL_3487;
  assign _EVAL_5067 = _EVAL_1745 & _EVAL_5850;
  assign _EVAL_334 = _EVAL_1316[31:24];
  assign _EVAL_4495 = _EVAL_1159[7:1];
  assign _EVAL_1818 = _EVAL_4222 & _EVAL_882;
  assign _EVAL_1360 = _EVAL_799 & _EVAL_6084;
  assign _EVAL_1966 = _EVAL_5074 & _EVAL_6076;
  assign _EVAL_6087 = _EVAL_2179 & _EVAL_3379;
  assign _EVAL_552 = ~_EVAL_5479;
  assign _EVAL_1784 = _EVAL_4841 & _EVAL_3261;
  assign _EVAL_3251 = _EVAL_5869 & _EVAL_3261;
  assign _EVAL_4877 = ~_EVAL_4065;
  assign _EVAL_440 = _EVAL_1500 & _EVAL_3418;
  assign _EVAL_3490 = _EVAL_4627 & _EVAL_5625;
  assign _EVAL_956 = _EVAL_5427 & _EVAL_882;
  assign _EVAL_3050 = _EVAL_3476 & _EVAL_2969;
  assign _EVAL_4399 = _EVAL_965 & _EVAL_1009;
  assign _EVAL_1062 = _EVAL_4689 & _EVAL_4108;
  assign _EVAL_1420 = _EVAL_1865 & _EVAL_3398;
  assign _EVAL_4028 = _EVAL_5074 & _EVAL_227;
  assign _EVAL_2769 = _EVAL_623 & _EVAL_1488;
  assign _EVAL_2191 = _EVAL_6059 & _EVAL_3261;
  assign _EVAL_3910 = _EVAL_5370 & _EVAL_6084;
  assign _EVAL_1411 = _EVAL_1145[525];
  assign _EVAL_4736 = _EVAL_5561 & _EVAL_3944;
  assign _EVAL_3156 = _EVAL_5700 & _EVAL_3379;
  assign _EVAL_5488 = _EVAL_1136 & _EVAL_4477;
  assign _EVAL_3740 = _EVAL_5561 & _EVAL_2394;
  assign _EVAL_2480 = _EVAL_1145[583];
  assign _EVAL_2464 = _EVAL_1281 & _EVAL_1009;
  assign _EVAL_1071 = _EVAL_751 & _EVAL_5543;
  assign _EVAL_2881 = _EVAL_298 & _EVAL_2382;
  assign _EVAL_2235 = _EVAL_5561 & _EVAL_4825;
  assign _EVAL_1743 = _EVAL_2592 & _EVAL_2748;
  assign _EVAL_3413 = ~_EVAL_4103;
  assign _EVAL_3151 = _EVAL_4856 & _EVAL_2969;
  assign _EVAL_3712 = _EVAL_5074 & _EVAL_5867;
  assign _EVAL_1025 = _EVAL_4149 & _EVAL_6084;
  assign _EVAL_949 = _EVAL_124[3];
  assign _EVAL_233 = _EVAL_5184 & _EVAL_3766;
  assign _EVAL_1741 = _EVAL_4755 & _EVAL_3170;
  assign _EVAL_168 = _EVAL_2065 & _EVAL_2362;
  assign _EVAL_3403 = _EVAL_1633 & _EVAL_5543;
  assign _EVAL_260 = _EVAL_688 & _EVAL_847;
  assign _EVAL_5122 = _EVAL_451 & _EVAL_4160;
  assign _EVAL_3822 = _EVAL_1622 & _EVAL_4775;
  assign _EVAL_845 = _EVAL_1145[541];
  assign _EVAL_3785 = _EVAL_4692 & _EVAL_3487;
  assign _EVAL_5100 = _EVAL_1996 & _EVAL_3379;
  assign _EVAL_2452 = _EVAL_2877 & _EVAL_1488;
  assign _EVAL_5955 = _EVAL_1689 & _EVAL_6084;
  assign _EVAL_2931 = _EVAL_3859 & _EVAL_3284;
  assign _EVAL_831 = _EVAL_5988 & _EVAL_3379;
  assign _EVAL_2399 = _EVAL_1620 & _EVAL_3170;
  assign _EVAL_4315 = _EVAL_251 & _EVAL_6084;
  assign _EVAL_4043 = _EVAL_4627 & _EVAL_1596;
  assign _EVAL_5246 = _EVAL_3075 & _EVAL_673;
  assign _EVAL_5707 = _EVAL_5869 & _EVAL_882;
  assign _EVAL_3238 = _EVAL_309 & _EVAL_3170;
  assign _EVAL_3581 = _EVAL_5866 & _EVAL_3379;
  assign _EVAL_2059 = _EVAL_3632 & _EVAL_5850;
  assign _EVAL_3700 = _EVAL_4042 & _EVAL_3508;
  assign _EVAL_3178 = _EVAL_4563 & _EVAL_2969;
  assign _EVAL_4686 = ~_EVAL_3374;
  assign _EVAL_3072 = _EVAL_3920 & _EVAL_5289;
  assign _EVAL_5618 = _EVAL_2305 & _EVAL_3379;
  assign _EVAL_4072 = _EVAL_4093 & _EVAL_3398;
  assign _EVAL_3815 = _EVAL_1424 & _EVAL_3379;
  assign _EVAL_5306 = _EVAL_3188 & _EVAL_5753;
  assign _EVAL_2469 = _EVAL_3706 & _EVAL_5543;
  assign _EVAL_876 = ~_EVAL_4922;
  assign _EVAL_5976 = _EVAL_3624 & _EVAL_2748;
  assign _EVAL_4104 = _EVAL_3945 < 4'h8;
  assign _EVAL_5810 = _EVAL_5193 & _EVAL_2969;
  assign _EVAL_3869 = _EVAL_5816 & _EVAL_3998;
  assign _EVAL_237 = _EVAL_5192 & _EVAL_5543;
  assign _EVAL_1594 = _EVAL_5155 & _EVAL_369;
  assign _EVAL_4114 = _EVAL_1145[519];
  assign _EVAL_1728 = _EVAL_2988 & _EVAL_5158;
  assign _EVAL_1338 = _EVAL_4141 & _EVAL_2969;
  assign _EVAL_4022 = _EVAL_5427 & _EVAL_3261;
  assign _EVAL_6048 = _EVAL_4783 & _EVAL_2748;
  assign _EVAL_4219 = _EVAL_3174 & _EVAL_3379;
  assign _EVAL_3282 = _EVAL_2842 & _EVAL_5299;
  assign _EVAL_314 = _EVAL_4141 & _EVAL_1488;
  assign _EVAL_620 = _EVAL_3281 & _EVAL_3379;
  assign _EVAL_4160 = _EVAL_5000 != 8'h0;
  assign _EVAL_3002 = _EVAL_5132 & _EVAL_3261;
  assign _EVAL_3216 = _EVAL_5510 & _EVAL_673;
  assign _EVAL_4570 = ~_EVAL_661;
  assign _EVAL_1322 = _EVAL_1202 & _EVAL_3418;
  assign _EVAL_708 = _EVAL_302 & _EVAL_2424;
  assign _EVAL_2939 = _EVAL_3421 & _EVAL_3398;
  assign _EVAL_2064 = _EVAL_2725 & _EVAL_3487;
  assign _EVAL_5461 = _EVAL_4627 & _EVAL_4703;
  assign _EVAL_2921 = ~_EVAL_5190;
  assign _EVAL_1047 = _EVAL_4944 & _EVAL_3413;
  assign _EVAL_257 = ~_EVAL_3589;
  assign _EVAL_5750 = _EVAL_4311 & _EVAL_5289;
  assign _EVAL_4630 = _EVAL_4627 & _EVAL_2695;
  assign _EVAL_5152 = _EVAL_3787 & _EVAL_5753;
  assign _EVAL_2460 = _EVAL_965 & _EVAL_4160;
  assign _EVAL_5760 = _EVAL_1145[657];
  assign _EVAL_5206 = _EVAL_3562 & _EVAL_3379;
  assign _EVAL_3480 = _EVAL_5246 & _EVAL_3154;
  assign _EVAL_4203 = _EVAL_905 & _EVAL_3487;
  assign _EVAL_2014 = _EVAL_6032 & _EVAL_2424;
  assign _EVAL_5663 = _EVAL_4235 & _EVAL_5543;
  assign _EVAL_1105 = _EVAL_2753[1];
  assign _EVAL_279 = _EVAL_807 & _EVAL_1009;
  assign _EVAL_4744 = _EVAL_4141 & _EVAL_6084;
  assign _EVAL_5341 = _EVAL_584 & _EVAL_4160;
  assign _EVAL_4329 = _EVAL_1917 & _EVAL_5814;
  assign _EVAL_4761 = _EVAL_2592 & _EVAL_2969;
  assign _EVAL_1108 = _EVAL_1344 & _EVAL_3398;
  assign _EVAL_4130 = _EVAL_4351 & _EVAL_2748;
  assign _EVAL_5630 = _EVAL_2192 & _EVAL_5543;
  assign _EVAL_3210 = _EVAL_1145[650];
  assign _EVAL_4666 = _EVAL_1730 & _EVAL_339;
  assign _EVAL_5486 = _EVAL_5521 & _EVAL_2950;
  assign _EVAL_2027 = _EVAL_1655 & _EVAL_3487;
  assign _EVAL_2476 = _EVAL_1067 & _EVAL_1009;
  assign _EVAL_5917 = _EVAL_2753[0];
  assign _EVAL_3381 = _EVAL_2335 & _EVAL_2956;
  assign _EVAL_1384 = _EVAL_5819 & _EVAL_5289;
  assign _EVAL_944 = _EVAL_5705 & _EVAL_2969;
  assign _EVAL_4726 = _EVAL_5077 & _EVAL_3154;
  assign _EVAL_318 = ~_EVAL_2847;
  assign _EVAL_686 = _EVAL_4462 & _EVAL_4664;
  assign _EVAL_1526 = _EVAL_2251 & _EVAL_6084;
  assign _EVAL_1102 = _EVAL_4257 & _EVAL_369;
  assign _EVAL_4773 = _EVAL_6032 & _EVAL_6084;
  assign _EVAL_2230 = _EVAL_3476 & _EVAL_1488;
  assign _EVAL_4529 = _EVAL_3451 & _EVAL_3418;
  assign _EVAL_5370 = _EVAL_5242 & _EVAL_3379;
  assign _EVAL_5381 = _EVAL_1082 & _EVAL_369;
  assign _EVAL_2453 = _EVAL_3996 & _EVAL_4664;
  assign _EVAL_5528 = _EVAL_1058 & _EVAL_673;
  assign _EVAL_5586 = _EVAL_2607 & _EVAL_1198;
  assign _EVAL_1079 = _EVAL_4254 & _EVAL_4775;
  assign _EVAL_2075 = _EVAL_594 & _EVAL_5753;
  assign _EVAL_5081 = _EVAL_407 & _EVAL_5543;
  assign _EVAL_2789 = _EVAL_5184 & _EVAL_5753;
  assign _EVAL_3453 = _EVAL_402 & _EVAL_5299;
  assign _EVAL_748 = _EVAL_309 & _EVAL_4109;
  assign _EVAL_2735 = _EVAL_2702 & _EVAL_5445;
  assign _EVAL_4099 = _EVAL_3844 & _EVAL_3702;
  assign _EVAL_4690 = _EVAL_5162 & _EVAL_5543;
  assign _EVAL_1395 = ~_EVAL_3789;
  assign _EVAL_4845 = _EVAL_589 & _EVAL_4109;
  assign _EVAL_3725 = _EVAL_2192 & _EVAL_2969;
  assign _EVAL_1290 = _EVAL_4213 != 4'h0;
  assign _EVAL_3402 = _EVAL_5074 & _EVAL_5438;
  assign _EVAL_816 = _EVAL_5148 & _EVAL_5543;
  assign _EVAL_4649 = _EVAL_778 & _EVAL_5753;
  assign _EVAL_2972 = _EVAL_5904 & _EVAL_673;
  assign _EVAL_2044 = _EVAL_1145[593];
  assign _EVAL_3540 = _EVAL_5561 & _EVAL_5782;
  assign _EVAL_4033 = _EVAL_5148 & _EVAL_2424;
  assign _EVAL_3926 = _EVAL_2986 & _EVAL_4751;
  assign _EVAL_4715 = ~_EVAL_5300;
  assign _EVAL_963 = _EVAL_3624 & _EVAL_5543;
  assign _EVAL_5988 = _EVAL_5074 & _EVAL_3509;
  assign _EVAL_1794 = _EVAL_3983 & _EVAL_4536;
  assign _EVAL_5482 = _EVAL_4141 & _EVAL_2748;
  assign _EVAL_1022 = _EVAL_2241 & _EVAL_2748;
  assign _EVAL_1063 = _EVAL_5561 & _EVAL_5308;
  assign _EVAL_4163 = ~_EVAL_5309;
  assign _EVAL_6084 = _EVAL_3820 != 7'h0;
  assign _EVAL_1947 = _EVAL_799 & _EVAL_3702;
  assign _EVAL_1870 = _EVAL_5155 & _EVAL_5543;
  assign _EVAL_1992 = _EVAL_2252 & _EVAL_847;
  assign _EVAL_4431 = _EVAL_5162 & _EVAL_2969;
  assign _EVAL_5845 = _EVAL_4093 & _EVAL_3261;
  assign _EVAL_4834 = _EVAL_3216 & _EVAL_882;
  assign _EVAL_1385 = _EVAL_4322 & _EVAL_5543;
  assign _EVAL_3528 = _EVAL_1145[653];
  assign _EVAL_2572 = _EVAL_774 & _EVAL_2748;
  assign _EVAL_4988 = _EVAL_4795 & _EVAL_2969;
  assign _EVAL_5365 = _EVAL_1536 & _EVAL_3702;
  assign _EVAL_1547 = _EVAL_1147 & _EVAL_4877;
  assign _EVAL_2200 = _EVAL_3188 & _EVAL_1290;
  assign _EVAL_3121 = _EVAL_4627 & _EVAL_5205;
  assign _EVAL_5338 = _EVAL_4187 & _EVAL_4788;
  assign _EVAL_2456 = _EVAL_1145[648];
  assign _EVAL_1884 = _EVAL_5478 & _EVAL_4477;
  assign _EVAL_2991 = _EVAL_1145[655];
  assign _EVAL_2252 = _EVAL_3565 & _EVAL_673;
  assign _EVAL_1980 = _EVAL_4627 & _EVAL_2975;
  assign _EVAL_4444 = _EVAL_2252 & _EVAL_3261;
  assign _EVAL_3608 = _EVAL_4007 & _EVAL_3519;
  assign _EVAL_2420 = _EVAL_5893 & _EVAL_3702;
  assign _EVAL_1974 = _EVAL_1146 & _EVAL_882;
  assign _EVAL_5599 = _EVAL_5074 & _EVAL_5205;
  assign _EVAL_3886 = _EVAL_2842 & _EVAL_3284;
  assign _EVAL_2078 = _EVAL_1145[526];
  assign _EVAL_5678 = _EVAL_778 & _EVAL_3766;
  assign _EVAL_4710 = _EVAL_2782 & _EVAL_2356;
  assign _EVAL_3041 = _EVAL_5816 & _EVAL_2320;
  assign _EVAL_513 = _EVAL_1655 & _EVAL_882;
  assign _EVAL_225 = _EVAL_1945 & _EVAL_5753;
  assign _EVAL_5956 = _EVAL_4627 & _EVAL_4114;
  assign _EVAL_5233 = _EVAL_688 & _EVAL_4477;
  assign _EVAL_1513 = _EVAL_3704 & _EVAL_5464;
  assign _EVAL_3755 = _EVAL_2972 & _EVAL_5289;
  assign _EVAL_2251 = _EVAL_2387 & _EVAL_3379;
  assign _EVAL_564 = _EVAL_5100 & _EVAL_3170;
  assign _EVAL_2144 = _EVAL_5788 & _EVAL_5464;
  assign _EVAL_2900 = _EVAL_1620 & _EVAL_4108;
  assign _EVAL_1364 = _EVAL_1966 & _EVAL_3379;
  assign _EVAL_5840 = _EVAL_3632 & _EVAL_4751;
  assign _EVAL_4218 = _EVAL_2972 & _EVAL_4775;
  assign _EVAL_2734 = _EVAL_5542 & _EVAL_3508;
  assign _EVAL_1975 = _EVAL_1649 & _EVAL_369;
  assign _EVAL_3377 = _EVAL_6032 & _EVAL_5543;
  assign _EVAL_3727 = _EVAL_4093 & _EVAL_4477;
  assign _EVAL_2388 = _EVAL_3574 & _EVAL_2320;
  assign _EVAL_2425 = _EVAL_1145[656];
  assign _EVAL_701 = _EVAL_1242 & _EVAL_847;
  assign _EVAL_1490 = _EVAL_4627 & _EVAL_3038;
  assign _EVAL_827 = _EVAL_1235 & _EVAL_1107;
  assign _EVAL_5471 = _EVAL_3052 & _EVAL_4477;
  assign _EVAL_725 = _EVAL_5642 & _EVAL_2748;
  assign _EVAL_3964 = _EVAL_1876 & _EVAL_847;
  assign _EVAL_1981 = _EVAL_386 & _EVAL_369;
  assign _EVAL_1810 = _EVAL_4757 & _EVAL_3261;
  assign _EVAL_5651 = _EVAL_1125 & _EVAL_847;
  assign _EVAL_3720 = _EVAL_3993 & _EVAL_3398;
  assign _EVAL_1786 = _EVAL_5054 & _EVAL_3487;
  assign _EVAL_1224 = _EVAL_5077 & _EVAL_3418;
  assign _EVAL_3082 = _EVAL_781 & _EVAL_3379;
  assign _EVAL_5404 = _EVAL_5148 & _EVAL_2748;
  assign _EVAL_3455 = _EVAL_5528 & _EVAL_3766;
  assign _EVAL_214 = _EVAL_537 & _EVAL_4160;
  assign _EVAL_4468 = _EVAL_1500 & _EVAL_3261;
  assign _EVAL_5625 = _EVAL_1145[254];
  assign _EVAL_3185 = _EVAL_4137 & _EVAL_3487;
  assign _EVAL_3448 = _EVAL_4795 & _EVAL_2424;
  assign _EVAL_3269 = _EVAL_4888 & _EVAL_5543;
  assign _EVAL_1081 = _EVAL_1625 & _EVAL_2748;
  assign _EVAL_5979 = _EVAL_5074 & _EVAL_4512;
  assign _EVAL_6088 = _EVAL_1316[31:1];
  assign _EVAL_4576 = _EVAL_5148 & _EVAL_1488;
  assign _EVAL_2006 = _EVAL_4314 & _EVAL_2620;
  assign _EVAL_2506 = _EVAL_2631 & _EVAL_3398;
  assign _EVAL_1404 = _EVAL_1677 & _EVAL_882;
  assign _EVAL_5087 = _EVAL_5561 & _EVAL_3647;
  assign _EVAL_5607 = _EVAL_5193 & _EVAL_369;
  assign _EVAL_871 = _EVAL_828 & _EVAL_2382;
  assign _EVAL_1729 = _EVAL_5561 & _EVAL_5829;
  assign _EVAL_3602 = _EVAL_828 & _EVAL_5464;
  assign _EVAL_3699 = _EVAL_1625 & _EVAL_2424;
  assign _EVAL_5588 = _EVAL_2972 & _EVAL_3766;
  assign _EVAL_1747 = _EVAL_4627 & _EVAL_2082;
  assign _EVAL_4664 = _EVAL_3236 != 4'h0;
  assign _EVAL_5132 = _EVAL_3295 & _EVAL_673;
  assign _EVAL_4073 = _EVAL_4187 & _EVAL_4160;
  assign _EVAL_1165 = _EVAL_688 & _EVAL_3398;
  assign _EVAL_1082 = _EVAL_787 & _EVAL_3379;
  assign _EVAL_376 = _EVAL_2241 & _EVAL_3702;
  assign _EVAL_619 = _EVAL_5766 & _EVAL_3766;
  assign _EVAL_2145 = _EVAL_5561 & _EVAL_5136;
  assign _EVAL_1850 = _EVAL_3815 & _EVAL_1735;
  assign _EVAL_3202 = _EVAL_3121 & _EVAL_3379;
  assign _EVAL_4379 = _EVAL_617 & _EVAL_3702;
  assign _EVAL_2726 = _EVAL_5068[513];
  assign _EVAL_1155 = _EVAL_5068[523];
  assign _EVAL_5517 = _EVAL_534 & _EVAL_5464;
  assign _EVAL_1745 = _EVAL_5351 & _EVAL_3379;
  assign _EVAL_5990 = _EVAL_668 & _EVAL_2969;
  assign _EVAL_2904 = _EVAL_4620 & _EVAL_2916;
  assign _EVAL_4767 = _EVAL_1920 & _EVAL_847;
  assign _EVAL_5141 = _EVAL_6080 & _EVAL_5850;
  assign _EVAL_2184 = _EVAL_5869 & _EVAL_4477;
  assign _EVAL_5239 = _EVAL_4419 & _EVAL_3261;
  assign _EVAL_3582 = _EVAL_5078 & _EVAL_4104;
  assign _EVAL_4241 = _EVAL_4916 & _EVAL_2382;
  assign _EVAL_5074 = _EVAL_933 & _EVAL_652;
  assign _EVAL_2892 = _EVAL_3264 == 22'h2cc0;
  assign _EVAL_5040 = _EVAL_3689 & _EVAL_2424;
  assign _EVAL_4661 = _EVAL_4393 & _EVAL_673;
  assign _EVAL_3687 = _EVAL_594 & _EVAL_5289;
  assign _EVAL_5015 = _EVAL_5068[528];
  assign _EVAL_4035 = _EVAL_3107 & _EVAL_1488;
  assign _EVAL_4461 = _EVAL_1876 & _EVAL_3487;
  assign _EVAL_3954 = _EVAL_6007 & _EVAL_3261;
  assign _EVAL_5216 = _EVAL_3225 & _EVAL_1226;
  assign _EVAL_4918 = _EVAL_4106 & _EVAL_1290;
  assign _EVAL_5610 = _EVAL_3898 & _EVAL_3702;
  assign _EVAL_1858 = _EVAL_534 & _EVAL_3170;
  assign _EVAL_3688 = _EVAL_2986 & _EVAL_4109;
  assign _EVAL_1832 = _EVAL_4499 & _EVAL_4751;
  assign _EVAL_2567 = _EVAL_3787 & _EVAL_5289;
  assign _EVAL_3033 = _EVAL_2292 & _EVAL_2382;
  assign _EVAL_1349 = _EVAL_5542 & _EVAL_3998;
  assign _EVAL_5079 = _EVAL_4322 & _EVAL_3702;
  assign _EVAL_1739 = _EVAL_2247 & _EVAL_476;
  assign _EVAL_3484 = _EVAL_1622 & _EVAL_3766;
  assign _EVAL_1807 = _EVAL_4219 & _EVAL_2424;
  assign _EVAL_4371 = _EVAL_620 & _EVAL_4109;
  assign _EVAL_566 = _EVAL_3322 & _EVAL_1198;
  assign _EVAL_5430 = _EVAL_5561 & _EVAL_1695;
  assign _EVAL_1601 = _EVAL_6022 & _EVAL_5543;
  assign _EVAL_1518 = _EVAL_6051 & _EVAL_5850;
  assign _EVAL_4900 = _EVAL_5561 & _EVAL_5269;
  assign _EVAL_3322 = _EVAL_590 & _EVAL_3379;
  assign _EVAL_3859 = _EVAL_375 & _EVAL_3379;
  assign _EVAL_2040 = _EVAL_5811 & _EVAL_3702;
  assign _EVAL_5276 = _EVAL_735 & _EVAL_4751;
  assign _EVAL_2002 = _EVAL_5074 & _EVAL_5625;
  assign _EVAL_5948 = _EVAL_2902 & _EVAL_2748;
  assign _EVAL_3626 = _EVAL_6032 & _EVAL_3702;
  assign _EVAL_1272 = _EVAL_528 & _EVAL_2382;
  assign _EVAL_1195 = _EVAL_857 & _EVAL_2748;
  assign _EVAL_2498 = _EVAL_3609 & _EVAL_552;
  assign _EVAL_2868 = _EVAL_792 & _EVAL_673;
  assign _EVAL_2192 = _EVAL_5243 & _EVAL_3379;
  assign _EVAL_3551 = _EVAL_4783 & _EVAL_1488;
  assign _EVAL_4987 = _EVAL_1667 & _EVAL_3379;
  assign _EVAL_3177 = _EVAL_402 & _EVAL_1198;
  assign _EVAL_3706 = _EVAL_1051 & _EVAL_3379;
  assign _EVAL_303 = _EVAL_4200 & _EVAL_882;
  assign _EVAL_1588 = _EVAL_2876 & _EVAL_2258;
  assign _EVAL_3984 = _EVAL_5450 & _EVAL_1735;
  assign _EVAL_646 = _EVAL_1039 & _EVAL_4477;
  assign _EVAL_4616 = _EVAL_4488 & _EVAL_3398;
  assign _EVAL_3663 = ~_EVAL_487;
  assign _EVAL_2555 = ~_EVAL_4119;
  assign _EVAL_2891 = _EVAL_5246 & _EVAL_3418;
  assign _EVAL_663 = _EVAL_284 & _EVAL_5543;
  assign _EVAL_1361 = _EVAL_947 & _EVAL_673;
  assign _EVAL_2723 = _EVAL_2005 & _EVAL_369;
  assign _EVAL_3816 = _EVAL_4507 & _EVAL_3284;
  assign _EVAL_5342 = _EVAL_2126 & _EVAL_3379;
  assign _EVAL_987 = _EVAL_1361 & _EVAL_3418;
  assign _EVAL_2599 = _EVAL_1370 & _EVAL_3154;
  assign _EVAL_5066 = _EVAL_3524 & _EVAL_369;
  assign _EVAL_5155 = _EVAL_793 & _EVAL_3379;
  assign _EVAL_1090 = _EVAL_5561 & _EVAL_2520;
  assign _EVAL_5271 = _EVAL_5795 & _EVAL_1009;
  assign _EVAL_5589 = _EVAL_5890 & _EVAL_318;
  assign _EVAL_5420 = _EVAL_5561 & _EVAL_2176;
  assign _EVAL_1603 = _EVAL_2753[8];
  assign _EVAL_578 = _EVAL_2170 & _EVAL_2748;
  assign _EVAL_6024 = _EVAL_5074 & _EVAL_5593;
  assign _EVAL_3049 = _EVAL_4499 & _EVAL_1735;
  assign TLMonitor__EVAL = _EVAL_88;
  assign _EVAL_410 = ~_EVAL_5878;
  assign _EVAL_3784 = _EVAL_6087 & _EVAL_2424;
  assign _EVAL_1782 = _EVAL_769 & _EVAL_3487;
  assign _EVAL_539 = ~_EVAL_5345;
  assign _EVAL_5888 = _EVAL_1920 & _EVAL_3487;
  assign _EVAL_352 = _EVAL_589 & _EVAL_1735;
  assign _EVAL_222 = _EVAL_5074 & _EVAL_731;
  assign _EVAL_2019 = _EVAL_5561 & _EVAL_5015;
  assign _EVAL_2260 = _EVAL_2859 & _EVAL_673;
  assign _EVAL_5114 = _EVAL_4689 & _EVAL_1735;
  assign _EVAL_1957 = _EVAL_5074 & _EVAL_3807;
  assign _EVAL_4647 = _EVAL_1622 & _EVAL_1009;
  assign _EVAL_4265 = _EVAL_2868 & _EVAL_3154;
  assign _EVAL_1911 = _EVAL_1620 & _EVAL_4751;
  assign _EVAL_4109 = _EVAL_1470 != 4'h0;
  assign _EVAL_2899 = _EVAL_5353 & _EVAL_3702;
  assign _EVAL_5217 = _EVAL_5068[545];
  assign _EVAL_5507 = _EVAL_3216 & _EVAL_847;
  assign _EVAL_3820 = _EVAL_1316[15:9];
  assign _EVAL_947 = _EVAL_5561 & _EVAL_786;
  assign _EVAL_3802 = _EVAL_1542 & _EVAL_847;
  assign _EVAL_5541 = _EVAL_5342 & _EVAL_1198;
  assign _EVAL_5123 = _EVAL_584 & _EVAL_801;
  assign _EVAL_4188 = _EVAL_2907 & _EVAL_3702;
  assign _EVAL_1944 = _EVAL_5788 & _EVAL_2382;
  assign _EVAL_206 = _EVAL_1145[589];
  assign _EVAL_1752 = _EVAL_1649 & _EVAL_2748;
  assign _EVAL_3863 = _EVAL_6080 & _EVAL_4108;
  assign _EVAL_3284 = _EVAL_2688 == 4'hf;
  assign _EVAL_698 = _EVAL_1281 & _EVAL_1290;
  assign _EVAL_1545 = _EVAL_2292 & _EVAL_4109;
  assign _EVAL_2405 = _EVAL_1145[539];
  assign _EVAL_4912 = _EVAL_298 & _EVAL_4993;
  assign _EVAL_1736 = _EVAL_5153 & _EVAL_2320;
  assign _EVAL_2041 = _EVAL_2585 & _EVAL_847;
  assign _EVAL_5144 = _EVAL_4627 & _EVAL_4428;
  assign _EVAL_2798 = _EVAL_1316[11:8];
  assign _EVAL_941 = _EVAL_5561 & _EVAL_3977;
  assign _EVAL_3579 = _EVAL_4525 & _EVAL_5464;
  assign _EVAL_3880 = _EVAL_3436 & _EVAL_4160;
  assign _EVAL_1428 = _EVAL_309 & _EVAL_5850;
  assign _EVAL_341 = _EVAL_735 & _EVAL_3170;
  assign _EVAL_2615 = ~_EVAL_1188;
  assign _EVAL_3794 = _EVAL_4627 & _EVAL_2465;
  assign _EVAL_1926 = _EVAL_1649 & _EVAL_2424;
  assign _EVAL_819 = _EVAL_4625 & _EVAL_3702;
  assign _EVAL_5240 = _EVAL_4783 & _EVAL_3702;
  assign _EVAL_2533 = _EVAL_251 & _EVAL_5543;
  assign _EVAL_6096 = _EVAL_5561 & _EVAL_2661;
  assign _EVAL_446 = _EVAL_4502 & _EVAL_3379;
  assign _EVAL_4086 = _EVAL_1145[516];
  assign _EVAL_4061 = _EVAL_2086 & _EVAL_5416;
  assign _EVAL_5570 = _EVAL_4219 & _EVAL_2748;
  assign _EVAL_574 = _EVAL_1145[659];
  assign _EVAL_1046 = _EVAL_4567 & _EVAL_3487;
  assign _EVAL_857 = _EVAL_3794 & _EVAL_3379;
  assign _EVAL_4909 = _EVAL_3490 & _EVAL_2892;
  assign _EVAL_1127 = _EVAL_3783 & _EVAL_3874;
  assign _EVAL_5456 = ~_EVAL_1826;
  assign _EVAL_3948 = _EVAL_4627 & _EVAL_2525;
  assign _EVAL_3830 = _EVAL_5618 & _EVAL_5543;
  assign _EVAL_2538 = _EVAL_5074 & _EVAL_413;
  assign _EVAL_3992 = _EVAL_5530 & _EVAL_3379;
  assign _EVAL_1867 = _EVAL_4618 & _EVAL_1009;
  assign _EVAL_3841 = _EVAL_3052 & _EVAL_3398;
  assign _EVAL_5854 = _EVAL_4145 & _EVAL_3379;
  assign _EVAL_3425 = _EVAL_529 & _EVAL_1198;
  assign _EVAL_2809 = _EVAL_1854 & _EVAL_882;
  assign _EVAL_4521 = _EVAL_3920 & _EVAL_1290;
  assign _EVAL_1262 = _EVAL_212 & _EVAL_1888;
  assign _EVAL_633 = _EVAL_1145[520];
  assign _EVAL_2280 = _EVAL_1312 & _EVAL_1488;
  assign _EVAL_777 = _EVAL_4042 & _EVAL_4993;
  assign _EVAL_3776 = _EVAL_3624 & _EVAL_6084;
  assign _EVAL_2383 = _EVAL_6059 & _EVAL_3487;
  assign _EVAL_2710 = _EVAL_2260 & _EVAL_3398;
  assign _EVAL_856 = ~_EVAL_4184;
  assign _EVAL_937 = _EVAL_2292 & _EVAL_1735;
  assign _EVAL_5055 = _EVAL_5854 & _EVAL_5299;
  assign _EVAL_5478 = _EVAL_3237 & _EVAL_673;
  assign _EVAL_1995 = _EVAL_4044 & _EVAL_4477;
  assign _EVAL_3640 = _EVAL_3188 & _EVAL_4664;
  assign _EVAL_4494 = _EVAL_2454 & _EVAL_4108;
  assign _EVAL_1332 = _EVAL_6087 & _EVAL_2969;
  assign _EVAL_3361 = _EVAL_3689 & _EVAL_2748;
  assign _EVAL_2433 = _EVAL_5561 & _EVAL_5711;
  assign _EVAL_3766 = _EVAL_3427 != 4'h0;
  assign _EVAL_1624 = _EVAL_3787 & _EVAL_3766;
  assign _EVAL_1096 = _EVAL_4144 & _EVAL_2956;
  assign _EVAL_3878 = _EVAL_1920 & _EVAL_3154;
  assign _EVAL_4682 = _EVAL_4144 & _EVAL_5299;
  assign _EVAL_4451 = _EVAL_3837 & _EVAL_2969;
  assign _EVAL_162 = _EVAL_4175 & _EVAL_3154;
  assign _EVAL_1076 = _EVAL_1408 & _EVAL_4854;
  assign _EVAL_3648 = _EVAL_5561 & _EVAL_5637;
  assign _EVAL_4137 = _EVAL_4432 & _EVAL_673;
  assign _EVAL_4280 = _EVAL_475 & _EVAL_5299;
  assign _EVAL_5082 = _EVAL_4841 & _EVAL_847;
  assign _EVAL_3321 = _EVAL_1316[31:25];
  assign _EVAL_4501 = _EVAL_5054 & _EVAL_4477;
  assign _EVAL_4627 = _EVAL_933 & _EVAL_4135;
  assign _EVAL_3973 = _EVAL_1677 & _EVAL_3398;
  assign _EVAL_5440 = _EVAL_5443 & _EVAL_673;
  assign _EVAL_377 = _EVAL_4577 & _EVAL_5753;
  assign _EVAL_469 = _EVAL_3837 & _EVAL_5543;
  assign _EVAL_3414 = _EVAL_4227 & _EVAL_3379;
  assign _EVAL_1716 = _EVAL_3935 & _EVAL_1488;
  assign _EVAL_5509 = _EVAL_2753[12];
  assign _EVAL_4069 = _EVAL_581 & _EVAL_5299;
  assign _EVAL_475 = _EVAL_1557 & _EVAL_3379;
  assign _EVAL_1207 = _EVAL_4462 & _EVAL_587;
  assign _EVAL_2376 = _EVAL_4844 & _EVAL_3379;
  assign _EVAL_5752 = _EVAL_668 & _EVAL_2748;
  assign _EVAL_1402 = _EVAL_5132 & _EVAL_3487;
  assign _EVAL_3288 = _EVAL_538 & _EVAL_5543;
  assign _EVAL_3701 = _EVAL_1145[512];
  assign _EVAL_467 = _EVAL_4187 & _EVAL_1290;
  assign _EVAL_888 = _EVAL_5074 & _EVAL_5656;
  assign _EVAL_6001 = _EVAL_617 & _EVAL_2748;
  assign _EVAL_4189 = _EVAL_6033 & _EVAL_5753;
  assign _EVAL_2274 = _EVAL_451 & _EVAL_801;
  assign _EVAL_2363 = _EVAL_2585 & _EVAL_882;
  assign _EVAL_3976 = _EVAL_486 & _EVAL_3702;
  assign _EVAL_4855 = _EVAL_4219 & _EVAL_6084;
  assign _EVAL_2142 = _EVAL_3837 & _EVAL_1488;
  assign _EVAL_4145 = _EVAL_5074 & _EVAL_5590;
  assign _EVAL_3485 = {_EVAL_2153,_EVAL_5509,_EVAL_2879,_EVAL_1603,_EVAL_5827,_EVAL_3759,_EVAL_1972,_EVAL_3315,_EVAL_1105,_EVAL_5917};
  assign _EVAL_3728 = _EVAL_4581 & _EVAL_2956;
  assign _EVAL_3996 = _EVAL_1439 & _EVAL_673;
  assign _EVAL_2810 = _EVAL_589 & _EVAL_4108;
  assign _EVAL_4423 = _EVAL_4661 & _EVAL_5753;
  assign _EVAL_1231 = _EVAL_2631 & _EVAL_847;
  assign _EVAL_1585 = ~_EVAL_1831;
  assign _EVAL_5640 = _EVAL_4222 & _EVAL_3418;
  assign _EVAL_398 = _EVAL_1145[662];
  assign _EVAL_2796 = _EVAL_3152 & _EVAL_1443;
  assign _EVAL_4586 = _EVAL_3364 & _EVAL_847;
  assign _EVAL_4527 = _EVAL_2205 & _EVAL_2382;
  assign _EVAL_692 = _EVAL_3632 & _EVAL_2382;
  assign _EVAL_1095 = _EVAL_2260 & _EVAL_847;
  assign _EVAL_3647 = _EVAL_5068[524];
  assign _EVAL_321 = ~_EVAL_3940;
  assign _EVAL_271 = _EVAL_4821 & _EVAL_2748;
  assign _EVAL_3512 = _EVAL_1747 & _EVAL_3379;
  assign _EVAL_1856 = _EVAL_5132 & _EVAL_3154;
  assign _EVAL_5564 = _EVAL_2592 & _EVAL_2424;
  assign _EVAL_4498 = _EVAL_1057 & _EVAL_1340;
  assign _EVAL_4890 = _EVAL_3787 & _EVAL_1290;
  assign _EVAL_5259 = _EVAL_3961 & _EVAL_2424;
  assign TLMonitor__EVAL_10 = Queue__EVAL_9;
  assign _EVAL_4333 = _EVAL_4175 & _EVAL_847;
  assign _EVAL_1965 = _EVAL_5994 & _EVAL_3487;
  assign _EVAL_4861 = _EVAL_3574 & _EVAL_4109;
  assign _EVAL_3375 = _EVAL_5440 & _EVAL_3418;
  assign _EVAL_5797 = _EVAL_3055 == 4'hf;
  assign _EVAL_5075 = ~_EVAL_4443;
  assign _EVAL_3224 = _EVAL_3706 & _EVAL_6084;
  assign _EVAL_2773 = _EVAL_1971 & _EVAL_1488;
  assign _EVAL_5196 = _EVAL_3826 & _EVAL_2956;
  assign _EVAL_5053 = _EVAL_1677 & _EVAL_4477;
  assign _EVAL_5310 = _EVAL_1312 & _EVAL_5543;
  assign _EVAL_5059 = _EVAL_1446 & _EVAL_369;
  assign _EVAL_5304 = ~_EVAL_2291;
  assign _EVAL_5856 = _EVAL_5561 & _EVAL_3694;
  assign _EVAL_996 = _EVAL_1689 & _EVAL_1488;
  assign _EVAL_1244 = _EVAL_4499 & _EVAL_5464;
  assign _EVAL_5356 = _EVAL_4137 & _EVAL_4477;
  assign _EVAL_3074 = _EVAL_3082 & _EVAL_1488;
  assign _EVAL_828 = _EVAL_4782 & _EVAL_3379;
  assign _EVAL_976 = _EVAL_4372 & _EVAL_2748;
  assign _EVAL_3301 = _EVAL_573 & _EVAL_3379;
  assign _EVAL_1212 = _EVAL_2725 & _EVAL_3261;
  assign _EVAL_4312 = _EVAL_3436 & _EVAL_801;
  assign _EVAL_774 = _EVAL_1590 & _EVAL_3379;
  assign _EVAL_1488 = _EVAL_709 != 7'h0;
  assign _EVAL_1097 = _EVAL_6087 & _EVAL_2748;
  assign _EVAL_390 = _EVAL_5561 & _EVAL_1093;
  assign _EVAL_1673 = _EVAL_1945 & _EVAL_4775;
  assign _EVAL_5954 = _EVAL_3704 & _EVAL_3170;
  assign _EVAL_2658 = _EVAL_5930 & _EVAL_1488;
  assign _EVAL_2657 = _EVAL_5561 & _EVAL_3200;
  assign _EVAL_6077 = _EVAL_5561 & _EVAL_2515;
  assign _EVAL_3302 = _EVAL_3107 & _EVAL_2424;
  assign _EVAL_5465 = _EVAL_4596 & _EVAL_4775;
  assign _EVAL_983 = _EVAL_617 & _EVAL_369;
  assign _EVAL_4971 = _EVAL_2260 & _EVAL_3261;
  assign _EVAL_2414 = _EVAL_1202 & _EVAL_4477;
  assign _EVAL_5982 = _EVAL_3156 & _EVAL_5543;
  assign _EVAL_3809 = _EVAL_2251 & _EVAL_5543;
  assign _EVAL_5313 = _EVAL_5561 & _EVAL_2052;
  assign _EVAL_4158 = _EVAL_5163 & _EVAL_4209;
  assign _EVAL_4094 = _EVAL_581 & _EVAL_3284;
  assign _EVAL_4920 = _EVAL_2170 & _EVAL_2424;
  assign _EVAL_936 = _EVAL_1145[645];
  assign _EVAL_1346 = _EVAL_4550 & _EVAL_3702;
  assign _EVAL_1962 = _EVAL_910 & _EVAL_3379;
  assign _EVAL_3511 = _EVAL_362 & _EVAL_1009;
  assign _EVAL_5455 = _EVAL_831 & _EVAL_2748;
  assign _EVAL_1897 = _EVAL_284 & _EVAL_2424;
  assign _EVAL_3476 = _EVAL_2593 & _EVAL_3379;
  assign _EVAL_3437 = _EVAL_5074 & _EVAL_4601;
  assign _EVAL_2262 = _EVAL_3993 & _EVAL_4477;
  assign _EVAL_562 = _EVAL_3032 & _EVAL_1009;
  assign _EVAL_5020 = _EVAL_1419 & _EVAL_2748;
  assign _EVAL_2037 = _EVAL_4028 & _EVAL_3379;
  assign _EVAL_1881 = _EVAL_2646 & _EVAL_5445;
  assign _EVAL_2204 = _EVAL_5819 & _EVAL_1009;
  assign _EVAL_1541 = _EVAL_1945 & _EVAL_3766;
  assign _EVAL_2712 = _EVAL_3574 & _EVAL_4751;
  assign _EVAL_2174 = _EVAL_5068[540];
  assign _EVAL_5587 = _EVAL_1067 & _EVAL_1290;
  assign _EVAL_1045 = _EVAL_4612 & _EVAL_2565;
  assign _EVAL_1107 = ~_EVAL_5696;
  assign _EVAL_5529 = _EVAL_4525 & _EVAL_4108;
  assign _EVAL_2548 = _EVAL_6022 & _EVAL_2969;
  assign _EVAL_2005 = _EVAL_2426 & _EVAL_3379;
  assign _EVAL_1199 = _EVAL_4627 & _EVAL_2456;
  assign _EVAL_1458 = _EVAL_4795 & _EVAL_2748;
  assign _EVAL_476 = ~_EVAL_3286;
  assign _EVAL_2179 = _EVAL_4627 & _EVAL_4512;
  assign _EVAL_2973 = _EVAL_2339 & _EVAL_856;
  assign _EVAL_5483 = _EVAL_1865 & _EVAL_3261;
  assign _EVAL_814 = _EVAL_4604 & _EVAL_3766;
  assign _EVAL_2066 = _EVAL_5598 & _EVAL_3398;
  assign _EVAL_4598 = _EVAL_6059 & _EVAL_3398;
  assign _EVAL_4326 = _EVAL_4083 & _EVAL_4477;
  assign _EVAL_4581 = _EVAL_4910 & _EVAL_3379;
  assign _EVAL_3010 = _EVAL_4093 & _EVAL_3487;
  assign _EVAL_2068 = _EVAL_5068[531];
  assign _EVAL_5900 = _EVAL_5353 & _EVAL_1488;
  assign _EVAL_1439 = _EVAL_5561 & _EVAL_3502;
  assign _EVAL_5302 = _EVAL_5662 & _EVAL_3398;
  assign _EVAL_4475 = _EVAL_3652 & _EVAL_2438;
  assign _EVAL_6036 = _EVAL_961 & _EVAL_3702;
  assign _EVAL_307 = _EVAL_3787 & _EVAL_4775;
  assign _EVAL_3888 = _EVAL_4916 & _EVAL_4109;
  assign _EVAL_3071 = _EVAL_1067 & _EVAL_4664;
  assign _EVAL_3505 = _EVAL_4235 & _EVAL_369;
  assign _EVAL_3412 = _EVAL_3055 != 4'h0;
  assign _EVAL_5549 = _EVAL_2255 & _EVAL_3379;
  assign _EVAL_5598 = _EVAL_2367 & _EVAL_673;
  assign _EVAL_933 = _EVAL_112 & _EVAL_2329;
  assign _EVAL_4623 = _EVAL_2304 & _EVAL_3379;
  assign _EVAL_5837 = _EVAL_1145[664];
  assign _EVAL_910 = _EVAL_5074 & _EVAL_4605;
  assign _EVAL_4392 = _EVAL_2205 & _EVAL_4108;
  assign _EVAL_591 = _EVAL_1040 & _EVAL_954;
  assign _EVAL_5352 = _EVAL_5795 & _EVAL_4775;
  assign _EVAL_2953 = _EVAL_5293 & _EVAL_1489;
  assign _EVAL_5500 = _EVAL_4525 & _EVAL_4751;
  assign _EVAL_6007 = _EVAL_249 & _EVAL_673;
  assign _EVAL_3237 = _EVAL_5561 & _EVAL_2068;
  assign _EVAL_1774 = _EVAL_774 & _EVAL_369;
  assign _EVAL_6059 = _EVAL_5420 & _EVAL_673;
  assign _EVAL_3369 = _EVAL_3052 & _EVAL_3487;
  assign _EVAL_4289 = _EVAL_5100 & _EVAL_5464;
  assign _EVAL_3630 = _EVAL_2873 & _EVAL_3284;
  assign _EVAL_2340 = _EVAL_5561 & _EVAL_923;
  assign _EVAL_5135 = _EVAL_3632 & _EVAL_5464;
  assign _EVAL_5647 = _EVAL_2725 & _EVAL_3418;
  assign _EVAL_6099 = _EVAL_3156 & _EVAL_3702;
  assign _EVAL_1553 = _EVAL_1008 & _EVAL_673;
  assign _EVAL_803 = _EVAL_2338 & _EVAL_369;
  assign _EVAL_5869 = _EVAL_2665 & _EVAL_673;
  assign _EVAL_4432 = _EVAL_5561 & _EVAL_1300;
  assign _EVAL_621 = _EVAL_5063 & _EVAL_3154;
  assign _EVAL_1631 = ~_EVAL_5558;
  assign _EVAL_5130 = _EVAL_2793 & _EVAL_3398;
  assign _EVAL_2736 = _EVAL_386 & _EVAL_2424;
  assign _EVAL_877 = _EVAL_5206 & _EVAL_1198;
  assign _EVAL_1246 = _EVAL_620 & _EVAL_5850;
  assign _EVAL_2999 = ~_EVAL_643;
  assign _EVAL_1783 = _EVAL_6075 & _EVAL_3261;
  assign _EVAL_5897 = _EVAL_3859 & _EVAL_5299;
  assign _EVAL_1792 = _EVAL_5662 & _EVAL_4477;
  assign _EVAL_2361 = _EVAL_2205 & _EVAL_5850;
  assign _EVAL_3008 = _EVAL_4083 & _EVAL_882;
  assign _EVAL_3409 = _EVAL_4841 & _EVAL_4477;
  assign _EVAL_5643 = _EVAL_4755 & _EVAL_4108;
  assign _EVAL_3598 = _EVAL_4175 & _EVAL_3487;
  assign _EVAL_927 = ~_EVAL_4810;
  assign _EVAL_3220 = _EVAL_1941 & _EVAL_3379;
  assign _EVAL_4202 = _EVAL_2733 & _EVAL_673;
  assign _EVAL_3300 = _EVAL_3226 & _EVAL_5464;
  assign _EVAL_1548 = _EVAL_4149 & _EVAL_2748;
  assign _EVAL_3347 = _EVAL_5561 & _EVAL_5169;
  assign _EVAL_1162 = _EVAL_3996 & _EVAL_5289;
  assign _EVAL_3179 = _EVAL_1125 & _EVAL_3418;
  assign _EVAL_4926 = _EVAL_897 & _EVAL_5299;
  assign TLMonitor__EVAL_2 = _EVAL_106;
  assign _EVAL_5380 = _EVAL_4627 & _EVAL_2117;
  assign _EVAL_565 = _EVAL_935 & _EVAL_2748;
  assign _EVAL_2430 = _EVAL_1364 & _EVAL_1198;
  assign _EVAL_3749 = _EVAL_5598 & _EVAL_882;
  assign _EVAL_5051 = _EVAL_302 & _EVAL_5543;
  assign _EVAL_3894 = _EVAL_1960 & _EVAL_587;
  assign _EVAL_5659 = _EVAL_3414 & _EVAL_2969;
  assign _EVAL_928 = _EVAL_2998 & _EVAL_882;
  assign _EVAL_1996 = _EVAL_4627 & _EVAL_6008;
  assign _EVAL_4628 = _EVAL_3451 & _EVAL_3261;
  assign _EVAL_1627 = _EVAL_5561 & _EVAL_6055;
  assign _EVAL_3817 = _EVAL_2241 & _EVAL_5543;
  assign _EVAL_587 = _EVAL_5905 != 4'h0;
  assign _EVAL_4052 = _EVAL_589 & _EVAL_5850;
  assign _EVAL_961 = _EVAL_3523 & _EVAL_3379;
  assign _EVAL_5662 = _EVAL_4727 & _EVAL_673;
  assign _EVAL_1915 = _EVAL_479 & _EVAL_1488;
  assign _EVAL_3488 = _EVAL_402 & _EVAL_2956;
  assign _EVAL_4253 = _EVAL_2312 & _EVAL_4715;
  assign _EVAL_5492 = _EVAL_4627 & _EVAL_5733;
  assign _EVAL_2129 = _EVAL_2877 & _EVAL_369;
  assign _EVAL_1489 = ~_EVAL_4348;
  assign _EVAL_3801 = _EVAL_4627 & _EVAL_2983;
  assign _EVAL_4200 = _EVAL_4668 & _EVAL_673;
  assign _EVAL_1854 = _EVAL_1696 & _EVAL_673;
  assign _EVAL_3514 = _EVAL_4462 & _EVAL_4775;
  assign _EVAL_3231 = _EVAL_1677 & _EVAL_3261;
  assign _EVAL_2969 = _EVAL_1989 != 7'h0;
  assign _EVAL_5590 = _EVAL_1145[652];
  assign _EVAL_4118 = _EVAL_4627 & _EVAL_622;
  assign _EVAL_4830 = _EVAL_5074 & _EVAL_3923;
  assign _EVAL_1170 = _EVAL_2725 & _EVAL_847;
  assign _EVAL_492 = _EVAL_4627 & _EVAL_1604;
  assign _EVAL_1707 = _EVAL_4627 & _EVAL_3210;
  assign _EVAL_4319 = _EVAL_4083 & _EVAL_3487;
  assign _EVAL_2023 = _EVAL_4462 & _EVAL_3766;
  assign _EVAL_5200 = _EVAL_4137 & _EVAL_847;
  assign _EVAL_1343 = _EVAL_5074 & _EVAL_2456;
  assign _EVAL_4205 = _EVAL_1536 & _EVAL_1488;
  assign _EVAL_4314 = _EVAL_768 & _EVAL_3379;
  assign _EVAL_4492 = ~_EVAL_1041;
  assign _EVAL_3616 = _EVAL_1145[528];
  assign _EVAL_2830 = _EVAL_1202 & _EVAL_3261;
  assign _EVAL_4904 = _EVAL_5561 & _EVAL_5491;
  assign _EVAL_2585 = _EVAL_1727 & _EVAL_673;
  assign _EVAL_2992 = _EVAL_3107 & _EVAL_2969;
  assign _EVAL_3704 = _EVAL_2043 & _EVAL_3379;
  assign _EVAL_5353 = _EVAL_4667 & _EVAL_3379;
  assign _EVAL_1019 = _EVAL_4755 & _EVAL_2382;
  assign _EVAL_183 = _EVAL_5561 & _EVAL_854;
  assign _EVAL_3195 = _EVAL_5940 & _EVAL_354;
  assign _EVAL_3593 = _EVAL_3826 & _EVAL_3284;
  assign _EVAL_1084 = _EVAL_5618 & _EVAL_6084;
  assign _EVAL_2375 = _EVAL_4083 & _EVAL_3418;
  assign _EVAL_2060 = _EVAL_3197 & _EVAL_3471;
  assign _EVAL_3063 = _EVAL_1865 & _EVAL_847;
  assign _EVAL_2356 = ~_EVAL_666;
  assign _EVAL_1044 = _EVAL_4200 & _EVAL_3154;
  assign _EVAL_699 = _EVAL_1145[672];
  assign _EVAL_3660 = _EVAL_3815 & _EVAL_4751;
  assign _EVAL_4210 = _EVAL_4625 & _EVAL_5543;
  assign _EVAL_2008 = _EVAL_1145[658];
  assign _EVAL_1933 = _EVAL_528 & _EVAL_5464;
  assign _EVAL_5616 = _EVAL_5074 & _EVAL_2525;
  assign _EVAL_1480 = _EVAL_3845 & _EVAL_5299;
  assign _EVAL_2402 = _EVAL_3032 & _EVAL_4775;
  assign _EVAL_946 = _EVAL_4254 & _EVAL_587;
  assign _EVAL_5474 = _EVAL_1103 & _EVAL_3702;
  assign _EVAL_409 = _EVAL_5063 & _EVAL_3418;
  assign _EVAL_3811 = _EVAL_3992 & _EVAL_5445;
  assign _EVAL_2965 = _EVAL_5193 & _EVAL_5543;
  assign _EVAL_570 = _EVAL_3512 & _EVAL_6084;
  assign _EVAL_1500 = _EVAL_5724 & _EVAL_673;
  assign _EVAL_1069 = _EVAL_1145[647];
  assign _EVAL_3565 = _EVAL_5561 & _EVAL_5241;
  assign _EVAL_6002 = _EVAL_1158 & _EVAL_847;
  assign _EVAL_449 = _EVAL_5561 & _EVAL_5050;
  assign _EVAL_4964 = _EVAL_4192 & _EVAL_369;
  assign _EVAL_1122 = _EVAL_4974 & _EVAL_4108;
  assign _EVAL_309 = _EVAL_641 & _EVAL_3379;
  assign _EVAL_2698 = _EVAL_3226 & _EVAL_3170;
  assign _EVAL_244 = _EVAL_1920 & _EVAL_3398;
  assign _EVAL_3394 = _EVAL_3130 & _EVAL_2748;
  assign _EVAL_4227 = _EVAL_4627 & _EVAL_3684;
  assign _EVAL_5676 = _EVAL_4736 & _EVAL_673;
  assign _EVAL_2500 = _EVAL_905 & _EVAL_4477;
  assign _EVAL_5344 = _EVAL_4936 & _EVAL_3379;
  assign _EVAL_1201 = _EVAL_4219 & _EVAL_369;
  assign _EVAL_3239 = _EVAL_2192 & _EVAL_1488;
  assign _EVAL_2656 = _EVAL_5618 & _EVAL_3702;
  assign _EVAL_5280 = _EVAL_4044 & _EVAL_3154;
  assign _EVAL_2540 = _EVAL_407 & _EVAL_2969;
  assign _EVAL_4485 = _EVAL_1865 & _EVAL_3487;
  assign _EVAL_3246 = _EVAL_2877 & _EVAL_5543;
  assign _EVAL_4589 = _EVAL_1620 & _EVAL_4109;
  assign _EVAL_1509 = _EVAL_5450 & _EVAL_5850;
  assign _EVAL_1530 = _EVAL_4419 & _EVAL_3418;
  assign _EVAL_429 = _EVAL_2631 & _EVAL_3487;
  assign _EVAL_3089 = _EVAL_4627 & _EVAL_699;
  assign _EVAL_3117 = _EVAL_4336 & _EVAL_4504;
  assign _EVAL_5778 = _EVAL_5528 & _EVAL_4775;
  assign _EVAL_3875 = _EVAL_2675 & _EVAL_6084;
  assign _EVAL_2395 = _EVAL_2717 & _EVAL_541;
  assign _EVAL_5223 = _EVAL_5561 & _EVAL_6004;
  assign _EVAL_335 = _EVAL_4627 & _EVAL_2078;
  assign _EVAL_360 = _EVAL_2842 & _EVAL_2956;
  assign _EVAL_4552 = _EVAL_1468 ? 8'hff : 8'h0;
  assign _EVAL_3175 = _EVAL_679 & _EVAL_369;
  assign _EVAL_4688 = _EVAL_5344 & _EVAL_4109;
  assign _EVAL_4039 = _EVAL_3183 & _EVAL_3702;
  assign _EVAL_205 = _EVAL_943 & _EVAL_2888;
  assign _EVAL_1183 = _EVAL_5440 & _EVAL_3154;
  assign _EVAL_407 = _EVAL_5602 & _EVAL_3379;
  assign _EVAL_3192 = _EVAL_446 & _EVAL_1198;
  assign _EVAL_2468 = _EVAL_891 & _EVAL_5424;
  assign _EVAL_3881 = _EVAL_2907 & _EVAL_369;
  assign _EVAL_2680 = _EVAL_5074 & _EVAL_4656;
  assign _EVAL_4522 = ~_EVAL_5600;
  assign _EVAL_2885 = _EVAL_3346 & _EVAL_4477;
  assign _EVAL_2329 = Queue__EVAL_9;
  assign _EVAL_2571 = _EVAL_2793 & _EVAL_3487;
  assign _EVAL_2333 = _EVAL_2484 & _EVAL_478;
  assign _EVAL_820 = _EVAL_3996 & _EVAL_3766;
  assign _EVAL_1717 = _EVAL_1633 & _EVAL_1488;
  assign _EVAL_1611 = _EVAL_3107 & _EVAL_3702;
  assign _EVAL_4587 = _EVAL_3216 & _EVAL_3487;
  assign _EVAL_3206 = _EVAL_5344 & _EVAL_4751;
  assign _EVAL_2243 = _EVAL_1962 & _EVAL_1198;
  assign _EVAL_3209 = _EVAL_1145[667];
  assign _EVAL_3329 = _EVAL_1145[257];
  assign _EVAL_3006 = _EVAL_5561 & _EVAL_5267;
  assign _EVAL_5679 = _EVAL_6007 & _EVAL_3398;
  assign _EVAL_4851 = _EVAL_4627 & _EVAL_6076;
  assign _EVAL_4302 = _EVAL_1493 & _EVAL_800;
  assign _EVAL_3258 = _EVAL_2550 & _EVAL_5753;
  assign _EVAL_2613 = _EVAL_4149 & _EVAL_5543;
  assign _EVAL_2246 = _EVAL_1344 & _EVAL_4477;
  assign _EVAL_2107 = _EVAL_4661 & _EVAL_1290;
  assign _EVAL_5264 = _EVAL_2607 & _EVAL_5299;
  assign _EVAL_6076 = _EVAL_1145[669];
  assign _EVAL_408 = _EVAL_1159[23:17];
  assign _EVAL_5975 = _EVAL_4462 & _EVAL_1290;
  assign _EVAL_2893 = _EVAL_1146 & _EVAL_3487;
  assign _EVAL_1050 = _EVAL_298 & _EVAL_5464;
  assign _EVAL_364 = ~_EVAL_2589;
  assign _EVAL_4817 = _EVAL_1145[536];
  assign _EVAL_3057 = _EVAL_5074 & _EVAL_2695;
  assign _EVAL_2304 = _EVAL_5074 & _EVAL_206;
  assign _EVAL_1663 = _EVAL_5370 & _EVAL_369;
  assign _EVAL_3698 = _EVAL_3961 & _EVAL_2969;
  assign _EVAL_4450 = _EVAL_4692 & _EVAL_3154;
  assign _EVAL_5458 = _EVAL_451 & _EVAL_5753;
  assign _EVAL_5401 = _EVAL_2341 & _EVAL_3447;
  assign _EVAL_911 = _EVAL_4987 & _EVAL_5299;
  assign _EVAL_5179 = _EVAL_3553 & _EVAL_3284;
  assign _EVAL_964 = _EVAL_3202 & _EVAL_3702;
  assign _EVAL_4435 = _EVAL_4311 & _EVAL_3766;
  assign _EVAL_3489 = _EVAL_2005 & _EVAL_5543;
  assign _EVAL_3778 = _EVAL_5100 & _EVAL_1735;
  assign _EVAL_4491 = _EVAL_2585 & _EVAL_3154;
  assign _EVAL_5747 = _EVAL_3992 & _EVAL_1924;
  assign _EVAL_1605 = _EVAL_831 & _EVAL_5543;
  assign _EVAL_984 = _EVAL_610 & _EVAL_3379;
  assign _EVAL_299 = _EVAL_3981 & _EVAL_3398;
  assign _EVAL_2924 = _EVAL_3451 & _EVAL_3398;
  assign _EVAL_3458 = _EVAL_5766 & _EVAL_1009;
  assign _EVAL_4559 = _EVAL_4224 & _EVAL_1735;
  assign _EVAL_5831 = ~_EVAL_1407;
  assign _EVAL_2478 = _EVAL_3456 & _EVAL_327;
  assign _EVAL_2863 = _EVAL_3651 & _EVAL_3702;
  assign _EVAL_1837 = _EVAL_965 & _EVAL_3313;
  assign _EVAL_710 = _EVAL_3451 & _EVAL_882;
  assign _EVAL_1574 = _EVAL_3935 & _EVAL_2748;
  assign _EVAL_1421 = _EVAL_4078 & _EVAL_2424;
  assign _EVAL_200 = _EVAL_5028 & _EVAL_4109;
  assign _EVAL_1936 = _EVAL_5132 & _EVAL_3398;
  assign _EVAL_3081 = _EVAL_251 & _EVAL_369;
  assign _EVAL_496 = _EVAL_4202 & _EVAL_801;
  assign _EVAL_207 = _EVAL_5528 & _EVAL_587;
  assign _EVAL_1193 = _EVAL_4604 & _EVAL_1290;
  assign _EVAL_3873 = _EVAL_921 & _EVAL_847;
  assign _EVAL_5454 = _EVAL_5561 & _EVAL_2077;
  assign _EVAL_4112 = _EVAL_309 & _EVAL_1735;
  assign _EVAL_1721 = _EVAL_921 & _EVAL_3398;
  assign _EVAL_4963 = _EVAL_529 & _EVAL_2956;
  assign _EVAL_3248 = _EVAL_1622 & _EVAL_5753;
  assign _EVAL_3066 = _EVAL_5074 & _EVAL_936;
  assign _EVAL_1642 = _EVAL_1655 & _EVAL_3154;
  assign _EVAL_4957 = _EVAL_5192 & _EVAL_369;
  assign _EVAL_645 = _EVAL_3436 & _EVAL_4788;
  assign _EVAL_4985 = _EVAL_434 & _EVAL_3261;
  assign _EVAL_5633 = _EVAL_961 & _EVAL_1488;
  assign _EVAL_3957 = _EVAL_3710 & _EVAL_1488;
  assign _EVAL_5914 = _EVAL_5246 & _EVAL_882;
  assign _EVAL_3754 = _EVAL_479 & _EVAL_3702;
  assign _EVAL_2370 = _EVAL_4627 & _EVAL_739;
  assign _EVAL_2471 = _EVAL_5912 & _EVAL_673;
  assign _EVAL_1103 = _EVAL_1386 & _EVAL_3379;
  assign _EVAL_4222 = _EVAL_6096 & _EVAL_673;
  assign _EVAL_862 = _EVAL_3130 & _EVAL_369;
  assign _EVAL_2923 = _EVAL_5450 & _EVAL_2382;
  assign _EVAL_4962 = _EVAL_984 & _EVAL_5299;
  assign _EVAL_282 = _EVAL_2260 & _EVAL_882;
  assign _EVAL_4121 = _EVAL_1745 & _EVAL_1735;
  assign _EVAL_3436 = _EVAL_5223 & _EVAL_1333;
  assign _EVAL_2126 = _EVAL_5074 & _EVAL_3038;
  assign _EVAL_380 = _EVAL_584 & _EVAL_4788;
  assign _EVAL_1363 = _EVAL_1145[518];
  assign _EVAL_938 = _EVAL_5068[530];
  assign _EVAL_2525 = _EVAL_1145[584];
  assign _EVAL_1977 = _EVAL_5074 & _EVAL_1426;
  assign _EVAL_5417 = _EVAL_1370 & _EVAL_4477;
  assign _EVAL_859 = _EVAL_3363 & _EVAL_704;
  assign _EVAL_5398 = _EVAL_2210 & _EVAL_3379;
  assign _EVAL_3826 = _EVAL_2327 & _EVAL_3379;
  assign _EVAL_5538 = _EVAL_4488 & _EVAL_882;
  assign _EVAL_4152 = _EVAL_1312 & _EVAL_369;
  assign _EVAL_1755 = _EVAL_5184 & _EVAL_5289;
  assign _EVAL_5650 = _EVAL_1971 & _EVAL_3702;
  assign _EVAL_3486 = _EVAL_1146 & _EVAL_3398;
  assign _EVAL_201 = _EVAL_4841 & _EVAL_3398;
  assign _EVAL_3536 = _EVAL_4499 & _EVAL_5850;
  assign _EVAL_1061 = _EVAL_5893 & _EVAL_2748;
  assign _EVAL_5722 = _EVAL_932 & _EVAL_2956;
  assign _EVAL_2271 = _EVAL_4795 & _EVAL_3702;
  assign _EVAL_5268 = _EVAL_2702 & _EVAL_5281;
  assign _EVAL_4283 = _EVAL_1971 & _EVAL_369;
  assign _EVAL_4146 = _EVAL_1312 & _EVAL_2424;
  assign _EVAL_4361 = _EVAL_2998 & _EVAL_3418;
  assign _EVAL_2297 = _EVAL_528 & _EVAL_1735;
  assign _EVAL_2466 = _EVAL_5924 & _EVAL_1395;
  assign _EVAL_5575 = _EVAL_5528 & _EVAL_4664;
  assign _EVAL_3932 = _EVAL_434 & _EVAL_3398;
  assign _EVAL_761 = _EVAL_124[0];
  assign _EVAL_5685 = _EVAL_3414 & _EVAL_1488;
  assign _EVAL_1811 = _EVAL_2335 & _EVAL_5299;
  assign _EVAL_3440 = _EVAL_4078 & _EVAL_2748;
  assign _EVAL_388 = _EVAL_4235 & _EVAL_3702;
  assign _EVAL_3586 = _EVAL_1316[3:0];
  assign _EVAL_2483 = _EVAL_4222 & _EVAL_3154;
  assign _EVAL_1313 = _EVAL_1920 & _EVAL_882;
  assign _EVAL_5987 = _EVAL_1446 & _EVAL_2748;
  assign _EVAL_4887 = _EVAL_4222 & _EVAL_4477;
  assign _EVAL_4310 = _EVAL_2376 & _EVAL_3702;
  assign _EVAL_4235 = _EVAL_1661 & _EVAL_3379;
  assign _EVAL_2242 = _EVAL_1006 & _EVAL_3379;
  assign _EVAL_3708 = _EVAL_5398 & _EVAL_2424;
  assign _EVAL_2750 = _EVAL_1553 & _EVAL_5289;
  assign _EVAL_2403 = _EVAL_2215 & _EVAL_4287;
  assign _EVAL_1916 = _EVAL_5618 & _EVAL_1488;
  assign _EVAL_2302 = _EVAL_1136 & _EVAL_847;
  assign _EVAL_3850 = _EVAL_2905 & _EVAL_1801;
  assign _EVAL_3323 = _EVAL_4627 & _EVAL_378;
  assign _EVAL_5739 = _EVAL_1145[577];
  assign _EVAL_3316 = _EVAL_3202 & _EVAL_2424;
  assign _EVAL_4334 = _EVAL_4141 & _EVAL_5543;
  assign _EVAL_2116 = _EVAL_1553 & _EVAL_4775;
  assign _EVAL_2649 = _EVAL_5023 & _EVAL_3418;
  assign _EVAL_3478 = _EVAL_5561 & _EVAL_1352;
  assign _EVAL_1447 = _EVAL_3220 & _EVAL_369;
  assign _EVAL_298 = _EVAL_2390 & _EVAL_3379;
  assign _EVAL_886 = _EVAL_6022 & _EVAL_369;
  assign _EVAL_4720 = _EVAL_4627 & _EVAL_3616;
  assign _EVAL_5414 = _EVAL_3220 & _EVAL_5543;
  assign _EVAL_4239 = _EVAL_4187 & _EVAL_3313;
  assign _EVAL_3004 = _EVAL_4692 & _EVAL_847;
  assign _EVAL_2768 = _EVAL_4577 & _EVAL_5289;
  assign _EVAL_793 = _EVAL_5074 & _EVAL_2082;
  assign _EVAL_3592 = _EVAL_5285 & _EVAL_369;
  assign _EVAL_3571 = ~_EVAL_1510;
  assign _EVAL_629 = _EVAL_2868 & _EVAL_882;
  assign _EVAL_4132 = _EVAL_2550 & _EVAL_1009;
  assign _EVAL_4391 = _EVAL_1202 & _EVAL_3487;
  assign _EVAL_2451 = _EVAL_5162 & _EVAL_6084;
  assign _EVAL_4836 = _EVAL_4029 & _EVAL_3379;
  assign _EVAL_5974 = _EVAL_1536 & _EVAL_2424;
  assign _EVAL_3611 = _EVAL_4149 & _EVAL_369;
  assign _EVAL_5911 = _EVAL_1344 & _EVAL_3418;
  assign _EVAL_5091 = _EVAL_4192 & _EVAL_3702;
  assign _EVAL_4048 = _EVAL_4078 & _EVAL_6084;
  assign _EVAL_4409 = _EVAL_1206 & _EVAL_1185;
  assign _EVAL_5798 = _EVAL_4745 & _EVAL_882;
  assign _EVAL_1149 = _EVAL_2673 & _EVAL_3379;
  assign _EVAL_3545 = _EVAL_4584 & _EVAL_1516;
  assign _EVAL_5755 = _EVAL_1962 & _EVAL_2956;
  assign _EVAL_2650 = _EVAL_3130 & _EVAL_2424;
  assign _EVAL_1657 = _EVAL_1136 & _EVAL_3418;
  assign _EVAL_1134 = _EVAL_4137 & _EVAL_3154;
  assign _EVAL_2039 = _EVAL_2986 & _EVAL_5464;
  assign _EVAL_5447 = _EVAL_5440 & _EVAL_847;
  assign _EVAL_5443 = _EVAL_5561 & _EVAL_4167;
  assign _EVAL_654 = _EVAL_263 & _EVAL_1198;
  assign _EVAL_590 = _EVAL_5074 & _EVAL_3209;
  assign _EVAL_4609 = _EVAL_690 & _EVAL_2079;
  assign _EVAL_1145 = 1024'h1 << _EVAL_3485;
  assign _EVAL_3421 = _EVAL_4806 & _EVAL_673;
  assign _EVAL_4507 = _EVAL_2897 & _EVAL_3379;
  assign _EVAL_1499 = _EVAL_1234 & _EVAL_3702;
  assign _EVAL_5444 = _EVAL_921 & _EVAL_3487;
  assign _EVAL_1426 = _EVAL_1145[604];
  assign _EVAL_5839 = _EVAL_2675 & _EVAL_2969;
  assign _EVAL_1133 = _EVAL_5869 & _EVAL_3418;
  assign _EVAL_5021 = _EVAL_3859 & _EVAL_2956;
  assign _EVAL_3961 = _EVAL_3948 & _EVAL_3379;
  assign _EVAL_3972 = _EVAL_1689 & _EVAL_2969;
  assign _EVAL_2124 = _EVAL_486 & _EVAL_2748;
  assign _EVAL_2552 = _EVAL_386 & _EVAL_5543;
  assign _EVAL_5192 = _EVAL_175 & _EVAL_3379;
  assign _EVAL_2770 = _EVAL_284 & _EVAL_2969;
  assign _EVAL_2906 = _EVAL_538 & _EVAL_369;
  assign _EVAL_5124 = _EVAL_5054 & _EVAL_847;
  assign _EVAL_2771 = _EVAL_4661 & _EVAL_5289;
  assign _EVAL_5498 = _EVAL_668 & _EVAL_6084;
  assign _EVAL_5971 = _EVAL_2592 & _EVAL_369;
  assign _EVAL_4545 = _EVAL_434 & _EVAL_3487;
  assign _EVAL_530 = _EVAL_1145[673];
  assign _EVAL_3679 = _EVAL_5344 & _EVAL_1735;
  assign _EVAL_3684 = _EVAL_1145[521];
  assign _EVAL_2634 = _EVAL_1393 & _EVAL_6084;
  assign _EVAL_4652 = _EVAL_799 & _EVAL_369;
  assign _EVAL_4135 = _EVAL_88 == 3'h4;
  assign _EVAL_4139 = _EVAL_5561 & _EVAL_1072;
  assign _EVAL_3968 = _EVAL_3476 & _EVAL_369;
  assign _EVAL_2285 = _EVAL_3421 & _EVAL_3261;
  assign _EVAL_3707 = _EVAL_4909 & _EVAL_3508;
  assign _EVAL_5092 = _EVAL_1393 & _EVAL_2748;
  assign _EVAL_1586 = _EVAL_3512 & _EVAL_369;
  assign _EVAL_3208 = _EVAL_4581 & _EVAL_5299;
  assign _EVAL_3340 = _EVAL_1633 & _EVAL_2748;
  assign _EVAL_3908 = _EVAL_5063 & _EVAL_882;
  assign _EVAL_4420 = _EVAL_4974 & _EVAL_2382;
  assign _EVAL_4859 = _EVAL_2631 & _EVAL_882;
  assign _EVAL_2497 = _EVAL_537 & _EVAL_801;
  assign _EVAL_2937 = _EVAL_2005 & _EVAL_2969;
  assign _EVAL_2560 = _EVAL_589 & _EVAL_4751;
  assign _EVAL_1536 = _EVAL_492 & _EVAL_3379;
  assign _EVAL_4194 = _EVAL_1039 & _EVAL_3487;
  assign _EVAL_549 = _EVAL_4795 & _EVAL_5543;
  assign _EVAL_1393 = _EVAL_3492 & _EVAL_3379;
  assign _EVAL_3354 = _EVAL_5427 & _EVAL_3418;
  assign _EVAL_2941 = _EVAL_1145[535];
  assign _EVAL_4608 = _EVAL_1419 & _EVAL_369;
  assign _EVAL_6086 = _EVAL_5074 & _EVAL_1596;
  assign _EVAL_608 = _EVAL_3710 & _EVAL_3702;
  assign _EVAL_2875 = _EVAL_2910 & _EVAL_1270;
  assign _EVAL_1453 = _EVAL_1633 & _EVAL_2424;
  assign _EVAL_1845 = _EVAL_5788 & _EVAL_3170;
  assign _EVAL_2165 = _EVAL_4689 & _EVAL_4109;
  assign _EVAL_5103 = _EVAL_2986 & _EVAL_2382;
  assign _EVAL_2416 = _EVAL_1533 & _EVAL_4751;
  assign _EVAL_2614 = _EVAL_434 & _EVAL_882;
  assign _EVAL_1528 = _EVAL_5068[517];
  assign _EVAL_1077 = _EVAL_5795 & _EVAL_1290;
  assign _EVAL_2273 = _EVAL_5206 & _EVAL_3284;
  assign _EVAL_2962 = _EVAL_778 & _EVAL_4664;
  assign _EVAL_1471 = _EVAL_3993 & _EVAL_3261;
  assign _EVAL_4225 = _EVAL_1145[580];
  assign _EVAL_1326 = _EVAL_4083 & _EVAL_3398;
  assign _EVAL_1538 = _EVAL_537 & _EVAL_4788;
  assign _EVAL_4472 = _EVAL_528 & _EVAL_4108;
  assign _EVAL_4750 = _EVAL_4627 & _EVAL_5590;
  assign _EVAL_3396 = _EVAL_4144 & _EVAL_3284;
  assign _EVAL_4503 = _EVAL_3935 & _EVAL_2969;
  assign _EVAL_4157 = _EVAL_5148 & _EVAL_3702;
  assign _EVAL_1887 = _EVAL_3188 & _EVAL_4775;
  assign _EVAL_6054 = _EVAL_2607 & _EVAL_2956;
  assign _EVAL_4378 = _EVAL_3082 & _EVAL_6084;
  assign _EVAL_5336 = _EVAL_1960 & _EVAL_5289;
  assign _EVAL_1958 = _EVAL_807 & _EVAL_4775;
  assign _EVAL_3470 = _EVAL_4856 & _EVAL_369;
  assign _EVAL_6011 = _EVAL_5427 & _EVAL_847;
  assign _EVAL_5251 = _EVAL_2170 & _EVAL_1488;
  assign _EVAL_3376 = _EVAL_4623 & _EVAL_369;
  assign _EVAL_3522 = _EVAL_4795 & _EVAL_6084;
  assign _EVAL_3837 = _EVAL_4118 & _EVAL_3379;
  assign _EVAL_651 = _EVAL_3996 & _EVAL_4775;
  assign _EVAL_4788 = _EVAL_350 != 8'h0;
  assign _EVAL_1468 = _EVAL_124[1];
  assign _EVAL_473 = _EVAL_5893 & _EVAL_5543;
  assign _EVAL_5502 = _EVAL_5994 & _EVAL_4477;
  assign _EVAL_2699 = _EVAL_1620 & _EVAL_5850;
  assign _EVAL_6039 = _EVAL_3624 & _EVAL_369;
  assign _EVAL_3923 = _EVAL_1145[665];
  assign _EVAL_752 = _EVAL_3216 & _EVAL_3398;
  assign _EVAL_1432 = _EVAL_1553 & _EVAL_3766;
  assign _EVAL_1619 = _EVAL_1159[15:9];
  assign _EVAL_3978 = _EVAL_4745 & _EVAL_847;
  assign _EVAL_659 = _EVAL_4219 & _EVAL_3702;
  assign _EVAL_4949 = _EVAL_5893 & _EVAL_369;
  assign _EVAL_2695 = _EVAL_1145[576];
  assign _EVAL_4140 = _EVAL_5068[527];
  assign _EVAL_4745 = _EVAL_5116 & _EVAL_673;
  assign _EVAL_3562 = _EVAL_5074 & _EVAL_699;
  assign _EVAL_4670 = _EVAL_5819 & _EVAL_4664;
  assign _EVAL_830 = _EVAL_3052 & _EVAL_3154;
  assign _EVAL_4613 = _EVAL_3346 & _EVAL_3487;
  assign _EVAL_3326 = _EVAL_5542 & _EVAL_2320;
  assign _EVAL_5819 = _EVAL_1090 & _EVAL_673;
  assign _EVAL_1470 = _EVAL_1316[27:24];
  assign _EVAL_790 = _EVAL_1865 & _EVAL_4477;
  assign _EVAL_4850 = _EVAL_761 ? 8'hff : 8'h0;
  assign _EVAL_544 = _EVAL_302 & _EVAL_1488;
  assign _EVAL_1808 = ~_EVAL_1777;
  assign _EVAL_2072 = _EVAL_3414 & _EVAL_3702;
  assign _EVAL_908 = _EVAL_5561 & _EVAL_3564;
  assign _EVAL_3523 = _EVAL_4627 & _EVAL_347;
  assign _EVAL_2511 = _EVAL_3710 & _EVAL_6084;
  assign _EVAL_3244 = _EVAL_1103 & _EVAL_5543;
  assign _EVAL_2588 = _EVAL_935 & _EVAL_5543;
  assign _EVAL_4565 = _EVAL_4627 & _EVAL_530;
  assign _EVAL_5737 = _EVAL_3704 & _EVAL_4751;
  assign _EVAL_3085 = _EVAL_4219 & _EVAL_5543;
  assign _EVAL_4703 = _EVAL_1145[607];
  assign _EVAL_5476 = _EVAL_4707 & _EVAL_5289;
  assign _EVAL_4764 = _EVAL_4627 & _EVAL_3186;
  assign _EVAL_2542 = _EVAL_6033 & _EVAL_5289;
  assign _EVAL_4141 = _EVAL_3054 & _EVAL_3379;
  assign _EVAL_177 = _EVAL_1145[544];
  assign _EVAL_2310 = _EVAL_5028 & _EVAL_2382;
  assign _EVAL_2409 = _EVAL_1675 & _EVAL_1488;
  assign _EVAL_3568 = _EVAL_1149 & _EVAL_369;
  assign _EVAL_5566 = _EVAL_4627 & _EVAL_1426;
  assign _EVAL_5927 = ~_EVAL_4397;
  assign _EVAL_3956 = _EVAL_1364 & _EVAL_5299;
  assign _EVAL_389 = _EVAL_2454 & _EVAL_4751;
  assign _EVAL_626 = _EVAL_124[2];
  assign _EVAL_2753 = _EVAL_4986[21:0];
  assign _EVAL_4419 = _EVAL_3648 & _EVAL_673;
  assign _EVAL_1824 = _EVAL_1145[532];
  assign _EVAL_4524 = _EVAL_5068[544];
  assign _EVAL_3462 = _EVAL_2868 & _EVAL_847;
  assign _EVAL_2975 = _EVAL_1145[649];
  assign _EVAL_1269 = _EVAL_5705 & _EVAL_5543;
  assign _EVAL_1152 = _EVAL_5148 & _EVAL_369;
  assign _EVAL_3497 = _EVAL_831 & _EVAL_369;
  assign _EVAL_3558 = ~_EVAL_1293;
  assign _EVAL_5194 = ~_EVAL_3914;
  assign _EVAL_757 = _EVAL_1146 & _EVAL_3418;
  assign _EVAL_529 = _EVAL_1355 & _EVAL_3379;
  assign _EVAL_5184 = _EVAL_4793 & _EVAL_673;
  assign _EVAL_2207 = _EVAL_4757 & _EVAL_3487;
  assign _EVAL_4006 = _EVAL_3928 & _EVAL_3398;
  assign _EVAL_2593 = _EVAL_4627 & _EVAL_413;
  assign _EVAL_2288 = _EVAL_4627 & _EVAL_5201;
  assign _EVAL_5226 = _EVAL_5162 & _EVAL_2748;
  assign _EVAL_1756 = _EVAL_475 & _EVAL_1198;
  assign _EVAL_5673 = _EVAL_3928 & _EVAL_847;
  assign _EVAL_6093 = _EVAL_5370 & _EVAL_2969;
  assign _EVAL_2362 = ~_EVAL_2766;
  assign _EVAL_1972 = _EVAL_2753[3];
  assign _EVAL_926 = ~_EVAL_5735;
  assign _EVAL_5543 = _EVAL_1316[8];
  assign _EVAL_5892 = _EVAL_362 & _EVAL_3766;
  assign _EVAL_6070 = _EVAL_2154 & _EVAL_4686;
  assign _EVAL_503 = _EVAL_4783 & _EVAL_5543;
  assign _EVAL_187 = _EVAL_4618 & _EVAL_587;
  assign _EVAL_555 = _EVAL_5819 & _EVAL_587;
  assign _EVAL_4097 = _EVAL_1145[546];
  assign _EVAL_1116 = _EVAL_3993 & _EVAL_3154;
  assign _EVAL_5387 = _EVAL_302 & _EVAL_2969;
  assign _EVAL_351 = _EVAL_2009 & _EVAL_3583;
  assign _EVAL_2886 = _EVAL_2170 & _EVAL_2969;
  assign _EVAL_1241 = _EVAL_4078 & _EVAL_5543;
  assign _EVAL_4896 = _EVAL_538 & _EVAL_2424;
  assign _EVAL_2290 = _EVAL_807 & _EVAL_587;
  assign _EVAL_5850 = _EVAL_5922 != 4'h0;
  assign _EVAL_3844 = _EVAL_4939 & _EVAL_3379;
  assign _EVAL_4300 = _EVAL_4219 & _EVAL_2969;
  assign _EVAL_6057 = _EVAL_5994 & _EVAL_3418;
  assign _EVAL_4091 = _EVAL_1500 & _EVAL_3398;
  assign _EVAL_5434 = _EVAL_2242 & _EVAL_6084;
  assign _EVAL_2724 = _EVAL_799 & _EVAL_2748;
  assign _EVAL_5656 = _EVAL_1145[660];
  assign _EVAL_4643 = _EVAL_5450 & _EVAL_4751;
  assign _EVAL_854 = _EVAL_5068[546];
  assign _EVAL_2675 = _EVAL_3695 & _EVAL_3379;
  assign _EVAL_4592 = _EVAL_2037 & _EVAL_3702;
  assign _EVAL_2298 = _EVAL_4083 & _EVAL_3261;
  assign _EVAL_3574 = _EVAL_1176 & _EVAL_3379;
  assign _EVAL_1226 = ~_EVAL_2301;
  assign _EVAL_3828 = _EVAL_616 & _EVAL_5456;
  assign _EVAL_2836 = _EVAL_3421 & _EVAL_3487;
  assign _EVAL_4063 = _EVAL_3188 & _EVAL_587;
  assign _EVAL_3998 = _EVAL_523 != 8'h0;
  assign _EVAL_1563 = _EVAL_3226 & _EVAL_5850;
  assign _EVAL_3328 = _EVAL_2254 & _EVAL_2748;
  assign _EVAL_3180 = _EVAL_1553 & _EVAL_4664;
  assign _EVAL_2732 = _EVAL_2037 & _EVAL_369;
  assign TLMonitor__EVAL_11 = Queue__EVAL_14;
  assign _EVAL_378 = _EVAL_1145[542];
  assign _EVAL_5284 = _EVAL_5795 & _EVAL_5289;
  assign _EVAL_4455 = _EVAL_4627 & _EVAL_1411;
  assign _EVAL_3167 = _EVAL_5998 & _EVAL_5464;
  assign _EVAL_4629 = _EVAL_5561 & _EVAL_4524;
  assign _EVAL_5025 = _EVAL_1039 & _EVAL_3261;
  assign _EVAL_4270 = _EVAL_3920 & _EVAL_3766;
  assign _EVAL_2125 = _EVAL_2868 & _EVAL_3418;
  assign _EVAL_262 = _EVAL_5930 & _EVAL_3702;
  assign _EVAL_4180 = _EVAL_4106 & _EVAL_5289;
  assign _EVAL_2475 = _EVAL_3837 & _EVAL_369;
  assign _EVAL_4232 = _EVAL_5440 & _EVAL_4477;
  assign _EVAL_3624 = _EVAL_5956 & _EVAL_3379;
  assign _EVAL_4674 = _EVAL_3866 & _EVAL_2612;
  assign _EVAL_688 = _EVAL_2340 & _EVAL_673;
  assign _EVAL_4191 = _EVAL_5930 & _EVAL_6084;
  assign _EVAL_2730 = _EVAL_921 & _EVAL_3154;
  assign _EVAL_3782 = _EVAL_3226 & _EVAL_4109;
  assign _EVAL_680 = _EVAL_5561 & _EVAL_1465;
  assign _EVAL_2612 = ~_EVAL_3196;
  assign _EVAL_4093 = _EVAL_4332 & _EVAL_673;
  assign _EVAL_4101 = _EVAL_1145[590];
  assign _EVAL_3803 = _EVAL_4311 & _EVAL_1290;
  assign _EVAL_1653 = _EVAL_334 == 8'hff;
  assign _EVAL_1029 = ~_EVAL_1670;
  assign _EVAL_2321 = _EVAL_4254 & _EVAL_3766;
  assign _EVAL_4223 = _EVAL_2260 & _EVAL_3154;
  assign _EVAL_4991 = _EVAL_386 & _EVAL_2969;
  assign _EVAL_5236 = _EVAL_1145[585];
  assign _EVAL_1876 = _EVAL_4439 & _EVAL_673;
  assign _EVAL_925 = _EVAL_1145[256];
  assign _EVAL_5343 = _EVAL_6007 & _EVAL_3418;
  assign _EVAL_6015 = _EVAL_2242 & _EVAL_2969;
  assign _EVAL_5418 = _EVAL_1229 & _EVAL_328;
  assign _EVAL_4856 = _EVAL_5043 & _EVAL_3379;
  assign _EVAL_2983 = _EVAL_1145[531];
  assign _EVAL_5229 = _EVAL_1223 & _EVAL_3702;
  assign _EVAL_768 = _EVAL_5074 & _EVAL_2397;
  assign _EVAL_4230 = _EVAL_2335 & _EVAL_1198;
  assign _EVAL_1380 = _EVAL_857 & _EVAL_3702;
  assign _EVAL_3955 = _EVAL_3524 & _EVAL_2748;
  assign _EVAL_2169 = _EVAL_1677 & _EVAL_3418;
  assign _EVAL_4917 = _EVAL_1675 & _EVAL_2424;
  assign _EVAL_6029 = _EVAL_4821 & _EVAL_369;
  assign _EVAL_268 = _EVAL_4137 & _EVAL_882;
  assign _EVAL_3276 = _EVAL_3202 & _EVAL_5543;
  assign _EVAL_2266 = _EVAL_4044 & _EVAL_882;
  assign _EVAL_4981 = ~_EVAL_454;
  assign _EVAL_4295 = _EVAL_362 & _EVAL_5753;
  assign _EVAL_331 = _EVAL_4042 & _EVAL_2320;
  assign _EVAL_2278 = _EVAL_4254 & _EVAL_1009;
  assign _EVAL_5412 = _EVAL_2585 & _EVAL_4477;
  assign _EVAL_3221 = _EVAL_4766 | _EVAL_24;
  assign _EVAL_3109 = ~_EVAL_484;
  assign _EVAL_491 = _EVAL_1865 & _EVAL_882;
  assign _EVAL_1446 = _EVAL_5016 & _EVAL_3379;
  assign _EVAL_5423 = _EVAL_1633 & _EVAL_2969;
  assign _EVAL_5734 = _EVAL_3928 & _EVAL_882;
  assign _EVAL_5882 = _EVAL_905 & _EVAL_3398;
  assign _EVAL_4975 = _EVAL_2731 & _EVAL_5543;
  assign _EVAL_1350 = _EVAL_5305 & _EVAL_3284;
  assign _EVAL_3240 = _EVAL_4224 & _EVAL_4751;
  assign _EVAL_4960 = _EVAL_1242 & _EVAL_3487;
  assign _EVAL_4422 = _EVAL_2254 & _EVAL_3702;
  assign _EVAL_4619 = _EVAL_1034 & _EVAL_5299;
  assign _EVAL_1394 = _EVAL_3070 & _EVAL_3284;
  assign _EVAL_577 = _EVAL_3052 & _EVAL_3261;
  assign _EVAL_5510 = _EVAL_5561 & _EVAL_2150;
  assign _EVAL_1483 = _EVAL_1876 & _EVAL_3261;
  assign _EVAL_801 = _EVAL_3048 != 8'h0;
  assign _EVAL_4044 = _EVAL_5252 & _EVAL_673;
  assign _EVAL_1006 = _EVAL_4627 & _EVAL_5739;
  assign _EVAL_2088 = _EVAL_5561 & _EVAL_1948;
  assign _EVAL_1243 = _EVAL_1745 & _EVAL_4109;
  assign _EVAL_2745 = _EVAL_2725 & _EVAL_882;
  assign _EVAL_631 = _EVAL_1393 & _EVAL_2969;
  assign _EVAL_2011 = _EVAL_1370 & _EVAL_3398;
  assign _EVAL_3077 = _EVAL_4627 & _EVAL_3528;
  assign _EVAL_5372 = _EVAL_1960 & _EVAL_4775;
  assign _EVAL_4910 = _EVAL_5074 & _EVAL_1558;
  assign _EVAL_6010 = _EVAL_4419 & _EVAL_4477;
  assign _EVAL_4366 = _EVAL_1655 & _EVAL_4477;
  assign _EVAL_4873 = _EVAL_3130 & _EVAL_3702;
  assign _EVAL_4625 = _EVAL_1418 & _EVAL_3379;
  assign _EVAL_4038 = _EVAL_4757 & _EVAL_3418;
  assign _EVAL_457 = _EVAL_4785 & _EVAL_1840;
  assign _EVAL_3065 = _EVAL_446 & _EVAL_3284;
  assign _EVAL_4790 = _EVAL_2471 & _EVAL_4477;
  assign _EVAL_5060 = _EVAL_1419 & _EVAL_5543;
  assign _EVAL_3245 = _EVAL_5549 & _EVAL_1198;
  assign _EVAL_1562 = _EVAL_1145[603];
  assign _EVAL_3552 = _EVAL_4909 & _EVAL_3998;
  assign _EVAL_1401 = _EVAL_4083 & _EVAL_3154;
  assign _EVAL_6069 = _EVAL_4627 & _EVAL_2941;
  assign _EVAL_2625 = _EVAL_4563 & _EVAL_1488;
  assign _EVAL_154 = _EVAL_2106 & _EVAL_369;
  assign _EVAL_5921 = _EVAL_3574 & _EVAL_3998;
  assign _EVAL_4635 = _EVAL_1067 & _EVAL_5289;
  assign _EVAL_3520 = _EVAL_5155 & _EVAL_2748;
  assign _EVAL_1558 = _EVAL_1145[671];
  assign _EVAL_3746 = _EVAL_828 & _EVAL_1735;
  assign _EVAL_950 = _EVAL_4689 & _EVAL_5850;
  assign _EVAL_1836 = _EVAL_1344 & _EVAL_882;
  assign _EVAL_1139 = _EVAL_4707 & _EVAL_5753;
  assign _EVAL_5083 = _EVAL_1625 & _EVAL_2969;
  assign _EVAL_4077 = ~_EVAL_506;
  assign _EVAL_1685 = _EVAL_3202 & _EVAL_2969;
  assign _EVAL_3095 = _EVAL_1234 & _EVAL_2748;
  assign _EVAL_894 = _EVAL_434 & _EVAL_847;
  assign _EVAL_2976 = _EVAL_5440 & _EVAL_3261;
  assign _EVAL_682 = _EVAL_4692 & _EVAL_3418;
  assign _EVAL_4111 = _EVAL_362 & _EVAL_587;
  assign _EVAL_2083 = _EVAL_5662 & _EVAL_3154;
  assign _EVAL_1801 = ~_EVAL_1544;
  assign _EVAL_868 = _EVAL_5598 & _EVAL_3261;
  assign _EVAL_2860 = _EVAL_4078 & _EVAL_369;
  assign _EVAL_1475 = _EVAL_1316[15:8];
  assign _EVAL_5028 = _EVAL_2582 & _EVAL_3379;
  assign _EVAL_5634 = _EVAL_2877 & _EVAL_2969;
  assign _EVAL_1340 = ~_EVAL_5307;
  assign _EVAL_1590 = _EVAL_4627 & _EVAL_241;
  assign _EVAL_191 = _EVAL_4856 & _EVAL_2424;
  assign _EVAL_2746 = _EVAL_3928 & _EVAL_4477;
  assign _EVAL_4196 = _EVAL_4870 & _EVAL_2956;
  assign _EVAL_3398 = _EVAL_1619 != 7'h0;
  assign _EVAL_3135 = _EVAL_6007 & _EVAL_847;
  assign _EVAL_5057 = _EVAL_1202 & _EVAL_847;
  assign _EVAL_4777 = _EVAL_2471 & _EVAL_847;
  assign _EVAL_2254 = _EVAL_5979 & _EVAL_3379;
  assign _EVAL_1478 = _EVAL_5063 & _EVAL_847;
  assign _EVAL_2850 = _EVAL_5074 & _EVAL_2991;
  assign _EVAL_3122 = _EVAL_4235 & _EVAL_1488;
  assign _EVAL_2021 = _EVAL_2292 & _EVAL_4751;
  assign _EVAL_172 = _EVAL_5023 & _EVAL_3261;
  assign _EVAL_3252 = _EVAL_3220 & _EVAL_2969;
  assign _EVAL_572 = _EVAL_5305 & _EVAL_2956;
  assign _EVAL_3818 = _EVAL_5353 & _EVAL_6084;
  assign _EVAL_4596 = _EVAL_680 & _EVAL_673;
  assign _EVAL_3461 = _EVAL_1145[644];
  assign _EVAL_386 = _EVAL_5525 & _EVAL_3379;
  assign _EVAL_4765 = _EVAL_5998 & _EVAL_5850;
  assign _EVAL_4681 = _EVAL_5998 & _EVAL_2382;
  assign _EVAL_2835 = _EVAL_2100 & _EVAL_3154;
  assign _EVAL_2236 = _EVAL_1316[31:28];
  assign _EVAL_2817 = _EVAL_5068[541];
  assign _EVAL_4211 = _EVAL_774 & _EVAL_1488;
  assign _EVAL_3166 = _EVAL_1082 & _EVAL_3702;
  assign _EVAL_2150 = _EVAL_5068[538];
  assign _EVAL_5328 = _EVAL_1689 & _EVAL_2748;
  assign _EVAL_4579 = _EVAL_3181 & _EVAL_462;
  assign _EVAL_5569 = _EVAL_6088 != 31'h0;
  assign _EVAL_4258 = _EVAL_3992 & _EVAL_1653;
  assign _EVAL_1324 = _EVAL_386 & _EVAL_6084;
  assign _EVAL_5736 = _EVAL_2583 & _EVAL_722;
  assign _EVAL_3295 = _EVAL_5561 & _EVAL_4162;
  assign _EVAL_1985 = _EVAL_5184 & _EVAL_4775;
  assign _EVAL_1734 = _EVAL_1620 & _EVAL_5464;
  assign _EVAL_5838 = _EVAL_5068[534];
  assign _EVAL_2799 = _EVAL_4625 & _EVAL_369;
  assign _EVAL_3677 = _EVAL_1149 & _EVAL_1488;
  assign _EVAL_3307 = _EVAL_434 & _EVAL_3418;
  assign _EVAL_4947 = _EVAL_4627 & _EVAL_633;
  assign _EVAL_4362 = _EVAL_5369 & _EVAL_5230;
  assign _EVAL_1931 = _EVAL_4757 & _EVAL_882;
  assign _EVAL_3029 = _EVAL_5028 & _EVAL_3170;
  assign _EVAL_5593 = _EVAL_1145[674];
  assign _EVAL_1830 = _EVAL_5398 & _EVAL_2748;
  assign _EVAL_3015 = ~_EVAL_5781;
  assign _EVAL_1009 = _EVAL_3882 != 4'h0;
  assign _EVAL_2015 = ~_EVAL_3327;
  assign _EVAL_842 = _EVAL_4596 & _EVAL_587;
  assign _EVAL_568 = _EVAL_1159[11:8];
  assign _EVAL_3787 = _EVAL_4139 & _EVAL_673;
  assign _EVAL_4557 = _EVAL_3844 & _EVAL_5543;
  assign _EVAL_6089 = _EVAL_5561 & _EVAL_3985;
  assign _EVAL_5652 = _EVAL_504 & _EVAL_1198;
  assign _EVAL_1161 = _EVAL_3837 & _EVAL_2424;
  assign _EVAL_6094 = _EVAL_3837 & _EVAL_3702;
  assign _EVAL_2814 = _EVAL_479 & _EVAL_2424;
  assign _EVAL_5733 = _EVAL_1145[524];
  assign _EVAL_1083 = _EVAL_3512 & _EVAL_2748;
  assign _EVAL_2295 = _EVAL_1039 & _EVAL_3398;
  assign TLMonitor__EVAL_1 = _EVAL_11;
  assign _EVAL_2902 = _EVAL_3445 & _EVAL_3379;
  assign _EVAL_4881 = _EVAL_668 & _EVAL_369;
  assign _EVAL_6097 = _EVAL_2725 & _EVAL_3154;
  assign _EVAL_1376 = _EVAL_5869 & _EVAL_3398;
  assign _EVAL_799 = _EVAL_1065 & _EVAL_3379;
  assign _EVAL_2733 = _EVAL_5561 & _EVAL_2706;
  assign _EVAL_3566 = _EVAL_1536 & _EVAL_5543;
  assign _EVAL_3198 = _EVAL_4987 & _EVAL_2956;
  assign _EVAL_2982 = _EVAL_4625 & _EVAL_2748;
  assign _EVAL_4673 = _EVAL_3476 & _EVAL_2748;
  assign _EVAL_4781 = _EVAL_6051 & _EVAL_1735;
  assign _EVAL_2504 = _EVAL_534 & _EVAL_4108;
  assign _EVAL_5702 = _EVAL_5676 & _EVAL_3487;
  assign _EVAL_1795 = _EVAL_581 & _EVAL_2956;
  assign _EVAL_3508 = _EVAL_1475 != 8'h0;
  assign _EVAL_3738 = _EVAL_4627 & _EVAL_5867;
  assign _EVAL_540 = _EVAL_284 & _EVAL_369;
  assign _EVAL_4488 = _EVAL_1000 & _EVAL_673;
  assign _EVAL_1946 = _EVAL_3364 & _EVAL_3398;
  assign _EVAL_1424 = _EVAL_4627 & _EVAL_1069;
  assign _EVAL_5148 = _EVAL_5879 & _EVAL_3379;
  assign _EVAL_5772 = _EVAL_4618 & _EVAL_5753;
  assign _EVAL_4293 = _EVAL_5068[514];
  assign _EVAL_4645 = _EVAL_3414 & _EVAL_369;
  assign _EVAL_1718 = _EVAL_3738 & _EVAL_3379;
  assign _EVAL_4220 = _EVAL_3183 & _EVAL_5543;
  assign _EVAL_4780 = _EVAL_1067 & _EVAL_587;
  assign _EVAL_464 = _EVAL_1145[654];
  assign _EVAL_2328 = _EVAL_4351 & _EVAL_3702;
  assign _EVAL_2536 = _EVAL_5561 & _EVAL_289;
  assign _EVAL_4439 = _EVAL_5561 & _EVAL_3211;
  assign _EVAL_5855 = _EVAL_4856 & _EVAL_3702;
  assign _EVAL_1234 = _EVAL_2655 & _EVAL_3379;
  assign _EVAL_287 = _EVAL_3421 & _EVAL_3418;
  assign _EVAL_4707 = _EVAL_4730 & _EVAL_673;
  assign _EVAL_3406 = _EVAL_3476 & _EVAL_3702;
  assign _EVAL_839 = _EVAL_3826 & _EVAL_5299;
  assign _EVAL_4601 = _EVAL_1145[610];
  assign _EVAL_622 = _EVAL_1145[578];
  assign _EVAL_4277 = _EVAL_932 & _EVAL_3284;
  assign _EVAL_1650 = _EVAL_2292 & _EVAL_5850;
  assign _EVAL_2662 = _EVAL_5598 & _EVAL_3487;
  assign _EVAL_5099 = _EVAL_2550 & _EVAL_4775;
  assign _EVAL_745 = _EVAL_528 & _EVAL_4109;
  assign _EVAL_2045 = _EVAL_4314 & _EVAL_5797;
  assign _EVAL_3112 = _EVAL_5077 & _EVAL_847;
  assign _EVAL_1033 = _EVAL_2192 & _EVAL_6084;
  assign _EVAL_2170 = _EVAL_1194 & _EVAL_3379;
  assign _EVAL_4506 = _EVAL_3226 & _EVAL_1735;
  assign _EVAL_6003 = _EVAL_897 & _EVAL_2956;
  assign _EVAL_2573 = _EVAL_5450 & _EVAL_4109;
  assign _EVAL_4862 = _EVAL_807 & _EVAL_5753;
  assign _EVAL_4691 = _EVAL_751 & _EVAL_369;
  assign _EVAL_5077 = _EVAL_2423 & _EVAL_673;
  assign _EVAL_3338 = _EVAL_1745 & _EVAL_3170;
  assign _EVAL_1991 = _EVAL_735 & _EVAL_1735;
  assign _EVAL_5228 = _EVAL_4577 & _EVAL_3766;
  assign _EVAL_5922 = _EVAL_1316[15:12];
  assign _EVAL_3161 = _EVAL_644 & _EVAL_4100;
  assign _EVAL_1798 = _EVAL_3421 & _EVAL_3154;
  assign _EVAL_5980 = _EVAL_1146 & _EVAL_847;
  assign _EVAL_1334 = _EVAL_4311 & _EVAL_1009;
  assign _EVAL_5578 = _EVAL_1533 & _EVAL_2320;
  assign _EVAL_2323 = _EVAL_5561 & _EVAL_1714;
  assign _EVAL_5761 = _EVAL_3981 & _EVAL_847;
  assign _EVAL_5796 = _EVAL_2702 & _EVAL_1924;
  assign _EVAL_5602 = _EVAL_4627 & _EVAL_210;
  assign _EVAL_3134 = _EVAL_251 & _EVAL_1488;
  assign _EVAL_3360 = _EVAL_1620 & _EVAL_2382;
  assign _EVAL_1661 = _EVAL_4627 & _EVAL_5932;
  assign _EVAL_3337 = _EVAL_5618 & _EVAL_369;
  assign _EVAL_418 = _EVAL_2242 & _EVAL_1488;
  assign _EVAL_1735 = _EVAL_323 != 4'h0;
  assign _EVAL_957 = _EVAL_2902 & _EVAL_5543;
  assign _EVAL_435 = _EVAL_2308 & _EVAL_3373;
  assign _EVAL_3279 = _EVAL_3624 & _EVAL_2424;
  assign _EVAL_1348 = _EVAL_2338 & _EVAL_2748;
  assign _EVAL_4931 = ~_EVAL_906;
  assign _EVAL_332 = _EVAL_1361 & _EVAL_882;
  assign _EVAL_4228 = _EVAL_1039 & _EVAL_882;
  assign _EVAL_5937 = _EVAL_1145[586];
  assign _EVAL_5991 = _EVAL_799 & _EVAL_1488;
  assign _EVAL_3500 = _EVAL_735 & _EVAL_4108;
  assign _EVAL_1094 = _EVAL_2592 & _EVAL_6084;
  assign _EVAL_2485 = _EVAL_5819 & _EVAL_5753;
  assign _EVAL_2205 = _EVAL_3089 & _EVAL_3379;
  assign _EVAL_5214 = _EVAL_4187 & _EVAL_1009;
  assign _EVAL_4060 = _EVAL_2335 & _EVAL_3284;
  assign _EVAL_2686 = _EVAL_1242 & _EVAL_4477;
  assign _EVAL_4193 = _EVAL_1149 & _EVAL_2424;
  assign _EVAL_1514 = _EVAL_5528 & _EVAL_5289;
  assign _EVAL_3032 = _EVAL_5036 & _EVAL_673;
  assign _EVAL_327 = ~_EVAL_5409;
  assign _EVAL_5968 = _EVAL_486 & _EVAL_5543;
  assign _EVAL_4454 = _EVAL_5353 & _EVAL_5543;
  assign _EVAL_5201 = _EVAL_1145[596];
  assign _EVAL_4655 = _EVAL_4707 & _EVAL_1290;
  assign _EVAL_2526 = _EVAL_4745 & _EVAL_3487;
  assign _EVAL_2842 = _EVAL_2850 & _EVAL_3379;
  assign _EVAL_1482 = _EVAL_4149 & _EVAL_2969;
  assign _EVAL_2334 = _EVAL_2148 & _EVAL_927;
  assign _EVAL_2665 = _EVAL_5561 & _EVAL_3230;
  assign _EVAL_2818 = _EVAL_2260 & _EVAL_4477;
  assign _EVAL_4891 = ~_EVAL_5255;
  assign _EVAL_867 = _EVAL_668 & _EVAL_1488;
  assign _EVAL_3370 = _EVAL_3130 & _EVAL_6084;
  assign _EVAL_1865 = _EVAL_4430 & _EVAL_673;
  assign _EVAL_4154 = _EVAL_1145[598];
  assign _EVAL_5666 = _EVAL_1876 & _EVAL_3418;
  assign _EVAL_967 = _EVAL_688 & _EVAL_3261;
  assign _EVAL_789 = _EVAL_6080 & _EVAL_4751;
  assign _EVAL_2679 = _EVAL_4974 & _EVAL_3170;
  assign _EVAL_5811 = _EVAL_3057 & _EVAL_3379;
  assign _EVAL_4259 = _EVAL_1145[640];
  assign _EVAL_2871 = _EVAL_4351 & _EVAL_5543;
  assign _EVAL_292 = _EVAL_3996 & _EVAL_1009;
  assign _EVAL_3632 = _EVAL_1980 & _EVAL_3379;
  assign _EVAL_4801 = _EVAL_309 & _EVAL_4751;
  assign _EVAL_1000 = _EVAL_5561 & _EVAL_3953;
  assign _EVAL_649 = _EVAL_3706 & _EVAL_2424;
  assign _EVAL_155 = _EVAL_4222 & _EVAL_3487;
  assign _EVAL_5789 = _EVAL_778 & _EVAL_1290;
  assign _EVAL_2032 = _EVAL_2251 & _EVAL_2748;
  assign _EVAL_5274 = _EVAL_5561 & _EVAL_1699;
  assign _EVAL_3159 = _EVAL_5998 & _EVAL_1735;
  assign _EVAL_2744 = _EVAL_4870 & _EVAL_1198;
  assign _EVAL_5880 = _EVAL_5246 & _EVAL_3487;
  assign _EVAL_5879 = _EVAL_4627 & _EVAL_2507;
  assign _EVAL_4082 = _EVAL_5023 & _EVAL_3398;
  assign _EVAL_1171 = _EVAL_4235 & _EVAL_6084;
  assign _EVAL_5320 = _EVAL_5023 & _EVAL_882;
  assign _EVAL_2269 = _EVAL_5370 & _EVAL_1488;
  assign _EVAL_5277 = _EVAL_6022 & _EVAL_3702;
  assign _EVAL_2209 = _EVAL_4692 & _EVAL_4477;
  assign _EVAL_5664 = _EVAL_6032 & _EVAL_2748;
  assign _EVAL_1459 = _EVAL_2550 & _EVAL_1290;
  assign _EVAL_1919 = _EVAL_2998 & _EVAL_847;
  assign _EVAL_3214 = _EVAL_5561 & _EVAL_3298;
  assign _EVAL_3160 = _EVAL_1234 & _EVAL_5543;
  assign _EVAL_4989 = _EVAL_778 & _EVAL_1009;
  assign _EVAL_4279 = ~_EVAL_3129;
  assign _EVAL_1525 = _EVAL_1718 & _EVAL_369;
  assign _EVAL_2617 = _EVAL_1945 & _EVAL_5289;
  assign _EVAL_5527 = _EVAL_5788 & _EVAL_4751;
  assign _EVAL_1487 = _EVAL_2242 & _EVAL_3702;
  assign _EVAL_4733 = _EVAL_3920 & _EVAL_5753;
  assign _EVAL_4380 = _EVAL_4567 & _EVAL_3154;
  assign _EVAL_585 = _EVAL_5994 & _EVAL_847;
  assign _EVAL_385 = _EVAL_6051 & _EVAL_3170;
  assign _EVAL_1448 = _EVAL_1649 & _EVAL_5543;
  assign _EVAL_4049 = _EVAL_2793 & _EVAL_3418;
  assign _EVAL_1841 = _EVAL_4627 & _EVAL_4341;
  assign _EVAL_1259 = _EVAL_2444 & _EVAL_2555;
  assign _EVAL_5466 = _EVAL_4149 & _EVAL_3702;
  assign _EVAL_3471 = ~_EVAL_1388;
  assign _EVAL_202 = _EVAL_5068[519];
  assign _EVAL_2890 = _EVAL_4563 & _EVAL_5543;
  assign _EVAL_613 = _EVAL_5676 & _EVAL_882;
  assign _EVAL_5241 = _EVAL_5068[526];
  assign _EVAL_4798 = _EVAL_2292 & _EVAL_3170;
  assign _EVAL_5376 = _EVAL_2675 & _EVAL_2748;
  assign _EVAL_1202 = _EVAL_3214 & _EVAL_673;
  assign _EVAL_3305 = _EVAL_2241 & _EVAL_2424;
  assign _EVAL_3768 = _EVAL_5854 & _EVAL_3284;
  assign _EVAL_997 = ~_EVAL_2825;
  assign _EVAL_2001 = _EVAL_4627 & _EVAL_4306;
  assign _EVAL_998 = _EVAL_3844 & _EVAL_2748;
  assign _EVAL_2570 = _EVAL_5561 & _EVAL_2377;
  assign _EVAL_1358 = _EVAL_4488 & _EVAL_3418;
  assign _EVAL_4639 = _EVAL_2607 & _EVAL_3284;
  assign _EVAL_2998 = _EVAL_1701 & _EVAL_673;
  assign _EVAL_740 = _EVAL_5930 & _EVAL_2748;
  assign _EVAL_5329 = _EVAL_3107 & _EVAL_5543;
  assign _EVAL_5281 = _EVAL_4551 == 8'hff;
  assign _EVAL_4812 = _EVAL_3346 & _EVAL_3154;
  assign _EVAL_2220 = _EVAL_620 & _EVAL_2382;
  assign _EVAL_4175 = _EVAL_5856 & _EVAL_673;
  assign _EVAL_5574 = _EVAL_1542 & _EVAL_3418;
  assign _EVAL_713 = _EVAL_4627 & _EVAL_4605;
  assign _EVAL_1561 = _EVAL_5766 & _EVAL_587;
  assign _EVAL_2292 = _EVAL_1199 & _EVAL_3379;
  assign _EVAL_972 = _EVAL_407 & _EVAL_1488;
  assign _EVAL_2000 = _EVAL_3052 & _EVAL_882;
  assign _EVAL_2646 = _EVAL_2002 & _EVAL_2892;
  assign _EVAL_5286 = _EVAL_1876 & _EVAL_3398;
  assign _EVAL_641 = _EVAL_4627 & _EVAL_3923;
  assign _EVAL_5576 = _EVAL_2252 & _EVAL_882;
  assign _EVAL_2653 = _EVAL_3070 & _EVAL_5299;
  assign _EVAL_2545 = _EVAL_4627 & _EVAL_2306;
  assign _EVAL_5814 = ~_EVAL_2669;
  assign _EVAL_2708 = _EVAL_6022 & _EVAL_2748;
  assign _EVAL_4689 = _EVAL_2455 & _EVAL_3379;
  assign _EVAL_4888 = _EVAL_2151 & _EVAL_3379;
  assign _EVAL_2705 = _EVAL_3414 & _EVAL_2424;
  assign _EVAL_5532 = _EVAL_479 & _EVAL_5543;
  assign _EVAL_263 = _EVAL_4830 & _EVAL_3379;
  assign _EVAL_4898 = _EVAL_2592 & _EVAL_3702;
  assign _EVAL_5497 = _EVAL_3632 & _EVAL_1735;
  assign _EVAL_2238 = _EVAL_4044 & _EVAL_3487;
  assign _EVAL_2581 = _EVAL_5788 & _EVAL_4109;
  assign _EVAL_4821 = _EVAL_2680 & _EVAL_3379;
  assign _EVAL_4002 = _EVAL_5795 & _EVAL_5753;
  assign _EVAL_5596 = _EVAL_5598 & _EVAL_4477;
  assign _EVAL_2927 = _EVAL_1553 & _EVAL_5753;
  assign _EVAL_2479 = _EVAL_4192 & _EVAL_5543;
  assign _EVAL_4934 = _EVAL_828 & _EVAL_3170;
  assign _EVAL_3781 = _EVAL_2100 & _EVAL_3261;
  assign _EVAL_213 = _EVAL_5054 & _EVAL_3398;
  assign _EVAL_1973 = _EVAL_1361 & _EVAL_4477;
  assign _EVAL_1971 = _EVAL_1274 & _EVAL_3379;
  assign _EVAL_2790 = _EVAL_2346 & _EVAL_4866;
  assign _EVAL_3267 = _EVAL_5074 & _EVAL_885;
  assign _EVAL_4714 = _EVAL_3032 & _EVAL_3766;
  assign _EVAL_579 = _EVAL_620 & _EVAL_5464;
  assign _EVAL_1600 = _EVAL_3624 & _EVAL_2969;
  assign _EVAL_1270 = ~_EVAL_582;
  assign _EVAL_3292 = _EVAL_1281 & _EVAL_4160;
  assign _EVAL_396 = _EVAL_5846 & _EVAL_5831;
  assign _EVAL_1635 = _EVAL_3032 & _EVAL_1290;
  assign _EVAL_3433 = _EVAL_2241 & _EVAL_2969;
  assign _EVAL_228 = _EVAL_2725 & _EVAL_4477;
  assign _EVAL_2879 = _EVAL_2753[9];
  assign _EVAL_2670 = _EVAL_1655 & _EVAL_3261;
  assign _EVAL_1893 = _EVAL_302 & _EVAL_3702;
  assign _EVAL_832 = _EVAL_3226 & _EVAL_4108;
  assign _EVAL_2934 = _EVAL_5930 & _EVAL_5543;
  assign _EVAL_3155 = _EVAL_961 & _EVAL_6084;
  assign _EVAL_4806 = _EVAL_5561 & _EVAL_4140;
  assign _EVAL_5565 = _EVAL_3512 & _EVAL_2969;
  assign _EVAL_266 = _EVAL_1500 & _EVAL_847;
  assign _EVAL_4243 = _EVAL_5398 & _EVAL_5543;
  assign _EVAL_372 = _EVAL_4235 & _EVAL_2969;
  assign _EVAL_3379 = _EVAL_3264 == 22'h0;
  assign _EVAL_4868 = _EVAL_5342 & _EVAL_2956;
  assign _EVAL_2783 = ~_EVAL_2690;
  assign _EVAL_1948 = _EVAL_5068[518];
  assign _EVAL_3529 = _EVAL_4567 & _EVAL_3418;
  assign _EVAL_2031 = _EVAL_4137 & _EVAL_3398;
  assign _EVAL_3884 = _EVAL_1419 & _EVAL_3702;
  assign _EVAL_1869 = _EVAL_4821 & _EVAL_5543;
  assign _EVAL_2917 = _EVAL_6051 & _EVAL_4108;
  assign _EVAL_1889 = _EVAL_4707 & _EVAL_587;
  assign _EVAL_2554 = _EVAL_2793 & _EVAL_847;
  assign _EVAL_1615 = _EVAL_4604 & _EVAL_5289;
  assign _EVAL_3382 = _EVAL_386 & _EVAL_3702;
  assign _EVAL_316 = _EVAL_2972 & _EVAL_587;
  assign _EVAL_2659 = _EVAL_4618 & _EVAL_1290;
  assign _EVAL_1375 = _EVAL_5100 & _EVAL_4109;
  assign _EVAL_4389 = _EVAL_3130 & _EVAL_5543;
  assign _EVAL_224 = _EVAL_479 & _EVAL_2748;
  assign _EVAL_5250 = _EVAL_3052 & _EVAL_3418;
  assign _EVAL_2725 = _EVAL_2536 & _EVAL_673;
  assign TLMonitor__EVAL_14 = _EVAL_34;
  assign _EVAL_2822 = _EVAL_3996 & _EVAL_5753;
  assign _EVAL_3825 = _EVAL_5074 & _EVAL_3461;
  assign _EVAL_184 = _EVAL_769 & _EVAL_4535;
  assign _EVAL_2123 = _EVAL_1854 & _EVAL_3487;
  assign _EVAL_5084 = _EVAL_5561 & _EVAL_5516;
  assign _EVAL_1182 = _EVAL_4916 & _EVAL_4751;
  assign _EVAL_1494 = _EVAL_2205 & _EVAL_4751;
  assign _EVAL_462 = ~_EVAL_887;
  assign _EVAL_2007 = _EVAL_1542 & _EVAL_882;
  assign _EVAL_4712 = _EVAL_2972 & _EVAL_4664;
  assign _EVAL_5360 = _EVAL_1945 & _EVAL_4664;
  assign _EVAL_758 = _EVAL_5192 & _EVAL_3702;
  assign _EVAL_630 = _EVAL_1202 & _EVAL_3398;
  assign _EVAL_2100 = _EVAL_2088 & _EVAL_673;
  assign _EVAL_2632 = _EVAL_5068[521];
  assign _EVAL_2651 = _EVAL_6051 & _EVAL_2382;
  assign _EVAL_2482 = _EVAL_2454 & _EVAL_5850;
  assign _EVAL_2873 = _EVAL_2172 & _EVAL_3379;
  assign _EVAL_4775 = _EVAL_568 != 4'h0;
  assign _EVAL_4594 = _EVAL_5528 & _EVAL_1290;
  assign _EVAL_2911 = _EVAL_3815 & _EVAL_5464;
  assign _EVAL_421 = _EVAL_735 & _EVAL_4109;
  assign _EVAL_4369 = _EVAL_3156 & _EVAL_369;
  assign _EVAL_2326 = _EVAL_2731 & _EVAL_369;
  assign _EVAL_3021 = _EVAL_4618 & _EVAL_4664;
  assign _EVAL_4357 = _EVAL_620 & _EVAL_1735;
  assign _EVAL_2518 = _EVAL_4525 & _EVAL_4109;
  assign _EVAL_1233 = _EVAL_5994 & _EVAL_3261;
  assign _EVAL_1268 = _EVAL_5854 & _EVAL_1198;
  assign _EVAL_5127 = _EVAL_4175 & _EVAL_882;
  assign _EVAL_4832 = _EVAL_1316[23:20];
  assign _EVAL_1578 = _EVAL_2731 & _EVAL_3702;
  assign _EVAL_369 = _EVAL_1316[0];
  assign _EVAL_3933 = _EVAL_1971 & _EVAL_2424;
  assign _EVAL_781 = _EVAL_4627 & _EVAL_4656;
  assign _EVAL_5786 = _EVAL_4757 & _EVAL_3398;
  assign _EVAL_1986 = _EVAL_5074 & _EVAL_2306;
  assign _EVAL_2043 = _EVAL_4627 & _EVAL_398;
  assign _EVAL_4214 = _EVAL_2986 & _EVAL_1735;
  assign _EVAL_4151 = _EVAL_617 & _EVAL_1488;
  assign _EVAL_3658 = _EVAL_4462 & _EVAL_5753;
  assign _EVAL_5419 = _EVAL_4419 & _EVAL_3487;
  assign _EVAL_1036 = _EVAL_5398 & _EVAL_3702;
  assign _EVAL_4383 = _EVAL_4692 & _EVAL_3398;
  assign _EVAL_3474 = _EVAL_2986 & _EVAL_3170;
  assign _EVAL_808 = _EVAL_475 & _EVAL_3284;
  assign _EVAL_2272 = _EVAL_1649 & _EVAL_6084;
  assign _EVAL_1888 = ~_EVAL_3280;
  assign _EVAL_4306 = _EVAL_1145[668];
  assign _EVAL_4460 = _EVAL_5561 & _EVAL_4375;
  assign _EVAL_1392 = _EVAL_5561 & _EVAL_2300;
  assign _EVAL_3689 = _EVAL_4764 & _EVAL_3379;
  assign _EVAL_1283 = _EVAL_5998 & _EVAL_4109;
  assign _EVAL_5119 = ~_EVAL_24;
  assign _EVAL_2950 = ~_EVAL_2918;
  assign _EVAL_5437 = _EVAL_4372 & _EVAL_369;
  assign _EVAL_3287 = _EVAL_4507 & _EVAL_2956;
  assign _EVAL_589 = _EVAL_4424 & _EVAL_3379;
  assign _EVAL_5930 = _EVAL_922 & _EVAL_3379;
  assign _EVAL_3075 = _EVAL_5561 & _EVAL_5997;
  assign _EVAL_171 = _EVAL_2252 & _EVAL_3487;
  assign _EVAL_1399 = _EVAL_6007 & _EVAL_882;
  assign _EVAL_2684 = _EVAL_1765 & _EVAL_5641;
  assign _EVAL_4394 = _EVAL_769 & _EVAL_1391;
  assign _EVAL_3669 = _EVAL_774 & _EVAL_2969;
  assign _EVAL_695 = _EVAL_5642 & _EVAL_369;
  assign _EVAL_3106 = _EVAL_4044 & _EVAL_3398;
  assign _EVAL_3107 = _EVAL_4630 & _EVAL_3379;
  assign _EVAL_4332 = _EVAL_5561 & _EVAL_938;
  assign _EVAL_4083 = _EVAL_2657 & _EVAL_673;
  assign _EVAL_3812 = _EVAL_3032 & _EVAL_5753;
  assign _EVAL_4555 = _EVAL_1622 & _EVAL_5289;
  assign _EVAL_4278 = _EVAL_4175 & _EVAL_4477;
  assign _EVAL_5754 = _EVAL_5766 & _EVAL_5753;
  assign _EVAL_361 = _EVAL_828 & _EVAL_4109;
  assign _EVAL_5289 = _EVAL_5913 != 4'h0;
  assign _EVAL_3672 = _EVAL_4563 & _EVAL_2748;
  assign _EVAL_2181 = _EVAL_2170 & _EVAL_3702;
  assign _EVAL_284 = _EVAL_3314 & _EVAL_3379;
  assign _EVAL_1725 = _EVAL_2675 & _EVAL_3702;
  assign _EVAL_4125 = _EVAL_807 & _EVAL_5289;
  assign _EVAL_3898 = _EVAL_3060 & _EVAL_3379;
  assign _EVAL_5773 = _EVAL_5184 & _EVAL_1009;
  assign _EVAL_3695 = _EVAL_4627 & _EVAL_4101;
  assign _EVAL_3407 = _EVAL_3130 & _EVAL_2969;
  assign _EVAL_1366 = _EVAL_5618 & _EVAL_2424;
  assign _EVAL_4514 = _EVAL_5819 & _EVAL_4775;
  assign _EVAL_3139 = _EVAL_2121 & _EVAL_5005;
  assign _EVAL_3655 = _EVAL_5398 & _EVAL_6084;
  assign _EVAL_5620 = _EVAL_4042 & _EVAL_3998;
  assign _EVAL_3346 = _EVAL_4460 & _EVAL_673;
  assign _EVAL_1742 = _EVAL_2998 & _EVAL_4477;
  assign _EVAL_1055 = _EVAL_807 & _EVAL_4664;
  assign _EVAL_5316 = _EVAL_4254 & _EVAL_5289;
  assign _EVAL_4533 = _EVAL_623 & _EVAL_5543;
  assign _EVAL_625 = _EVAL_1370 & _EVAL_3261;
  assign _EVAL_4079 = _EVAL_3981 & _EVAL_882;
  assign _EVAL_4543 = _EVAL_3450 & _EVAL_2015;
  assign _EVAL_1316 = {_EVAL_3136,_EVAL_3420,_EVAL_4552,_EVAL_4850};
  assign _EVAL_4701 = _EVAL_3082 & _EVAL_2424;
  assign _EVAL_2305 = _EVAL_4627 & _EVAL_2093;
  assign _EVAL_1227 = _EVAL_407 & _EVAL_369;
  assign _EVAL_5088 = _EVAL_2252 & _EVAL_3418;
  assign _EVAL_712 = _EVAL_5077 & _EVAL_3398;
  assign _EVAL_2397 = _EVAL_1145[704];
  assign _EVAL_5945 = _EVAL_751 & _EVAL_2969;
  assign _EVAL_1988 = _EVAL_2585 & _EVAL_3261;
  always @(posedge _EVAL_106) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_429 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6a6f668)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1334 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb9fa6b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1741 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dfb8083)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5372 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8473bc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5135 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b8fc6f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_482 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1756 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55b9c162)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2498 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(758cb958)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3892 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8c89a8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4280 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d8b3251)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6071 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8be114b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_424 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4527 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee6422e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3853 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bdaca1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_465 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1460666a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2407 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66a12bf5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_659 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddb7c8c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2129 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6becc217)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4928 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5588 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aba328ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4422 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81879cd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4018 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39d8ad9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2758 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d545d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5127 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2105 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c027e865)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5282 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ea80ad6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4391 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d9e4e95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5188 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f752a53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b89b08a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_442 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c0bc693)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5671 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a50766e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6054 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71f8565b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1180 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a72668cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1940 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31d19c4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_884 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(813fb7e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_638 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80e60562)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4063 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2745630)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2851 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5667ba3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3094 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b91ad1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86798a6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4437 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3508578)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2499 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a92f191b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d207baf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1406 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b079f431)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4016 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3cd1912)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1909 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9b2e95e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3bc9634)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5362 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1851 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f59d898)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3434 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(364e0f9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5666 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3250 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1384 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fec9d68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1225 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(387eed1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2718 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2ee545)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2724 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65364693)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4294 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ca5c29c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2714 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2360bfc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2575 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a27e3b58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2613 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd98bba6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5331 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c744dda7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4787 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb027efe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5196 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(432f8743)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2345 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fca47b00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_825 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a65d57e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4691 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8417f0eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_900 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8622a0e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_380 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1289ef5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1283 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b5854b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5887 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd8d2fd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5259 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4790 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67332c04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2919 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2608 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64407b02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4739 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e79e7df5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1879 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9e0a23d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2022 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94518058)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5029 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df56667a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4011 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3feecab8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4876 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc6e7eda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5138 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5041 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e7d4061)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5993 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c92590a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3737 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a198bca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4996 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34b74e41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1122 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(160ddfcf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2789 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22c486ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5498 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2923 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a88bf7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2011 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5018 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45863aae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3a5aa13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4110 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23e2ec4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2222 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2908 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b707cc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3177 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9477f2f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1725 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d754e11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2103 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(497ecc0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2023 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1069a9f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1692 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(183c765b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4868 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(529a847e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3235 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4592 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6246761)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5959 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb886b9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4675 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7075f7b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5759 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd8af9c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3781 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3422 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(160d0932)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5326 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8161b9f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1916 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5082 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7622bd4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1697 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2849 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1884 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(310eb9bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1409 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5dcdbfe6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5730 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(221fd06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1259 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(513694be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1588 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3489b4b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1913 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b53e60b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1811 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(caed19c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1724 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa5fdfa9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2223 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68a7fe7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3138 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47330d18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1133 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1548 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f97fc8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5756 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21b2f0c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5357 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17312b2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3954 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1086 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc44a16e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5215 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a7f8a93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4423 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2368aeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3109 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2d4cd28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_987 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_389 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be173732)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1004 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ad1e6c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3457 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3720 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4737 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f99556d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4346 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_695 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(379bd7d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3285 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9e75e32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2630 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb445ec0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4413 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5857 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2723 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccc9041)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2266 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce30b9e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5643 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc80ae6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4295 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6f8c890)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5773 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28294c17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_200 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d7ed84c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4934 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f59052be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5340 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d2f8fc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5764 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e894bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5182 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ebecb08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5129 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96853bd3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1513 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d85dfcb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3999 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdb8992f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4113 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_914 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3030 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca3f3403)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_388 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20392bff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3788951b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4379 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(904f5055)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1169 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4887 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da29b4d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5559 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(186dc231)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_755 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cee6da3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9edf2d02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_819 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a25f9ddc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3296 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a05c069)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_764 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c16f1c62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_754 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ae473c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4381 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(875c1551)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b6ed464)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2965 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13b625f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1871 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(196e0307)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2116 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20b7446d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2833 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18865441)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5897 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d33bfb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1595 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18d7326d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4506 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c046015c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6c30e04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2445 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23b8fd88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2195 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5108 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbdc901c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4724 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3178 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_467 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1888bd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4039 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fc87e23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2510 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20f121d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1182 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e15c62f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2687 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d8594f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_985 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96e9fa52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1365 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e8c3a1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2097 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48ad49d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4305 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99bfcd5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2622 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86bb3730)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2494 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2795 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9660cf31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3061 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e38514e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5754 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96944c51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3835 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bc47eae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3792 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3da78d15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1405 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3241 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(685ebbd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4652 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a5f6880)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1247 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce97226c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5818 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(812200e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4270 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69de10c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5845 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1214 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(603b963a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1837 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1458 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b358728)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3360 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f552e03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_770 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4353 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5a07d06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4516 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2310 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84656c1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1743 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f0b2a49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2346 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac3155b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4138 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4871 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96588dc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3440 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd73a559)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3503 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e74128c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1911 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8833631)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2773 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3258 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd7ec13f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4814 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7dee0437)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3933 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4299 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1637 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(baf1d064)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1031 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7419803f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3014 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_698 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f476ae9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1428 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1458332)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5877 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(976c63b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5546 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e2b0676)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1049 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3830 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f56a5b86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_619 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e50eebb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3002 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2552 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf50f6cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2059 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f26c589a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1586 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7aaebf1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1905 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd54d5ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2249 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a36b68d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1717 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1786 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85277bd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5652 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f6542d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3758 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(880e14cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3354 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3705 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecf19022)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5412 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eafe3597)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5627 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(191fb36c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2290 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bc34919)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_348 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13bfa7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_797 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8936074)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1070 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_725 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ea4ac36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2460 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1728 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9f67483)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3803 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad078e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5790 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2677 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d09e290d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5889 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e999dddd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4748 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b710a83f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4966 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f16aeed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2297 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46162427)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_696 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84851fb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4896 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4819 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(852bd17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5978 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a59e190)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a79824de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4759 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5375660)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5723 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cab5e8be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1162 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eaaa0d9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2670 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1547 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b0990e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2035 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2517 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5589 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b03d197)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1867 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b186961)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2830 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3537 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4516ac3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3924 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c10d719)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_391 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3014bff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4594 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84c69b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3410 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(337239e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6074 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72d71d83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4435 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d298745)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3053 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a81bf58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1742 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c6940ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3260 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(780b05f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_458 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fad1ffd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5834 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8038da26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1798 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3894ded4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4111 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3a55e7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1591 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2213 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cca505b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2750 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3625d753)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_860 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80a8f305)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97b1de0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3358 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(561b8b76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3462 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70aa9dcd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4547 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(167ce1f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2184 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1dfc885)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3802 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b86d6f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1993 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d9df1de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3976 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3aa37b93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4950 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3349 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(911483dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4075 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12312d2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2284 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3c5bf36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3873 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e7a9d26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1081 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c14bc87e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1782 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9e82e78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3959 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5336 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(941fcab8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4157 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9dcd769)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1776 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba275eff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1856 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39739948)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1062 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(237f6a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5200 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ed82521)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2063 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(783e910b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5587 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf1f41ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3926 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb9f30fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1297 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4206 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_651 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(711a6e8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2489 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f0cd75c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4491 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29fd31bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5517 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(650d082e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1723 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb60e9d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3723 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_663 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e7d1b97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3744 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1660 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(806f7364)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5896 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0f12da6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1895 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71d9f483)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1568 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2294 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_803 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1cfa453)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4962 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8194cc9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_710 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_345 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cfdcfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4278 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7277e66f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3699 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1919 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(721e7b3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5920 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_481 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(688351fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2160 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13d7ac53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3406 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7aa1e172)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2737 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f313c12e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1459 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a962101)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_956 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4228 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3829 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce645ead)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5880 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e9fac35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1580 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1076 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57dce7ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1607 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2808 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ada68189)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3760 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4467 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc697f07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5034 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86f201e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3287 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b2c6124)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3370 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_3157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2768 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8206d29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4917 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3577 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b890b1f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4183 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d2abc3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2013 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f0db8df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4350 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3539 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5955 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e684bf7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4471 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1862 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe5f13f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1992 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bc30e55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2668 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fe01424)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3746 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3f90f88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5296 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24d718f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3166 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee999b87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1530 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1015 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fc651af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4599 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(455d82af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5541 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(190424da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_455 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62795e06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1007 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_656 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4069 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60d134f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6083 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7deffb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_474 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(739e7945)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5060 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b699e09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4449 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cbe6d22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5072 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4188 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d5cb61a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1685 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2187 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e93a71da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4472 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e7e1818)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1084 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3342 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b407a98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4545 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60bf4c5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35e788b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4956 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0cc1f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1687 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76fe371a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2299 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf9e73d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1978 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de4ca397)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2420 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cfc7f9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2246 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe7819be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1328 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b753a8ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5507 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9c6fee4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4359 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32400a7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2275 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6047cf52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1639 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1567 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19142047)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2870 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33782ba2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2395 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b72bb19a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1514 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45c5fa12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3690 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a0b4b43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4373 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c041b590)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2730 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efbd6faf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_669 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db1b1faa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1010 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2167 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4225e009)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_457 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5fdcaa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5882 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1802 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d36675a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1709 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7ca0761)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1910 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3636 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(968dc709)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_330 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f6d32fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2572 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7446c6a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2799 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a5ccb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3888 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cd7255e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_580 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5428 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7461bf0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(741c3d2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1933 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd93d8b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2966 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4362 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3655e6a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2500 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(239510d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6062 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dc2ae97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4038 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1518 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48270edf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4091 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5607 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(928afd55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5371 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(275bb00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_946 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b02c6f75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4648 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(decb907d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3084 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe510702)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_827 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b892f4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4236 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7960a2e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4645 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faccd179)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4035 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4881 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57cd8122)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3952 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a19e98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1847 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1600 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1193 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1023eb98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2685 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_721 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1734 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1ba000d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1505 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3768 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb168eee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1471 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4324 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3034 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b415de29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5400 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1988 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4164 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(613c0b0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3582 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21291691)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2700 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd6fce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5919 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1985 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(178cea19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5391 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c08527bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_473 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b7bee80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_871 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10fb7f21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3167 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d2a5235)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1285 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f967e9bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3543 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c418d2bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4914 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1949 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e872f5e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_844 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb819b8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4451 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3292 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_367 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d54726)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1036 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb140c1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2392 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3776b075)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3536 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36ca3ece)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4589 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12686b6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3473 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5216 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3e136f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1360 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1404 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4682 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c6b265c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5046 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce4697c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5175 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3484 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff526162)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2482 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(817d2996)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4034 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3162 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41f3e20f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5574 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_555 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd185708)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3968 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88428257)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5673 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(559c44d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_832 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19647cbf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1901 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2d91609)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4494 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(781a2613)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4756 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d988ea8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1462 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(374423ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4833 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b3d3efe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5888 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa64d8f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44a969bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3245 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ace7ac92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1794 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a9ccf93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3266 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c27e829f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3345 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e77ad6b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3033 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29fc6285)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3381 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c0a3aba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1682 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f542cf1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4333 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1fc14d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4561 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2930 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64b74339)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4363 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ac76443)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5081 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bd892db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5514 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5911 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5974 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1059 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(589b1f76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_867 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3455 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3245b39c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5131 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70fc116b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3337 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1360f029)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2775 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ca96dc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2245 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6587535)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2358 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ea44b5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3659 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2645 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4436 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d05f3bc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3238 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4665b00f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4271 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d255c5fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_441 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba7370a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3769 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6f58acb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1116 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3863 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99e6507c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3195 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43953da1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4765 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1c7139a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5679 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6092 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98d5edd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3664 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de9eb172)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1313 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4427 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96bdcc12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5841 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1942cb5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5214 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0e471ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4185 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6eab9b15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3432 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fc800bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3074 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4168 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba08d73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3424 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a32f0a19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2295 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85c0fee3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5170 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(457607ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1480 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c952b61d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5360 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(241dd748)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3683 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2523acb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4898 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0d47bbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_775 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7780564d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_682 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4059 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fc89a14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_463 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db9ba861)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2253 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(680db966)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3300 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(365ad8aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5895 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2635 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b936a9ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4005 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5a500fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1814 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(807cd8a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2025 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8b98568)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5703 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f980d2f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2194 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5982 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e228e13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4196 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e986bd8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5596 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb62d04f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5744 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39c1680c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3691 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4695 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3af249f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_547 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(587d486)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3029 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cfde3fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb7c2b05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3028 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42adb1a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3367 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a40b25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4743 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e017bb8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4619 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1e54053)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1369 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3943 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4768 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8af02569)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1450 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8f1387d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3263 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2195dd55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2926 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5672 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cfb481d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1212 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4676 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff1c7258)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4212 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61e44f4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_934 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a257600)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2432 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a0e0f09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_331 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15c9e33f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2169 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4521 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7aca3f84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_418 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1711 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(769d16cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3967 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(890a35ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5786 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1844 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(541156c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2652 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5750 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e9986e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4585 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5948 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c72ea818)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2745 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2886 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5968 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ff0eaac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3049 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4c4405c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1165 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2581 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8155f70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5483 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_621 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c55f55d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5986 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4008ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4591 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3438 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f8a065)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4792 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6aaeb468)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_527 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c03ac8ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1579 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1994 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3840 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e05d87e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4468 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1755 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7cd3fed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1861 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a28f64a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4203 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d5ae90d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3592 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30ab8fa4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4712 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7fbf49b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2363 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1838 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33227aa6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1326 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2953 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3d940bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1833 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8849c4fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1606 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9c9f98d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1434 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be08fe1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3179 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1694 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b416ad6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1278 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(208321e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2836 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a05bf275)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2324 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db7cdd96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5212 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1244 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec32b3c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3630 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63769f5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5953 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b707211)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3333 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4896f25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2403 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c248c967)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4315 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4429 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_585 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f0564c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(586be7ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_859 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f2c5431)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4343 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c41b001)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3087 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6a587d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5303 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3185 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b81e3a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2656 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(268d749e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3206 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbe832e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1210 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69fa017)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5030 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7ee120b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5024 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(143ba796)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5990 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6047 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5c40830)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2835 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a25a2933)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1094 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1201 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7af101f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3091 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(468cec1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4968 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f537cc32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3966 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4ea6c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4907 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5771 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14497212)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2069 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2372aeca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5355 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1038 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2e52301)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5284 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c21808b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2872 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a7e87ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3336 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d536cf83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4608 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64cf600e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3175 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db2c545)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3101 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67b6c7d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3391 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(492277d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5014 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f158713)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1083 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27ac170)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1809 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90050d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1014 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5124 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ebdd48e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1170 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23d5b088)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_629 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3677 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3964 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0bfe4ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1509 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5be6128d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5141 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2461d054)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1691 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ade26640)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5414 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4415950)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c4a3a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1951 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3547fd2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_771 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5015bd30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3700 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e2444e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4392 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fb034eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1981 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1247c15d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1525 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ec43d02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6002 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5b35b21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4960 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b51c705)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_591 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9d3c7b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_814 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1d92f89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1447 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca592ab0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4529 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3307 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4991 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2881 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(503baaa8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2560 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27f1d068)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_572 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7281957)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2895 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68badf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4773 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1463 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96bb874d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1754 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a37aa3f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4926 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa083844)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3727 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98fb3d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1432 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4625dfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2414 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77ec11ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2108 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2906be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3910 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_996 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3224 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3159 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0a769f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_776 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2421 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5a3bb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2960 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa007e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1207 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc2f8beb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2144 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b161d466)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_358 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(138343e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5692 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5544 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bbaf1173)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1448 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a97e349a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1327 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbf00eb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1877 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da2e43e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5238 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9019ccd2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3730 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4357 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6525af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2402 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46af6c1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4655 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a354968)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4047 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5071 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12b81111)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6015 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4464 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2797b85e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1179 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4230 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2167550)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2141 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7657c671)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3135 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(520f079c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5631 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(177b772b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2651 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33c1e939)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4006 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5796 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c50ceaac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2815 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(557291c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1615 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ade6f738)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2060 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43fcf796)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_631 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3007 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45a34a95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1003 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2443 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ede83568)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2903 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(163e2d91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2891 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5722 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9795e30e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2973 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c08d5026)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11b6aa96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6011 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dcedede1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4180 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c98346c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3276 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96926d21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5868 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f0d2190)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3566 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95427f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2977 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35572b55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4930 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd58b528)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_734 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ca2241)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1324 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d2a8ad5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3813 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3785 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a069f78d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3316 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1736 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35043ad7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_877 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be0a8bba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2931 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1a0c712)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6081 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dcf141)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3134 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5226 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0f83796)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3375 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_826 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2985 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d18b8300)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2643 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(300b4a8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5575 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5e9569)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_849 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c873916c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3777 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa272e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1708 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5eddf1c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50e4fd2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2496 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4933c54c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1203 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd171d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5639 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9c6e7ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(463ea659)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2274 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_624 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99ccf6b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2509 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ccf3ebd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5356 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2fc0fbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2792 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13d274de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4242 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c09d9be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3104 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d33b38a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2049 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5199 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5067 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c8be89b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4394 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ea83cc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_453 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(782f87e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2523 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d2d1db5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1111 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c722d5d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3748 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adb19040)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2311 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(beccf062)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5502 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ba99a2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4702 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5be6894d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3199 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eba4f141)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3588 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(782a6d4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_488 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5246dbb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5668 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdaaa72a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5810 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(826dc468)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5840 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0401767)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2704 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1810 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2814 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4414 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(165ae724)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5524 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a61a4bea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1650 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8362b44b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5802 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b86edc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4999 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9acb7952)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1537 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cf14f36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2518 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7ac51ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1663 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f7bbfc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_909 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5251 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1394 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdca3a3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4838 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5255edb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_583 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6a9f45a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1795 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3013318)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2314 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32b0516d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4616 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2171 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7ef80c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_435 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee0e8623)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5118 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6a8c9d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4281 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dcf137af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1100 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3490fe45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_658 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7be5177f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2468 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a808a53c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_810 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf98a3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3908 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_373 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8c26277)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2809 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5833 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2580d5b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5288 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17fa6208)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2713 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c759d762)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2790 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9b3ce6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3486 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5458 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75450b91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4513 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fae33d78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3112 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f586c82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_562 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd4d9f72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2464 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6488c6b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5848 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd38e6e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3764 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4f9caf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2909 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4241 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f020309)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2168 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35336603)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2598 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d908047d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2388 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5620 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eff6d374)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1061 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(caecf886)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3854 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e80806a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5094 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1eacea3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87f9be83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2666 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6e9970d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6038 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6043 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c3126be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1291 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3500 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecb53c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_982 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcd8d5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4329 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af8a8600)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2033 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3628 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_586 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2612161)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_684 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6014 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eae55c82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3306 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1845 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1d18857)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2804 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fed8ee0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_968 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ffb4ef5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3949 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac25197d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2987 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e23844a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1012 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3569 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6e8e270)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5448 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(704775e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1455 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1781 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1183 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5166406)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5055 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e308c3fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1215 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2182ca55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1807 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6095 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a547140e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4211 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4690 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7848cf5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5451 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2110 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(901e72eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5900 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1126 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f636c09f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2349 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(273b20de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2221 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b39f131c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4662 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d016e21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4207 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f7c1d40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5973 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f4debde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2834 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_972 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ceee5c8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_916 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4f92be8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4587 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c7681f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4300 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5022 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fddb77c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_950 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(705007cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4920 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4389 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1535 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c198ed09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3602 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1165aa66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2539 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(338e484c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3718 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b835f53b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5686 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf65935a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4334 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3633e9f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1005 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69505fee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4052 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(964a8735)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3116 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21825144)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5745 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19afc78b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5271 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b674825)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4514 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(484e79a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5560 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1053 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d98eab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1769 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4271950f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1387 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1233 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3201 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2741 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e20c221a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2513 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4ce84d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3147 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b17dfdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2209 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5e78a59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2893 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3435 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(894b952e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3231 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_503 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2deeb2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3026 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aaf1384c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1772 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23e4d992)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5651 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d097b804)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_510 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96ddb71a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2935 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3c8fc47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4369 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f6c6c01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4680 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43eefcaf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5964 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0b875)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3369 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74e9aea3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3991 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80f6ce9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3386 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94a0e2f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1109 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e22f6086)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3782 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44384c53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1444 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de708a04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5476 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed3e3974)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2239 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4daea2eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5678 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(427cb36e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4879 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15099aec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_654 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1e5d3b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4901 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f15d846d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4617 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3852 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6628db51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2553 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b40a313)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1380 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41447f2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a522acd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4498 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af4e9ce6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3678 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed8fde40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2280 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3474 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8857854d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5576 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3817 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f40b6b50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79f5059d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1478 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d315fab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3282 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc80ea61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1178 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b29c5caa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5037 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b55eb3dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6036 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d95931eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2650 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5702 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb5bbbaf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5649 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35731a40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1487 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f02e1c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3850 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56e50597)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2863 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80d81a24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5208 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_608 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5187 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4886 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_813 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a85c33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5209 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1454 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d92435)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2075 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(767980e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2378 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5012 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdb0b287)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1921 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(643d3210)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2644 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(632152de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3646 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fbe612d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_948 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d262bda7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_830 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7d76cde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_967 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2929 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa3663a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1902 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5999 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3939 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d38ceac1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3638 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96eeabcc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1719 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(216ccb8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2437 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4eb642c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2839 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c2ad167)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96f219cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1721 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4696 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da5c1915)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2149 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8da60e57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4975 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62050cfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3572 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a131d522)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2441 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bace6656)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1601 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b672edd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3257 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bef547e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_759 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15c81c6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3688 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(293e071)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3902 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccca6948)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4283 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5737 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4554a38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3942 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4c1382f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3603 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3da8f598)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_637 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b4526ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_875 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb8168a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3657 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e39d98ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6009 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4865ef0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_579 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7331baa5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5387 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4670 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ad6d860)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1338 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4802 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5469 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9043c58b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5083 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4501 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b07f4065)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4319 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9901e7d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5283 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1213 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94d52c66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4027 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67c882e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1640 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5976 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a71efab0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2243 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c03be73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_649 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1294 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a37b90b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4248 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25d9e4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4420 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d449dd56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2272 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1773 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd27e1b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2200 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f82141)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1793 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1b7575d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2528 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68aab53d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2328 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d600b9a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5368 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68363bf3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1479 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e041721a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1684 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0eb28dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5292 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4847 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df9b0b69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3480 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8424aed7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_461 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9aeddca2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5310 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60b2e1d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4189 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9effb938)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6045 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5280 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc2f0316)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_790 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ead206a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5894 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5f9435c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2230 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3809 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(346552db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3841 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5591 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb6f2fe7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3187 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f5440b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1893 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(542cc6aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_817 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33675f1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3279 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4447 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3e1dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1376 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3069 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6093ede7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2605 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26b10acf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2127 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f48b5800)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1774 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37b9f6ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_821 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2762 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_422 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64146fb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4171 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64ba8a90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1974 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2271 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8131ef04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2495 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46175ea8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1647 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7f61fe3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2556 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3489 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a10c9db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_357 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5245e2c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_843 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b75ce7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1243 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7dd730b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5159 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23ab018b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1958 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2e04643)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3050 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2371 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3917 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2ae8870)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_377 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3b7c0f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_196 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e286d50a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1078 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6efc757c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2325 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cac92e4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2759 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1673 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc955384)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3488 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8d4ab20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2602 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7519442)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3868 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34dba21b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4049 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_975 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e23ccdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3601 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eda7e229)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_893 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2f0c880)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1296 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33ba118f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3078 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(180b1da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3409 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6010 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5991 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2734 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3517 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdab9614)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1984 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5365 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(763c6142)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5529 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cad0887b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6085 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(183bdaba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3878 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5941f67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1990 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14684dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5114 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(471db8f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4801 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cd4a757)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3065 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2d641e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2915 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a71af01c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3044 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab684226)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3495 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3531 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f27573ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1991 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9a19898)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1752 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f1689cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3505 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4202248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5021 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4875200b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4678 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c411e5e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3972 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1332 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_978 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82124d3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4378 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2708 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0e0884)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4431 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5134 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdb91af3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2860 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f836b76b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3371 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9304df4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5320 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1642 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(336bf02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2900 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dcead0bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1835 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ffe00be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4609 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9a27d9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2032 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd2c90da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_886 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9c1f390)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4669 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcc8b059)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1922 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f4fdedf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3085 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(740f079d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3896 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6732b3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3610 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed2e2799)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4073 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5482 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb5a8010)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3784 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2571 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5167fde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3155 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5774 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9043957b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1095 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b12ebe82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5693 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(562c9882)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5736 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d548588c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3169 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(590f7a0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5477 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b141bf3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2732 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7807e296)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5630 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34f44a6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2412 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2982 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61aebaa8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5059 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b86083c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5680 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49d8efab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4008 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a693014e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3433 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3510 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73d63c4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2606 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5832 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c42d59c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3608 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f091516c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4857 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(736df8a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_928 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5111 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6469f89a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5695 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e779bd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4984 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59ff9cc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1467 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19b80982)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2974 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72047530)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2256 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e87347e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1358 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_983 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb56f085)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3208 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cfdce38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_952 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8ae6943)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2530 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(136aa091)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2436 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1262 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34b5aa44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2124 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fb49a43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2574 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fed99956)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3145 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc1234d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2992 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_913 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f113f97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df76f06b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1852 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_409 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_889 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1ea4703)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5130 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4399 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5a3ef13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5444 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c54a5efc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4132 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52556c9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2658 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3071 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d803a93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4326 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a7f8059)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5417 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56ef5852)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1189 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e3a0f24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2698 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cca1d63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2334 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af4ba4e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3858 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_415 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(842e5499)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2634 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1449 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b578f83b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3747 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd969604)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5354 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c691b983)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3389 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3695ad2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3252 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3139 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2361 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35292e27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1139 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(142f163d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2399 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81fc24e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3640 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd3b279a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2262 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4576 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3361 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed3b4a0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2083 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a46b36c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4205 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4784 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2313 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5957 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17905fa7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1526 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3153 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5431 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5564 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5298 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18986e50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5789 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff038850)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2946 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b765626)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2540 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1565 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f4cbb48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2343 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88bfcaa5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4983 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2659 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85ec50c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5003 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ee423a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1305 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(121f03f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4121 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c18468a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3247 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86de25f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2542 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e438f1c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1635 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af43b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5648 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95ab95f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4628 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2070 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(133b7906)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1142 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad8eefe7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5907 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b604c26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5240 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c2b0c52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3780 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2579530c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5042 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74263f90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4276 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11a4565)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4964 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(204616dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3530 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2eee967a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5497 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9de25fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1836 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1077 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec8d5fea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5855 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76f02d0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3348 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14d02faa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5234 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac7a72e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2712 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82b33d7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_829 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_862 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b7b12b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2939 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2810 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b027053b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5625e99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2268 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a6f5363)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2123 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4872b5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_670 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3401 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8560caa5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3881 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7e240f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_484 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a0a735d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3025 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e54a3abe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2383 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41554a38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4731 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f237811)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5531 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2a3be7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3816 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15ab0e0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_779 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8abbaf1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2084 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8571e4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1350 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1029a2f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1529 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(235119ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4822 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16965a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1816 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e13663)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4245 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e034110c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4706 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0fb3591)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4385 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b11daa0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2584 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58c37a41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_964 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb87a4cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1561 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb9b45e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3249 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47d53a9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_341 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97d227c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2175 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61605821)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5329 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1784 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2682 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78a10587)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2922 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a90f5a18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4062 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88f8dc86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2066 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2890 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27d08dbf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1043 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_627 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73dd549d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3778 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec090c0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3545 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25e7d18b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5040 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2720 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e3199e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1348 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a15d12e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2729 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77b5bce3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5102 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f18f98f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2072 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e247986)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4463 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2503 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd6c00c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5035 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1025 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1850 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ee86147)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3009 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e291153)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5264 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a49e7e5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1995 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d995e53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef600cd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2430 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76a8fec5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2785 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce72ee70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3137 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f811b2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5489 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6005 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5cb1adb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1965 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b995755)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4072 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2318 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74a4bfa5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4033 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2822 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cef9abe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1975 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edff2e3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5568 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0cb5681)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4560 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2458 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3856 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_564 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fa55b25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4979 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4166 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa1c9bed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_477 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f64cdfcf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2067 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23afa6f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_839 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea18b29a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1096 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7def3c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5276 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbfa3325)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3828 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3851b01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2885 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2a768d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6090 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5839 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1401 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fce9082)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5404 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2220 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc8fe53c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4060 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42dd3015)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1055 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9378903f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4543 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(134231a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_740 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f07c54b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1669 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(343ee801)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3714 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4568 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f16b434a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1783 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5954 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(188a148b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5851 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26b7f0eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4297 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa58a5ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_957 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cc8e158)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1017 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f9543d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4967 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9046f56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_332 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_920 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4094 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44b6e5eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5664 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8517c92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5349 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2133 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_630 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3897 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(558e650f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4057 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6264fe3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5376 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a494201d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3660 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce2f8b83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5947 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84c7feb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1117 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8205882)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5402 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4102 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4971 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2457 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bfdea3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3117 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(985c942f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2551 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3068 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(924eff48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3331 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4146 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4794 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3399 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1715 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51fbc41b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4988 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3265 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9846241)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4607 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7855b078)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3542 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(689789ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1453 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_757 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1938 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea5048d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2142 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_536 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(578dbe49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_879 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17f4ca65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2763 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5613 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7753db82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_515 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39ab6817)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3124 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3501 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f060324b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_421 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f972144d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4673 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df3d0107)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3557 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5103 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(391554f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9caaf9f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4361 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1538 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(251f09f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5167 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1016 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3160 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fde753e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3721 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd47cb00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5975 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bda5162)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_911 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2e06089)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2526 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3600 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1104 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9b9469)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4255 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9af87a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5640 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3163 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2653 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(222ef853)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5121 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2270 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bdc1347)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2475 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4834 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4302 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc23012b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4344 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56380227)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5239 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1722 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1224b9a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5650 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afe11fcc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1926 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1624 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b1d19b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_376 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc3d4fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4288 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8386eec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4158 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3f1e8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_724 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f149afb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_837 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6bf9560)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1227 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b956c669)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_306 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3157b69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5699 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26616b89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3860 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(970aee12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4239 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4760 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70d41a22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4151 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1251 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46d26e16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1152 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4761 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3118 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3143 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f265394f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3679 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5acc9bfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_760 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7fdee73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3734 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12484089)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd9adfc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3931 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bdbc05b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2089 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99642548)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1733 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3468 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4537 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75cd7782)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4327 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2181 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9776db8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1413 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2ae02e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5272 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_745 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2712a354)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4688 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(106d79a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1085 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f07959b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da89ffb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1001 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(931f254)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3725 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2770 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_406 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48cfe32a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5858 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6347f379)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4216 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31bacbd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_758 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed2f2e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2533 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(847f702)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4573 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2259 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(583c739d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3822 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb291941)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2062 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8539373)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3076 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e84cee3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5597 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4207174)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2678 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3812038e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4722 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5512 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9daa0528)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3459 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c40cb18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5057 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22201739)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3811 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0fb8eb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5592 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1778 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3884 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30d082a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2265 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ade9f0a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5822 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3394 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3010 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42a460a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5775 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bbdc38c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5172 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e32133c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5506 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34c6e74c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3617 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4500 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c720dad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3525 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3387 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4873 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3251 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4767 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc2eb4ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2466 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81fbc8b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3228 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5726 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dab54871)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2846 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2746 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb2d1736)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_752 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1241 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d328459)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5328 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab2443ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5557 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a658af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5945 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_570 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4201 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5053 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a61c185)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4855 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3876 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95b10217)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5707 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_480 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef45c7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1864 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(872c6352)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_820 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a75204b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5853 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_554 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3240 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4730fce5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3239 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3227 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1e04bd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2302 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a3fe03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5447 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc87efb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5210 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2684 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc1435e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2191 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3269 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6acb9861)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5534 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_625 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4461 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42a41d41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1612 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2333 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(918aa604)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1934 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbe04cfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3595 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5020 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68326ff5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1947 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7df1c7af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3e48056)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3590 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4af0c2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5221 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0cfa927)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4839 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef9aee23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_470 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4096 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(301c1eb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1764 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1022 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d4cc392)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_955 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3556 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(728392cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4575 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4a3f6c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4099 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92c0ab03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4650 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77a3f1b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_322 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee83fd65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4937 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0514bdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1592 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12e3f7b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5437 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9d9c356)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5361 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2628 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(408e7656)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5980 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9588e34e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4214 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39382ef7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2278 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c524211)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2934 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41f4a860)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1255 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58457bc7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5381 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afcede63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4115 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa22bbe4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1789 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a50d0821)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5734 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5261 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5092 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c788b6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3441 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62288438)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5755 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c54fd2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2821 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bbf8058)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3377 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7518ffe4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2524 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3362 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5457 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4273 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8e674f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3243 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30fae625)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5500 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(814adb36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_387 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61aac666)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5601 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2957 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6708cf45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4815 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7ae71af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4976 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5c50a97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5946 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1412 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86e1f5e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3417 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(142f3fcf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4842 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fc6f651)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2064 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7245bea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2163 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e18de450)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1319 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87e7ff78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4544 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc10fb75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2107 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a039d240)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3515 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2367cf62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5527 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f53a229)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5250 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5473 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7e8f69f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5363 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6ad51fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4174 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(288429cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2573 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(527bed14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2326 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce0a73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5422 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5323e45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3021 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(189072d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1936 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42f92751)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2627 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fabdff6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2469 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2286727d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2599 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63ee2c55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5570 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27bdd7e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4641 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1050 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18982a08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2841 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4c1f328)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3672 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b9aa725)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5343 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5921 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1163 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a138e57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2207 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3da8f055)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4191 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3198 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7be1c2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1341 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cff90e74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3376 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ba291a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5085 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f102d069)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1127 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca04e2db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3326 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1261 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10bd2d90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1024 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14d46a5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4409 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3e9c4fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6050 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbaf01a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3774 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a31110a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3901 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(837dbca6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4380 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2567476b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1482 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2911 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1161b10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4002 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26c3fd8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5486 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e98e4bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2906 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3864e06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_691 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(add21105)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2769 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4644 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5053dae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_469 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_744 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3382 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a5684e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4342 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4310 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e680b99f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1896 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4811 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2663 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0a36c82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5720 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3302 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1097 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84c9a3f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3575 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1033 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3886 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(216f523d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2529 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(422fa863)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2875 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb8a2ef8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5532 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3df1d2ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5565 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3911 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c871cee3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_508 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a38da8b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4473 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b458ed7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1955 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3974 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffd5b7d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2567 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(574c772e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1373 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_535 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1329 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(811a4958)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6101 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dac3dc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2521 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3058441)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3978 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(123d632f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2577 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ee1ccb1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2899 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2464cfa0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5647 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5685 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5316 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b17f9fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2519 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee2c25f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5843 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c32a422)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4330 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d46eea83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2742 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1250 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76a7ee11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1246 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54fc963e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2904 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2bb10c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5622 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b60bec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d00a0980)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5481 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(803f5fce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1310 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89b7bc29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5099 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69aa06ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6042 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80fdafc4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1605 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(942cdcf9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3511 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b45438b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6039 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22215a4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4208 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9ddbc12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5682 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0968c75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2449 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fa25267)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4729 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_711 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(716c966e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4218 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51b1a50b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4068 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2ba1f6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2942 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3017ac2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_917 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fca052b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2755 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a43f28f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4371 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bac79b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3008 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_804 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2472 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(719e8665)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4243 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34a93a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4714 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f040b9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2417 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6699f086)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2674 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(346d46d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4798 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5e6df81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1894 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8251a0c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2051 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd91821c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2118 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44cc5966)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3795 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b70088e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3875 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4470 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(565cd9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5488 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9a83336)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4780 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6db32c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4312 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(103bbb5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3063 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f711269a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1830 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce4e4695)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_540 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28000fc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3041 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88369f8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_694 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5341 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88baed20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3776 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bbfe70f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2427 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1594 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d000ce7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2250 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1195 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e0c7279)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_777 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7edcc65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1702 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc62c838)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2861 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(750b16df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4403 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d19e2a2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_701 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ead9d70c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17c36f2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4781 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51765527)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2478 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c04442d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3579 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ecc25a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2736 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_628 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3db44ed2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_509 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efffd05e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4444 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3328 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8e4cde3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5033 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7afdc28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4079 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5152 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94ecdaa6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2672 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5862 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf7a5ab5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4598 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5395 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(542d11a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4777 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5919697)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3994 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5302 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3642 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddea5b76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4593 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a2ed325)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1839 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25f3905a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4454 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(587039cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_557 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac2dd825)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1268 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a6c78bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1700 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2744 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7d1ee14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5229 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e68a735)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4951 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f22b78d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4649 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(206bdc5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1047 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de338be3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5088 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2476 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(655cc895)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4862 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e21844e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2816 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(906bc69c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_998 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b803ec0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3303 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2791c765)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5798 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1019 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1f8d738)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5740 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f90856)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5347 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(741219d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3491 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fadb848)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5379 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3262 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41096e2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1071 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3364bec2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_692 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d0110d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2594 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a77371d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4025 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10771b54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4918 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c64337ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3932 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1415 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26832fc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4232 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faee6b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_773 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_596 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a740783)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_571 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93bc1724)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3593 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2afa000)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5634 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b56c58b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2401 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4253 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee8299fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3649 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4453 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2119 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff4818de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2624 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd2d8c59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_678 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8be92b34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5076 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32769c0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5654 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad3b877a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_316 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(126a60d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6017 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5d06170)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5179 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(171beb45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3481 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3812 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad1eb7f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1349 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2373 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9be8125)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4694 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5421 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f23b1c9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5319 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5fa5422)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4082 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4519 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb11b0a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1385 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26702761)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_816 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3288 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26e3e668)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4017 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3922 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bb614e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1757 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2368 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(169de992)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5032 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e6ec607)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4762 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4278047)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4957 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77d17fab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3390 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50a5eaf1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5538 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3655 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4946 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a2a0a59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6023 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d48ee71f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2057 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee3daff0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4193 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2289 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63f866f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1066 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4f102e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7313391)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1079 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3074059)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_363 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4586 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93a976b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1231 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6955e887)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_937 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c80815e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2689 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1906 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77496d0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d68e094)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4989 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b062e67c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3990 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17d6f9be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3458 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7105baac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1870 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87b58332)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2760 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb295e10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2844 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b663d94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3439 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a6302f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5207 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ac563f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3833 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(430c11b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b5513ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_396 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4eb87fc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3340 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7f14132)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2298 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1954 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ef03549)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2548 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5721 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2224 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f06e89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4874 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_351 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a510b1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_566 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96c1561)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5090 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb38b118)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2354 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63fcbf24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3728 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(558baf42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3849 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f42d26b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2459 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b30de12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1615f719)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3988 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(858e3318)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2384 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93e63869)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5470 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d1dd2c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4220 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3dbb445)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3248 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(643d6e47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3514 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb2d88be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4155 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(748958d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2531 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4309 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_512 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(888d5ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5966 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dab5daa5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_808 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4890506a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1739 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d54863c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5273 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4aaaed2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4938 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2244 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c8e880)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2554 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c82ca22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_565 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(122f6b9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3641 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edec3f8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3894 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad6eeb1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4613 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d83a9fc7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2962 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33f0e818)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5348 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96e1b5dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1832 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8b7f092)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5390 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34d105)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_314 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2649 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5452 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c49f7af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1045 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2b94fb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2413 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37f1f001)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd2c8f15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_951 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7f31b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4130 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa6fb72f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2442 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb41f4fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_989 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afa02b5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3749 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3176 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe9328c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2614 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_553 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b981b05c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4048 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5b1ff7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2686 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f9f7731)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3151 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1371 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5610 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2a7c434)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2355 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5825 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bc15c10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3158 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34bc313c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5434 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5433 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d697ac02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5466 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbfcd850)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4485 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5341f60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_556 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16403328)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5474 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fad07b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fc1405f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_944 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4733 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13cd9ce2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2140 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80e35ba0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3013 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b627164e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4744 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2404 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3095 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(749974cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3698 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_578 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(315a5056)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1375 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6832d647)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4071 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5245 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(652b3573)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4666 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9842af3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1501 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd3129a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3773 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(272e83a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5729 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9adce45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5938 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3874345e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_963 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d00d3bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1399 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3551 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4261 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e500ee5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4013 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5769a989)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1574 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10bd9f2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4861 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5186284c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2497 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6867cbfd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6029 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b71f5c83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5291 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1599 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9db4ea6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5268 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f20b5ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4813 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4654 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(588f112c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_428 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1269 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9f2dd12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1512 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b3549ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2165 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6289bcfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5657 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87828a82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3831 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2341aa44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1666 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47273e82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1317 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(969f5d33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1611 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9499a24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5225 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93aa40f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3955 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d45b495)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1307 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(598526c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3735 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(febdcc19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_868 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1881 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc937802)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2705 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d279ee0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1367 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4a096c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5688 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3754 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a4cfe57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5987 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(775ffca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4223 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cf3a782)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2721 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45ac00e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1483 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2699 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff53ed11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5110 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2422139f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4457 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(234e348)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2134 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2400 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a02f2889)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1485 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50a86404)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_588 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b0f64ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_444 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe442064)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5367 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0985d38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1931 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_865 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2379 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0140b68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3425 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0b9d782)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4892 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3db9230c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_874 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(336d3f4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4406 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc7da7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2006 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ad6fc09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2296 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e65c4ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1421 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4925 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e23a2cc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2955 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35fd657d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2715 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d1d2b7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2041 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25b74a43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2871 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(704a2551)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2453 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfb280a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2451 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1451 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bab5c9d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5350 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8dfe2b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5449 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae672067)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4882 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46f1dfc4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5971 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21205bd8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5809 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb641502)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2796 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91f0db94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2914 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30788eff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2095 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d918663)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1652 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(759f5159)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5772 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc9ca7f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_976 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93428057)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1638 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4480 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(767c60f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(730113d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5178 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14d30d2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4915 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ab6a212)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2321 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8260679)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_660 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_789 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6271de5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_798 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2660 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43485148)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3598 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f32694d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3246 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a95c8c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1915 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3305 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3396 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(251ed9f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3106 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2740 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed37ac5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3529 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4635 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8aa0ea29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3443 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71cc9f8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2479 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(699e7d81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3051 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(228690e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5218 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b3ea1ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4503 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4726 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b4530d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5105 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcb9ce7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_491 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4caeef8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1887 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c6ba419)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5154 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21b9c005)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_440 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2214 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56c05f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5051 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3770 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_788 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(519de1cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5149 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9f65589)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_372 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4442 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2434fefb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3736 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b6708e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_836 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e0ec6c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3073 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fa60370)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3081 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f7916e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5778 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80b3d1c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5583 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f39107c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1539 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17cb8a7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2771 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0625995)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2990 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2081 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f8ad0bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4316 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5539 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5b06a94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1616 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ed52626)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4339 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0861c13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1834 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(109bbfa3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3192 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4dd49f39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3708 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5752 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2037bde7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6046 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b79ee6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4317 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eee6ea5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4481 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0cbc97d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3193 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99c8f06e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5017 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37708200)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_892 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf38e3c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4066 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcfc4c84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4092 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2818 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(252daeda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2386 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee315726)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2710 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5812 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2661475)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1928 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91af208c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6068 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5025 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3799 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bb74287)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3448 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4320 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9054be6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3520 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af2aaf0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3957 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6057 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5160 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4db3cc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6003 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8af54850)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3622 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1102 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0604d58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5586 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d87cfc16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1750 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85ff57a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3568 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccce5deb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_599 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46807db8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1575 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ebbfc90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1628 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba25dff8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2269 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4301 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6376792)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5228 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1391a8b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2130 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56957473)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1073 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33e2f0dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2791 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2b84a25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5195 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44814c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4112 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3836ebe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1044 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff5ca33c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1197 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62610ef0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2735 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a817c38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5425 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88b46593)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4061 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcba9195)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4231 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0408b7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3453 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bbf8a9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2619 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3861 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6e719c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2409 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_612 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1c6515f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4366 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6995e13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2431 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2014 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2039 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b952f6ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4282 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83b62eaa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4952 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ff424c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2679 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27bd7c60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1196 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4684 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a56cdc4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_842 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74765d43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2028 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a3b51f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2662 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9f01e7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3506 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1524 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd3d4dcc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1366 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4859 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1209 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee10d4ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4440 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee43713)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79a05503)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4476 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1e0723f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1800 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49ae7fe7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1346 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(464da7e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1869 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(794327de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5659 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1150 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92c4956b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2924 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4133 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1272 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3f38a52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5860 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ae8b304)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3407 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5306 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95662fe0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1118 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(661aa7a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4129 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3739 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7caec6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1578 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a0d1db7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1792 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e96c776)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5914 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3366 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6065 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3311 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2e59c8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1046 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19beac4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4095 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b42a56e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1541 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb617c92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5902 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5161 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b08a9178)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1973 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f453429)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3620 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(541fb518)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3132 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(863f073e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3180 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b136d4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5408 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2416 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bb781f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2202 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a27e3f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3182 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_894 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81e92806)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3753 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3c882d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5327 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e53de990)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2711 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba0bae7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_618 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5afd4b51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1224 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_471 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3313831e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5761 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(957126e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2087 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7719ac96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4364 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41c9d40b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_496 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f50f4ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4610 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(749dbe0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1779 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b33d6105)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_748 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba5e117c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2640 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4554 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81200c83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4800 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57132ea2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1452 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ec726f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6060 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecf3be18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2285 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3951 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba1930c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4265 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba6fb343)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_513 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2927 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41542b46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3716 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1b11c4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5604 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c26c8e49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2021 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d307bb88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b6b1bfd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1266 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4150 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7469a4b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2807 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e22334cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4949 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6ac9a31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6099 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ca88122)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6048 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b835094)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1651 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(156f341f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3899 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4faead0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a34ffb22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1982 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78dcabb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_864 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b637d507)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1818 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_824 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ad2d842)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_521 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bc9352b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5338 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_873 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3886f19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3475 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7faae2fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5128 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3705cfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_895 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13c3c7fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5490 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b5ea83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4023 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(626ef657)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3004 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7375109f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3072 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b187f411)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2485 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f9247ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3244 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29d8a790)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2411 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e881f2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3680 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(478ca91e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2452 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5418 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af221a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2007 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2198 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40080e22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5941 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11082284)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1037 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15c03d13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4555 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3949ae6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1322 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4674 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45a7cbb1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4643 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bae4250d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3470 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87b0538d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1543 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f372d0da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3904 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d264c53c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5439 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ea517a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4797 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1e8b912)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4923 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fb9dba2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2483 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a4547d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3122 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5823 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(695e2989)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2578 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4082bd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5133 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2858 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f13b2f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_490 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29f966f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2204 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2430161a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3207 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8f61b4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2031 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5294 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d0e1942)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5943 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c1ba44a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_940 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f35739d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4693 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a618dec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2506 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3707 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56a03a40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1137 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3611 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f97a190d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1420 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2027 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(184cc901)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2219 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72c92ba0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_756 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c19a0d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4532 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c35158a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4487 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1819 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2238 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cae487ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3338 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14b8f4db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4117 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d284354)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2558 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2504 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6150dd57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2831 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be842a17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_697 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36a39535)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2829 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4993edb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3097 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20502c72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5419 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a60d7f59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3479 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9a6c09f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4647 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aad4a8c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4639 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5ee8ba0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5633 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4194 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a993f7b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3400 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3669 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_397 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(444cb7a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5886 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6c66b18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5352 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76bd3e3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_870 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4022 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4796 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9326ff6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6001 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc0bb5a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2754 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1679 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1088 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(965971e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2000 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2647 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4959 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa90f6ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5632 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2d3f445)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4289 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e286784)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4031 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8942b3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5603 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b001e64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5235 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1701ce7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3142 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdeb2017)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4681 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b0a33f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5950 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(809754e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4963 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73844fe6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1325 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e138b13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3472 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c058b7a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4579 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb7427d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1546 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3880 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8ebb5ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4125 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46008419)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5401 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89d94b93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1897 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5122 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3522 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_802 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c74a019d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4533 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21df778f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5027 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c55f6ac0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1302 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3552 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2aaa307)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1511 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2012 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fdbcd12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3493 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb81106f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2440 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76e1d92c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1171 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4557 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dae3aa7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3516 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c752c1bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4942 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d33d9a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2738 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa647f1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3919 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cadaa911)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2020 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5a5db2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1853 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa522001)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3755 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53cf3799)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1200 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5e0d99e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5619 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c44eb08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_791 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38dcff3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_601 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(761b2f04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5578 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2511 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_577 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1634 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ef2d0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5385 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5594 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40e06319)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2217 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1767 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68e28d3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5213 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1999 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63778ced)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5091 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cf2f3b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2502 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5150 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffa74571)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_973 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2917 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67d0919c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5663 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6347ba80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2406 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86368ce0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3103 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13eaeb4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2045 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89317d9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6097 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16de76f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5813 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13ad2836)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5874 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45833346)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5086 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9331fb7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5286 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_708 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5455 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f111ef58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_317 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69744720)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4559 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb477b60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3561 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8611a29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5079 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a36b710d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6094 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e50115c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3079 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91747d43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5748 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9960769)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2576 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6037 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f866224)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1521 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6764cd8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5277 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a271706)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3631 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96478066)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_650 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60e2bff8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2091 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4600a53f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2803 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7f93872)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4323 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d31c8e83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2347 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c764e2d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4335 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(884994c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1499 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adc032cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3980 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efa265a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4020 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8479e3f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2364 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2dee117)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3626 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b65aea8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9aa7d55c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4531 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98df2e99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2611 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(941efd30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3984 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e47c544d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6102 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(879f79f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2617 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9be209c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3869 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a27b0bac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3658 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5fbeb45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5892 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f370f99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_878 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6070 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4810ce3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2317 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45783ba9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4210 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b495c19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4240 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1108 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4912 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3842 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48cc4a0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_342 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fe46ced)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2604 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a256e70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4890 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b0554e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1589 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d82e3f6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5508 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec24ff9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2273 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73aea036)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_765 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(667e2aa1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5066 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a98173f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4723 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(140cf884)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e32fde3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1545 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(402c3d1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2073 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(114e906)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1907 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ebbd9bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2344 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3056 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e6a6e98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1657 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3547 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31ea9358)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3290 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73e32a5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3969 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab6ce8ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1559 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a186b6a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4383 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1134 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5985df18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1946 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3973 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3644 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef447485)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_809 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(296dea86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1402 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2beac267)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1551 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80e9d358)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4710 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70c00437)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4258 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8a8d99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4382 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14cfdb96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1532 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57304025)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5233 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5056 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3da0e62a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4475 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ca2282c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5909 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bef51244)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2040 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1218789a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4812 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21427601)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3958 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3882c67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4459 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26e93cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1944 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59ddd6a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1494 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5264b2dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1858 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(192d1110)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4152 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a28dbd26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4985 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5842 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3818 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1563 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d0fb860)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4878 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5260faf3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5123 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46a80df9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4405 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69f11ec6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3687 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63135215)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2976 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4365 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(431f54b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4277 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de7e134e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c685fb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4845 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4130034b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98843882)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4395 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb81fa87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4701 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2588 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3850940d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6093 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b01e3d25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4753 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ea0fde7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3497 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d40981dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5423 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5465 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b2c3325)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3403 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d34f8a44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3161 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90a771c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_712 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5471 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48123347)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2947 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c42bb1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4450 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6819469c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4803 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8c1154d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5747 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dff34a15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4804 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2c1f16f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2125 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_767 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1716 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_549 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8869319)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2625 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_385 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d50acb11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2937 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1703 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79dc42bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1064 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(331b54c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1161 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b46c9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d5e1796)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1889 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14a44f99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5189 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2375 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ff86d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3000 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46917d6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_686 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d28ca09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5646 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(449a72b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2193 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b55edaa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3956 & _EVAL_5119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4343ce13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
