//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: b21cef66-00f3-44d5-a188-807f478b1270, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_69(
  output        _EVAL,
  input  [31:0] _EVAL_0,
  output        _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  output        _EVAL_4,
  input  [2:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  output [2:0]  _EVAL_7,
  input  [1:0]  _EVAL_8,
  input         _EVAL_9,
  output        _EVAL_10,
  output [31:0] _EVAL_11,
  input  [31:0] _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  output        _EVAL_15,
  output        _EVAL_16,
  output        _EVAL_17,
  input  [29:0] _EVAL_18,
  input         _EVAL_19,
  input         _EVAL_20,
  input         _EVAL_21,
  output        _EVAL_22,
  output [1:0]  _EVAL_23,
  output [2:0]  _EVAL_24,
  output [3:0]  _EVAL_25,
  output [3:0]  _EVAL_26,
  input         _EVAL_27,
  input  [3:0]  _EVAL_28,
  output        _EVAL_29,
  output [2:0]  _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  output [2:0]  _EVAL_33,
  input         _EVAL_34,
  input  [2:0]  _EVAL_35,
  output [2:0]  _EVAL_36,
  input  [3:0]  _EVAL_37,
  output        _EVAL_38,
  input         _EVAL_39,
  output [3:0]  _EVAL_40,
  output [31:0] _EVAL_41,
  input         _EVAL_42,
  input         _EVAL_43,
  input         _EVAL_44,
  input  [2:0]  _EVAL_45,
  input         _EVAL_46,
  output        _EVAL_47,
  output        _EVAL_48,
  input         _EVAL_49,
  output [29:0] _EVAL_50,
  input  [3:0]  _EVAL_51
);
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire [1:0] _EVAL_54;
  wire  _EVAL_55;
  reg  _EVAL_56;
  reg [31:0] _RAND_0;
  wire [2:0] _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire [3:0] _EVAL_61;
  wire  _EVAL_62;
  wire [2:0] _EVAL_63;
  wire  _EVAL_65;
  wire [15:0] _EVAL_66;
  wire [1:0] _EVAL_67;
  wire  _EVAL_68;
  wire [3:0] _EVAL_69;
  wire [1:0] _EVAL_70;
  wire  _EVAL_71;
  wire [1:0] _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire [31:0] _EVAL_76;
  wire [22:0] _EVAL_77;
  wire  _EVAL_78;
  wire [7:0] _EVAL_79;
  reg  _EVAL_80;
  reg [31:0] _RAND_1;
  wire [1:0] _EVAL_81;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_86;
  reg [31:0] _EVAL_87;
  reg [31:0] _RAND_2;
  wire [3:0] _EVAL_88;
  reg  _EVAL_89;
  reg [31:0] _RAND_3;
  wire [3:0] _EVAL_90;
  reg [1:0] _EVAL_91;
  reg [31:0] _RAND_4;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire [7:0] _EVAL_94;
  wire [1:0] _EVAL_95;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire [40:0] _EVAL_100;
  wire [1:0] _EVAL_101;
  wire [1:0] _EVAL_102;
  wire [3:0] _EVAL_103;
  wire  _EVAL_104;
  wire [31:0] _EVAL_105;
  wire  _EVAL_107;
  wire [3:0] _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire [2:0] _EVAL_111;
  wire  _EVAL_112;
  wire [1:0] _EVAL_113;
  wire  _EVAL_114;
  wire [7:0] _EVAL_115;
  wire [3:0] _EVAL_116;
  wire [4:0] _EVAL_117;
  wire [3:0] _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire [1:0] _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  reg [31:0] _EVAL_127;
  reg [31:0] _RAND_5;
  wire [4:0] _EVAL_128;
  reg [2:0] _EVAL_129;
  reg [31:0] _RAND_6;
  wire [7:0] _EVAL_130;
  wire [1:0] _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  reg [2:0] _EVAL_134;
  reg [31:0] _RAND_7;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire [31:0] _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  reg [2:0] _EVAL_140;
  reg [31:0] _RAND_8;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [31:0] _EVAL_143;
  wire [31:0] _EVAL_144;
  wire [86:0] _EVAL_145;
  wire [3:0] _EVAL_146;
  wire [7:0] _EVAL_147;
  wire [1:0] _EVAL_148;
  wire [3:0] _EVAL_149;
  wire [3:0] _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_153;
  wire [31:0] _EVAL_154;
  wire  _EVAL_155;
  wire [1:0] _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_167;
  wire [30:0] _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire [86:0] _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire [3:0] _EVAL_178;
  wire  _EVAL_179;
  wire [1:0] _EVAL_180;
  wire  _EVAL_181;
  wire [3:0] _EVAL_182;
  wire  _EVAL_183;
  wire [1:0] _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire [3:0] _EVAL_187;
  wire [1:0] _EVAL_188;
  wire  _EVAL_189;
  wire [3:0] _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire [3:0] _EVAL_198;
  wire  _EVAL_199;
  wire [29:0] _EVAL_200;
  wire  _EVAL_201;
  wire [7:0] _EVAL_202;
  wire [1:0] _EVAL_203;
  wire  _EVAL_205;
  wire [3:0] _EVAL_206;
  wire [5:0] _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire [1:0] _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  reg  _EVAL_215;
  reg [31:0] _RAND_9;
  wire  _EVAL_216;
  wire [3:0] _EVAL_217;
  wire  _EVAL_218;
  wire [5:0] _EVAL_219;
  wire  _EVAL_221;
  wire [3:0] _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_225;
  wire [6:0] _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire [2:0] _EVAL_230;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire [1:0] _EVAL_236;
  wire [3:0] _EVAL_237;
  wire [31:0] _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire [1:0] _EVAL_245;
  wire  _EVAL_246;
  wire [3:0] _EVAL_247;
  wire [3:0] _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire [4:0] _EVAL_252;
  wire [4:0] _EVAL_253;
  wire  _EVAL_254;
  wire [3:0] _EVAL_255;
  wire  _EVAL_256;
  wire [1:0] _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire [30:0] _EVAL_261;
  wire [22:0] _EVAL_262;
  wire [3:0] _EVAL_263;
  wire [1:0] _EVAL_264;
  wire [2:0] _EVAL_265;
  wire [86:0] _EVAL_266;
  wire  _EVAL_267;
  wire [31:0] _EVAL_268;
  wire  _EVAL_269;
  wire [3:0] _EVAL_270;
  wire [7:0] _EVAL_271;
  wire  _EVAL_273;
  wire [1:0] _EVAL_274;
  wire [3:0] _EVAL_275;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_282;
  wire [5:0] _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire [3:0] _EVAL_291;
  wire  _EVAL_292;
  wire [31:0] _EVAL_293;
  wire [1:0] _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire [31:0] _EVAL_297;
  wire [30:0] _EVAL_300;
  wire [1:0] _EVAL_301;
  reg [5:0] _EVAL_302;
  reg [31:0] _RAND_10;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire [3:0] _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire [86:0] _EVAL_310;
  reg [5:0] _EVAL_311;
  reg [31:0] _RAND_11;
  wire [1:0] _EVAL_312;
  wire  _EVAL_313;
  wire [3:0] _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire [3:0] _EVAL_318;
  wire  _EVAL_319;
  wire [1:0] _EVAL_320;
  wire  _EVAL_321;
  wire  _EVAL_322;
  wire [1:0] _EVAL_323;
  wire [3:0] _EVAL_324;
  wire  _EVAL_325;
  wire [3:0] _EVAL_326;
  wire  _EVAL_327;
  wire  _EVAL_328;
  wire  _EVAL_329;
  wire  _EVAL_330;
  reg  _EVAL_331;
  reg [31:0] _RAND_12;
  wire [3:0] _EVAL_332;
  wire [1:0] _EVAL_333;
  wire  _EVAL_334;
  wire [3:0] _EVAL_335;
  reg [29:0] _EVAL_337;
  reg [31:0] _RAND_13;
  wire [7:0] _EVAL_338;
  wire  _EVAL_339;
  wire [3:0] _EVAL_340;
  wire  _EVAL_341;
  wire  _EVAL_342;
  wire [7:0] _EVAL_343;
  wire  _EVAL_344;
  wire [7:0] _EVAL_345;
  wire [7:0] _EVAL_346;
  wire [1:0] _EVAL_347;
  wire  _EVAL_348;
  wire [3:0] _EVAL_349;
  wire  _EVAL_350;
  wire  _EVAL_351;
  wire  _EVAL_352;
  wire [3:0] _EVAL_353;
  wire  _EVAL_354;
  wire [1:0] _EVAL_355;
  wire [32:0] _EVAL_356;
  reg  _EVAL_358;
  reg [31:0] _RAND_14;
  wire [1:0] _EVAL_359;
  wire  _EVAL_360;
  wire  _EVAL_361;
  reg  _EVAL_363;
  reg [31:0] _RAND_15;
  wire  _EVAL_364;
  wire [7:0] _EVAL_365;
  reg  _EVAL_366;
  reg [31:0] _RAND_16;
  wire [31:0] _EVAL_367;
  wire [3:0] _EVAL_368;
  wire [7:0] _EVAL_369;
  wire [7:0] _EVAL_370;
  wire  _EVAL_371;
  reg  _EVAL_375;
  reg [31:0] _RAND_17;
  wire  _EVAL_376;
  wire  _EVAL_377;
  wire [1:0] _EVAL_378;
  wire  _EVAL_380;
  wire [1:0] _EVAL_381;
  wire [3:0] _EVAL_382;
  wire  _EVAL_383;
  wire  _EVAL_384;
  reg [3:0] _EVAL_385;
  reg [31:0] _RAND_18;
  reg [3:0] _EVAL_386;
  reg [31:0] _RAND_19;
  wire  _EVAL_387;
  wire  _EVAL_388;
  wire  _EVAL_389;
  wire [1:0] _EVAL_390;
  wire  _EVAL_391;
  wire  _EVAL_392;
  wire  _EVAL_393;
  reg  _EVAL_394;
  reg [31:0] _RAND_20;
  wire  _EVAL_395;
  wire [1:0] _EVAL_397;
  wire [3:0] _EVAL_398;
  wire [31:0] _EVAL_399;
  wire  _EVAL_400;
  wire [7:0] _EVAL_401;
  wire [86:0] _EVAL_402;
  wire  _EVAL_403;
  reg [3:0] _EVAL_404;
  reg [31:0] _RAND_21;
  wire [3:0] _EVAL_405;
  wire  _EVAL_406;
  wire  _EVAL_407;
  wire [40:0] _EVAL_408;
  wire [31:0] _EVAL_409;
  wire [1:0] _EVAL_410;
  wire  _EVAL_411;
  wire [3:0] _EVAL_412;
  wire [5:0] _EVAL_414;
  wire [5:0] _EVAL_415;
  wire  _EVAL_416;
  wire  _EVAL_417;
  wire [3:0] _EVAL_418;
  wire [7:0] _EVAL_419;
  wire  _EVAL_420;
  wire [1:0] _EVAL_421;
  wire [2:0] _EVAL_422;
  wire  _EVAL_423;
  wire  _EVAL_424;
  wire [3:0] _EVAL_425;
  wire  _EVAL_426;
  wire [7:0] _EVAL_427;
  wire  _EVAL_428;
  wire  _EVAL_429;
  wire  _EVAL_430;
  wire  _EVAL_431;
  wire [1:0] _EVAL_432;
  wire  _EVAL_433;
  wire  _EVAL_435;
  wire  _EVAL_436;
  wire [7:0] _EVAL_437;
  wire [6:0] _EVAL_438;
  wire [3:0] _EVAL_439;
  wire  _EVAL_440;
  wire  _EVAL_442;
  wire  _EVAL_443;
  wire  _EVAL_444;
  reg  _EVAL_446;
  reg [31:0] _RAND_22;
  wire  _EVAL_447;
  wire  _EVAL_449;
  wire  _EVAL_450;
  wire  _EVAL_451;
  wire  _EVAL_452;
  wire [3:0] _EVAL_453;
  wire  _EVAL_454;
  wire  _EVAL_455;
  wire [3:0] _EVAL_458;
  reg  _EVAL_459;
  reg [31:0] _RAND_23;
  wire [3:0] _EVAL_460;
  wire  _EVAL_461;
  wire  _EVAL_462;
  wire  _EVAL_463;
  wire  _EVAL_464;
  wire  _EVAL_465;
  wire  _EVAL_468;
  wire [3:0] _EVAL_470;
  wire  _EVAL_471;
  wire  _EVAL_473;
  wire  _EVAL_474;
  wire  _EVAL_475;
  wire [5:0] _EVAL_476;
  wire  _EVAL_477;
  wire [3:0] _EVAL_478;
  wire [5:0] _EVAL_479;
  wire [31:0] _EVAL_480;
  wire [1:0] _EVAL_482;
  assign _EVAL_93 = _EVAL_127[27];
  assign _EVAL_274 = _EVAL_57[1:0];
  assign _EVAL_184 = _EVAL_265[1:0];
  assign _EVAL_10 = _EVAL_135 ? _EVAL_183 : _EVAL_44;
  assign _EVAL_211 = ~_EVAL_273;
  assign _EVAL_453 = _EVAL_386 >> _EVAL_359;
  assign _EVAL_476 = _EVAL_438[5:0];
  assign _EVAL_409 = _EVAL_92 ? _EVAL_87 : _EVAL_127;
  assign _EVAL_116 = _EVAL_386 >> _EVAL_397;
  assign _EVAL_243 = _EVAL_425[0];
  assign _EVAL_482 = {_EVAL_286,_EVAL_313};
  assign _EVAL_391 = _EVAL_311 == 6'h0;
  assign _EVAL_320 = {_EVAL_256,_EVAL_278};
  assign _EVAL_131 = {_EVAL_316,_EVAL_403};
  assign _EVAL_52 = _EVAL_275[0];
  assign _EVAL_122 = _EVAL_304 & _EVAL_273;
  assign _EVAL_174 = _EVAL_167 & _EVAL_234;
  assign _EVAL_16 = _EVAL_266[39];
  assign _EVAL_344 = _EVAL_144[31];
  assign _EVAL_418 = _EVAL_326 | _EVAL_190;
  assign _EVAL_86 = _EVAL_385[0];
  assign _EVAL_48 = _EVAL_21 | _EVAL_205;
  assign _EVAL_334 = _EVAL_206[0];
  assign _EVAL_479 = _EVAL_345[7:2];
  assign _EVAL_133 = _EVAL_35[2];
  assign _EVAL_71 = _EVAL_127[24];
  assign _EVAL_429 = _EVAL_439[0];
  assign _EVAL_108 = ~_EVAL_404;
  assign _EVAL_378 = _EVAL_70 | 2'h1;
  assign _EVAL_1 = _EVAL_2 & _EVAL_330;
  assign _EVAL_465 = _EVAL_87[16];
  assign _EVAL_97 = _EVAL_302 == 6'h0;
  assign _EVAL_474 = _EVAL_391 ? _EVAL_176 : _EVAL_363;
  assign _EVAL_29 = _EVAL_135 ? _EVAL_109 : _EVAL_46;
  assign _EVAL_306 = _EVAL_140 == _EVAL_3;
  assign _EVAL_68 = _EVAL_127[13];
  assign _EVAL_164 = _EVAL_91 == 2'h3;
  assign _EVAL_328 = _EVAL_358 | _EVAL_375;
  assign _EVAL_67 = {_EVAL_136,_EVAL_83};
  assign _EVAL_70 = 2'h1 << _EVAL_86;
  assign _EVAL_69 = _EVAL_314 & _EVAL_335;
  assign _EVAL_367 = _EVAL_87 & _EVAL_399;
  assign _EVAL_173 = _EVAL_170 ? _EVAL_145 : 87'h0;
  assign _EVAL_4 = _EVAL_19;
  assign _EVAL_307 = _EVAL_128[3:0];
  assign _EVAL_146 = _EVAL_386 >> _EVAL_381;
  assign _EVAL_463 = _EVAL_150[0];
  assign _EVAL_247 = {_EVAL_249,_EVAL_153,_EVAL_288,_EVAL_417};
  assign _EVAL_312 = {_EVAL_461,_EVAL_194};
  assign _EVAL_92 = _EVAL_201 == _EVAL_99;
  assign _EVAL_423 = _EVAL_255[0];
  assign _EVAL_230 = {{1'd0}, _EVAL_355};
  assign _EVAL_301 = {_EVAL_416,_EVAL_139};
  assign _EVAL_15 = _EVAL_391 ? _EVAL_110 : _EVAL_195;
  assign _EVAL_126 = _EVAL_87[12];
  assign _EVAL_195 = _EVAL_319 | _EVAL_151;
  assign _EVAL_171 = _EVAL_129[2];
  assign _EVAL_371 = 3'h1 == _EVAL_230;
  assign _EVAL_395 = _EVAL_91 == 2'h2;
  assign _EVAL_147 = _EVAL_292 ? 8'hff : 8'h0;
  assign _EVAL_304 = _EVAL_378[1];
  assign _EVAL_415 = _EVAL_226[5:0];
  assign _EVAL_59 = _EVAL_91 != 2'h0;
  assign _EVAL_149 = _EVAL_386 >> _EVAL_156;
  assign _EVAL_316 = _EVAL_87[14];
  assign _EVAL_159 = _EVAL_308 & _EVAL_384;
  assign _EVAL_120 = _EVAL_162 | _EVAL_282;
  assign _EVAL_135 = _EVAL_114 & _EVAL_181;
  assign _EVAL_342 = _EVAL_127[16];
  assign _EVAL_290 = _EVAL_118[0];
  assign _EVAL_163 = _EVAL_198[0];
  assign _EVAL_79 = _EVAL_468 ? 8'hff : 8'h0;
  assign _EVAL_284 = _EVAL_222[0];
  assign _EVAL_393 = _EVAL_87[9];
  assign _EVAL_333 = _EVAL_101 | _EVAL_184;
  assign _EVAL_145 = {_EVAL_111,_EVAL_422,_EVAL_51,_EVAL_6,_EVAL_18,_EVAL_43,_EVAL_14,_EVAL_9,_EVAL_100};
  assign _EVAL_100 = {_EVAL_27,_EVAL_13,_EVAL_31,_EVAL_32,_EVAL_37,_EVAL_12,_EVAL_39};
  assign _EVAL_101 = {_EVAL_53,_EVAL_395};
  assign _EVAL_400 = _EVAL_127[26];
  assign _EVAL_104 = _EVAL_127[2];
  assign _EVAL_426 = _EVAL_91 == 2'h0;
  assign _EVAL_294 = {_EVAL_126,_EVAL_244};
  assign _EVAL_24 = _EVAL_266[86:84];
  assign _EVAL_309 = _EVAL_75 | _EVAL_174;
  assign _EVAL_473 = _EVAL_127[0];
  assign _EVAL_475 = _EVAL_404[0];
  assign _EVAL_462 = _EVAL_87[4];
  assign _EVAL_449 = _EVAL_412[0];
  assign _EVAL_98 = _EVAL_275[3];
  assign _EVAL_200 = _EVAL_18 ^ 30'h2000;
  assign _EVAL_417 = _EVAL_127[7];
  assign _EVAL_142 = _EVAL_391 ? _EVAL_444 : _EVAL_80;
  assign _EVAL_228 = _EVAL_344 == _EVAL_213;
  assign _EVAL_414 = _EVAL_94[7:2];
  assign _EVAL_81 = {_EVAL_295,_EVAL_473};
  assign _EVAL_55 = 3'h3 == _EVAL_230;
  assign _EVAL_319 = _EVAL_80 & _EVAL_395;
  assign _EVAL_138 = _EVAL_181 & _EVAL_260;
  assign _EVAL_401 = _EVAL_262[7:0];
  assign _EVAL_105 = _EVAL_356[31:0];
  assign _EVAL_437 = _EVAL_155 ? 8'hff : 8'h0;
  assign _EVAL = _EVAL_259 & _EVAL_241;
  assign _EVAL_148 = {_EVAL_218,_EVAL_192};
  assign _EVAL_123 = _EVAL_405[0];
  assign _EVAL_383 = _EVAL_87[10];
  assign _EVAL_47 = _EVAL_266[43];
  assign _EVAL_114 = _EVAL_97 & _EVAL_208;
  assign _EVAL_353 = _EVAL_386 >> _EVAL_264;
  assign _EVAL_440 = _EVAL_97 & _EVAL_260;
  assign _EVAL_41 = _EVAL_266[32:1];
  assign _EVAL_427 = _EVAL_223 ? 8'hff : 8'h0;
  assign _EVAL_248 = _EVAL_386 >> _EVAL_410;
  assign _EVAL_419 = _EVAL_77[7:0];
  assign _EVAL_207 = {{5'd0}, _EVAL_193};
  assign _EVAL_26 = _EVAL_28;
  assign _EVAL_390 = {_EVAL_84,_EVAL_350};
  assign _EVAL_295 = _EVAL_87[0];
  assign _EVAL_210 = {_EVAL_443,_EVAL_411};
  assign _EVAL_381 = {_EVAL_471,_EVAL_197};
  assign _EVAL_150 = _EVAL_386 >> _EVAL_294;
  assign _EVAL_99 = _EVAL_228 ? _EVAL_227 : _EVAL_305;
  assign _EVAL_156 = {_EVAL_393,_EVAL_229};
  assign _EVAL_155 = _EVAL_404[1];
  assign _EVAL_266 = _EVAL_402 | _EVAL_173;
  assign _EVAL_124 = {_EVAL_107,_EVAL_417};
  assign _EVAL_110 = _EVAL_395 | _EVAL_53;
  assign _EVAL_213 = _EVAL_480[31];
  assign _EVAL_162 = _EVAL_329 | _EVAL_420;
  assign _EVAL_242 = _EVAL_164 | _EVAL_395;
  assign _EVAL_11 = _EVAL_135 ? _EVAL_127 : _EVAL_0;
  assign _EVAL_112 = _EVAL_87[26];
  assign _EVAL_205 = _EVAL_440 & _EVAL_181;
  assign _EVAL_377 = _EVAL_87[18];
  assign _EVAL_255 = _EVAL_386 >> _EVAL_180;
  assign _EVAL_153 = _EVAL_127[23];
  assign _EVAL_407 = _EVAL_418[0];
  assign _EVAL_338 = _EVAL_98 ? 8'hff : 8'h0;
  assign _EVAL_57 = {_EVAL_333, 1'h0};
  assign _EVAL_410 = {_EVAL_377,_EVAL_141};
  assign _EVAL_125 = _EVAL_389 & _EVAL_97;
  assign _EVAL_464 = _EVAL_387 ? _EVAL_251 : _EVAL_189;
  assign _EVAL_221 = _EVAL_391 ? _EVAL_110 : _EVAL_195;
  assign _EVAL_297 = {_EVAL_147,_EVAL_130,_EVAL_427,_EVAL_202};
  assign _EVAL_72 = {_EVAL_431,_EVAL_78};
  assign _EVAL_132 = _EVAL_61[0];
  assign _EVAL_356 = _EVAL_144 + _EVAL_76;
  assign _EVAL_111 = _EVAL_384 ? 3'h4 : _EVAL_35;
  assign _EVAL_189 = _EVAL_285 ? _EVAL_251 : 1'h1;
  assign _EVAL_234 = _EVAL_273 & _EVAL_121;
  assign _EVAL_73 = _EVAL_418[2];
  assign _EVAL_53 = _EVAL_20 & _EVAL_241;
  assign _EVAL_40 = _EVAL_266[36:33];
  assign _EVAL_109 = _EVAL_56 | _EVAL_46;
  assign _EVAL_128 = {_EVAL_187, 1'h0};
  assign _EVAL_361 = _EVAL_182[0];
  assign _EVAL_428 = _EVAL_105[31];
  assign _EVAL_50 = _EVAL_266[73:44];
  assign _EVAL_340 = _EVAL_386 >> _EVAL_81;
  assign _EVAL_322 = _EVAL_127[6];
  assign _EVAL_421 = {_EVAL_296,_EVAL_288};
  assign _EVAL_137 = ~_EVAL_480;
  assign _EVAL_175 = _EVAL_332[0];
  assign _EVAL_25 = _EVAL_266[80:77];
  assign _EVAL_107 = _EVAL_87[7];
  assign _EVAL_206 = _EVAL_386 >> _EVAL_323;
  assign _EVAL_384 = ~_EVAL_464;
  assign _EVAL_188 = {_EVAL_112,_EVAL_400};
  assign _EVAL_460 = _EVAL_386 >> _EVAL_67;
  assign _EVAL_190 = _EVAL_219[3:0];
  assign _EVAL_246 = _EVAL_87[6];
  assign _EVAL_271 = _EVAL_214 ? 8'hff : 8'h0;
  assign _EVAL_232 = _EVAL_248[0];
  assign _EVAL_203 = {_EVAL_279,_EVAL_93};
  assign _EVAL_154 = {_EVAL_338,_EVAL_365,_EVAL_271,_EVAL_369};
  assign _EVAL_214 = _EVAL_275[1];
  assign _EVAL_259 = _EVAL_49 & _EVAL_474;
  assign _EVAL_277 = 3'h0 == _EVAL_230;
  assign _EVAL_439 = _EVAL_386 >> _EVAL_390;
  assign _EVAL_335 = ~_EVAL_178;
  assign _EVAL_222 = _EVAL_386 >> _EVAL_102;
  assign _EVAL_288 = _EVAL_127[15];
  assign _EVAL_323 = {_EVAL_250,_EVAL_60};
  assign _EVAL_293 = _EVAL_171 ? _EVAL_105 : _EVAL_409;
  assign _EVAL_77 = 23'hff << _EVAL_51;
  assign _EVAL_223 = _EVAL_418[1];
  assign _EVAL_451 = _EVAL_391 ? _EVAL_254 : _EVAL_80;
  assign _EVAL_345 = ~_EVAL_401;
  assign _EVAL_387 = _EVAL_35 == 3'h3;
  assign _EVAL_33 = _EVAL_266[83:81];
  assign _EVAL_236 = ~_EVAL_274;
  assign _EVAL_412 = _EVAL_386 >> _EVAL_301;
  assign _EVAL_250 = _EVAL_87[11];
  assign _EVAL_7 = _EVAL_3;
  assign _EVAL_403 = _EVAL_127[14];
  assign _EVAL_280 = _EVAL_49 & _EVAL_451;
  assign _EVAL_103 = {{1'd0}, _EVAL_63};
  assign _EVAL_382 = _EVAL_386 >> _EVAL_72;
  assign _EVAL_130 = _EVAL_73 ? 8'hff : 8'h0;
  assign _EVAL_76 = _EVAL_171 ? _EVAL_480 : _EVAL_137;
  assign _EVAL_54 = {_EVAL_462,_EVAL_364};
  assign _EVAL_17 = _EVAL_266[0];
  assign _EVAL_408 = {_EVAL_366,_EVAL_394,_EVAL_446,_EVAL_215,_EVAL_348,_EVAL_309,_EVAL_267,_EVAL_120,_EVAL_143,_EVAL_328};
  assign _EVAL_226 = _EVAL_302 - 6'h1;
  assign _EVAL_194 = _EVAL_127[8];
  assign _EVAL_88 = _EVAL_386 >> _EVAL_113;
  assign _EVAL_442 = $signed(_EVAL_300) == 31'sh0;
  assign _EVAL_256 = _EVAL_87[5];
  assign _EVAL_185 = _EVAL_129[1];
  assign _EVAL_305 = _EVAL_185 == _EVAL_344;
  assign _EVAL_267 = _EVAL_162 | _EVAL_289;
  assign _EVAL_425 = _EVAL_386 >> _EVAL_148;
  assign _EVAL_349 = _EVAL_117[3:0];
  assign _EVAL_364 = _EVAL_127[4];
  assign _EVAL_66 = {_EVAL_163,_EVAL_341,_EVAL_435,_EVAL_463,_EVAL_334,_EVAL_123,_EVAL_186,_EVAL_290,_EVAL_115};
  assign _EVAL_192 = _EVAL_127[22];
  assign _EVAL_183 = _EVAL_375 | _EVAL_46;
  assign _EVAL_468 = _EVAL_404[2];
  assign _EVAL_201 = _EVAL_129[0];
  assign _EVAL_180 = {_EVAL_433,_EVAL_452};
  assign _EVAL_263 = _EVAL_283[3:0];
  assign _EVAL_219 = {_EVAL_326, 2'h0};
  assign _EVAL_113 = {_EVAL_199,_EVAL_212};
  assign _EVAL_198 = _EVAL_386 >> _EVAL_421;
  assign _EVAL_117 = {_EVAL_69, 1'h0};
  assign _EVAL_144 = _EVAL_367 | _EVAL_297;
  assign _EVAL_289 = _EVAL_167 & _EVAL_327;
  assign _EVAL_402 = _EVAL_142 ? _EVAL_310 : 87'h0;
  assign _EVAL_262 = 23'hff << _EVAL_28;
  assign _EVAL_330 = ~_EVAL_205;
  assign _EVAL_244 = _EVAL_127[12];
  assign _EVAL_376 = _EVAL_340[0];
  assign _EVAL_36 = _EVAL_266[76:74];
  assign _EVAL_182 = _EVAL_386 >> _EVAL_210;
  assign _EVAL_292 = _EVAL_418[3];
  assign _EVAL_350 = _EVAL_127[1];
  assign _EVAL_258 = {_EVAL_380,_EVAL_71};
  assign _EVAL_406 = _EVAL_458[0];
  assign _EVAL_380 = _EVAL_87[24];
  assign _EVAL_265 = {_EVAL_101, 1'h0};
  assign _EVAL_392 = _EVAL_176 & _EVAL_53;
  assign _EVAL_74 = _EVAL_324[0];
  assign _EVAL_399 = {_EVAL_370,_EVAL_79,_EVAL_437,_EVAL_343};
  assign _EVAL_355 = _EVAL_5[1:0];
  assign _EVAL_327 = _EVAL_211 & _EVAL_287;
  assign _EVAL_187 = _EVAL_247 & _EVAL_335;
  assign _EVAL_365 = _EVAL_119 ? 8'hff : 8'h0;
  assign _EVAL_346 = {_EVAL_284,_EVAL_243,_EVAL_423,_EVAL_58,_EVAL_216,_EVAL_232,_EVAL_352,_EVAL_158};
  assign _EVAL_325 = _EVAL_87[31];
  assign _EVAL_443 = _EVAL_87[28];
  assign _EVAL_254 = _EVAL_236[0];
  assign _EVAL_461 = _EVAL_87[8];
  assign _EVAL_324 = _EVAL_386 >> _EVAL_245;
  assign _EVAL_416 = _EVAL_87[29];
  assign _EVAL_63 = _EVAL_404[3:1];
  assign _EVAL_296 = _EVAL_87[15];
  assign _EVAL_196 = _EVAL_211 & _EVAL_121;
  assign _EVAL_313 = _EVAL_127[20];
  assign _EVAL_351 = _EVAL_237[0];
  assign _EVAL_197 = _EVAL_127[19];
  assign _EVAL_458 = _EVAL_386 >> _EVAL_258;
  assign _EVAL_169 = $signed(_EVAL_261) & 31'sh22002000;
  assign _EVAL_455 = _EVAL_453[0];
  assign _EVAL_94 = ~_EVAL_419;
  assign _EVAL_424 = _EVAL_460[0];
  assign _EVAL_339 = _EVAL_127[25];
  assign _EVAL_269 = _EVAL_464 | _EVAL_426;
  assign _EVAL_167 = _EVAL_378[0];
  assign _EVAL_318 = _EVAL_386 >> _EVAL_95;
  assign _EVAL_251 = _EVAL_233 & _EVAL_442;
  assign _EVAL_444 = _EVAL_254 & _EVAL_395;
  assign _EVAL_283 = {_EVAL_398, 2'h0};
  assign _EVAL_102 = {_EVAL_191,_EVAL_153};
  assign _EVAL_422 = _EVAL_384 ? 3'h0 : _EVAL_5;
  assign _EVAL_119 = _EVAL_275[2];
  assign _EVAL_75 = _EVAL_329 | _EVAL_122;
  assign _EVAL_261 = {1'b0,$signed(_EVAL_200)};
  assign _EVAL_352 = _EVAL_88[0];
  assign _EVAL_433 = _EVAL_87[21];
  assign _EVAL_329 = _EVAL_385 >= 4'h2;
  assign _EVAL_310 = {6'h0,_EVAL_385,_EVAL_140,_EVAL_337,_EVAL_89,_EVAL_331,_EVAL_459,_EVAL_408};
  assign _EVAL_450 = _EVAL_167 & _EVAL_315;
  assign _EVAL_143 = _EVAL_209 ? _EVAL_240 : _EVAL_293;
  assign _EVAL_471 = _EVAL_87[19];
  assign _EVAL_65 = _EVAL_127[10];
  assign _EVAL_240 = {_EVAL_455,_EVAL_424,_EVAL_449,_EVAL_361,_EVAL_351,_EVAL_132,_EVAL_74,_EVAL_406,_EVAL_346,_EVAL_66};
  assign _EVAL_332 = _EVAL_386 >> _EVAL_54;
  assign _EVAL_83 = _EVAL_127[30];
  assign _EVAL_95 = {_EVAL_161,_EVAL_68};
  assign _EVAL_470 = _EVAL_386 >> _EVAL_432;
  assign _EVAL_202 = _EVAL_407 ? 8'hff : 8'h0;
  assign _EVAL_121 = ~_EVAL_287;
  assign _EVAL_279 = _EVAL_87[27];
  assign _EVAL_61 = _EVAL_386 >> _EVAL_188;
  assign _EVAL_436 = _EVAL_353[0];
  assign _EVAL_118 = _EVAL_386 >> _EVAL_312;
  assign _EVAL_347 = {_EVAL_383,_EVAL_65};
  assign _EVAL_176 = _EVAL_236[1];
  assign _EVAL_216 = _EVAL_146[0];
  assign _EVAL_285 = _EVAL_35 == 3'h2;
  assign _EVAL_388 = ~_EVAL_242;
  assign _EVAL_241 = _EVAL_388 & _EVAL_269;
  assign _EVAL_249 = _EVAL_127[31];
  assign _EVAL_300 = _EVAL_169;
  assign _EVAL_30 = _EVAL_135 ? 3'h1 : _EVAL_45;
  assign _EVAL_84 = _EVAL_87[1];
  assign _EVAL_227 = ~_EVAL_428;
  assign _EVAL_38 = _EVAL_266[37];
  assign _EVAL_389 = _EVAL_477 & _EVAL_2;
  assign _EVAL_370 = _EVAL_447 ? 8'hff : 8'h0;
  assign _EVAL_225 = _EVAL_470[0];
  assign _EVAL_179 = _EVAL_270[0];
  assign _EVAL_208 = _EVAL_45 == 3'h0;
  assign _EVAL_360 = _EVAL_87[25];
  assign _EVAL_158 = _EVAL_116[0];
  assign _EVAL_348 = _EVAL_75 | _EVAL_450;
  assign _EVAL_275 = _EVAL_398 | _EVAL_263;
  assign _EVAL_405 = _EVAL_386 >> _EVAL_347;
  assign _EVAL_58 = _EVAL_368[0];
  assign _EVAL_438 = _EVAL_311 - _EVAL_207;
  assign _EVAL_170 = _EVAL_391 ? _EVAL_392 : _EVAL_363;
  assign _EVAL_432 = {_EVAL_246,_EVAL_322};
  assign _EVAL_62 = ~_EVAL_133;
  assign _EVAL_270 = _EVAL_386 >> _EVAL_124;
  assign _EVAL_398 = _EVAL_307 | _EVAL_217;
  assign _EVAL_229 = _EVAL_127[9];
  assign _EVAL_452 = _EVAL_127[21];
  assign _EVAL_321 = 3'h2 == _EVAL_230;
  assign _EVAL_136 = _EVAL_87[30];
  assign _EVAL_253 = {_EVAL_349, 1'h0};
  assign _EVAL_454 = _EVAL_391 & _EVAL_49;
  assign _EVAL_420 = _EVAL_304 & _EVAL_211;
  assign _EVAL_268 = _EVAL_127 & _EVAL_399;
  assign _EVAL_141 = _EVAL_127[18];
  assign _EVAL_343 = _EVAL_475 ? 8'hff : 8'h0;
  assign _EVAL_431 = _EVAL_87[3];
  assign _EVAL_193 = _EVAL_49 & _EVAL_221;
  assign _EVAL_233 = _EVAL_51 <= 4'h2;
  assign _EVAL_291 = _EVAL_386 >> _EVAL_131;
  assign _EVAL_260 = _EVAL_45 == 3'h1;
  assign _EVAL_90 = _EVAL_253[3:0];
  assign _EVAL_218 = _EVAL_87[22];
  assign _EVAL_317 = _EVAL_280 & _EVAL_395;
  assign _EVAL_60 = _EVAL_127[11];
  assign _EVAL_245 = {_EVAL_360,_EVAL_339};
  assign _EVAL_287 = _EVAL_337[0];
  assign _EVAL_315 = _EVAL_273 & _EVAL_287;
  assign _EVAL_212 = _EVAL_127[17];
  assign _EVAL_273 = _EVAL_337[1];
  assign _EVAL_286 = _EVAL_87[20];
  assign _EVAL_217 = _EVAL_252[3:0];
  assign _EVAL_22 = _EVAL_266[42];
  assign _EVAL_397 = {_EVAL_465,_EVAL_342};
  assign _EVAL_252 = {_EVAL_307, 1'h0};
  assign _EVAL_199 = _EVAL_87[17];
  assign _EVAL_447 = _EVAL_404[3];
  assign _EVAL_157 = _EVAL_478[0];
  assign _EVAL_314 = {_EVAL_325,_EVAL_191,_EVAL_296,_EVAL_107};
  assign _EVAL_115 = {_EVAL_179,_EVAL_225,_EVAL_157,_EVAL_175,_EVAL_354,_EVAL_436,_EVAL_429,_EVAL_376};
  assign _EVAL_78 = _EVAL_127[3];
  assign _EVAL_411 = _EVAL_127[28];
  assign _EVAL_23 = _EVAL_8;
  assign _EVAL_326 = _EVAL_349 | _EVAL_90;
  assign _EVAL_282 = _EVAL_167 & _EVAL_196;
  assign _EVAL_359 = {_EVAL_325,_EVAL_249};
  assign _EVAL_139 = _EVAL_127[29];
  assign _EVAL_430 = _EVAL_87[2];
  assign _EVAL_435 = _EVAL_318[0];
  assign _EVAL_172 = _EVAL_45[0];
  assign _EVAL_341 = _EVAL_291[0];
  assign _EVAL_264 = {_EVAL_430,_EVAL_104};
  assign _EVAL_478 = _EVAL_386 >> _EVAL_320;
  assign _EVAL_181 = _EVAL_306 & _EVAL_59;
  assign _EVAL_278 = _EVAL_127[5];
  assign _EVAL_368 = _EVAL_386 >> _EVAL_482;
  assign _EVAL_191 = _EVAL_87[23];
  assign _EVAL_308 = _EVAL_259 & _EVAL_53;
  assign _EVAL_480 = _EVAL_268 | _EVAL_154;
  assign _EVAL_354 = _EVAL_382[0];
  assign _EVAL_161 = _EVAL_87[13];
  assign _EVAL_477 = _EVAL_21 | _EVAL_205;
  assign _EVAL_237 = _EVAL_386 >> _EVAL_203;
  assign _EVAL_151 = _EVAL_363 & _EVAL_53;
  assign _EVAL_369 = _EVAL_52 ? 8'hff : 8'h0;
  assign _EVAL_178 = _EVAL_108 | _EVAL_103;
  assign _EVAL_186 = _EVAL_149[0];
  assign _EVAL_209 = _EVAL_134[0];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_56 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _EVAL_80 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _EVAL_87 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_89 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _EVAL_91 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _EVAL_127 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_129 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _EVAL_134 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _EVAL_140 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _EVAL_215 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _EVAL_302 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _EVAL_311 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _EVAL_331 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _EVAL_337 = _RAND_13[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _EVAL_358 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _EVAL_363 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _EVAL_366 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _EVAL_375 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _EVAL_385 = _RAND_18[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _EVAL_386 = _RAND_19[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _EVAL_394 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _EVAL_404 = _RAND_21[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _EVAL_446 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _EVAL_459 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge _EVAL_34) begin
    if (_EVAL_125) begin
      if (_EVAL_138) begin
        _EVAL_56 <= _EVAL_46;
      end
    end
    if (_EVAL_42) begin
      _EVAL_80 <= 1'h0;
    end else if (_EVAL_391) begin
      _EVAL_80 <= _EVAL_444;
    end
    if (_EVAL_159) begin
      if (_EVAL_426) begin
        _EVAL_87 <= _EVAL_12;
      end
    end
    if (_EVAL_159) begin
      if (_EVAL_426) begin
        _EVAL_89 <= _EVAL_43;
      end
    end
    if (_EVAL_42) begin
      _EVAL_91 <= 2'h0;
    end else if (_EVAL_125) begin
      if (_EVAL_181) begin
        if (_EVAL_260) begin
          _EVAL_91 <= 2'h2;
        end else begin
          _EVAL_91 <= 2'h0;
        end
      end else if (_EVAL_317) begin
        if (_EVAL_395) begin
          _EVAL_91 <= 2'h1;
        end else if (_EVAL_159) begin
          if (_EVAL_426) begin
            _EVAL_91 <= 2'h3;
          end
        end
      end else if (_EVAL_159) begin
        if (_EVAL_426) begin
          _EVAL_91 <= 2'h3;
        end
      end
    end else if (_EVAL_317) begin
      if (_EVAL_395) begin
        _EVAL_91 <= 2'h1;
      end else if (_EVAL_159) begin
        if (_EVAL_426) begin
          _EVAL_91 <= 2'h3;
        end
      end
    end else if (_EVAL_159) begin
      if (_EVAL_426) begin
        _EVAL_91 <= 2'h3;
      end
    end
    if (_EVAL_125) begin
      if (_EVAL_138) begin
        _EVAL_127 <= _EVAL_0;
      end
    end
    if (_EVAL_159) begin
      if (_EVAL_426) begin
        _EVAL_129 <= _EVAL_5;
      end
    end
    if (_EVAL_159) begin
      if (_EVAL_426) begin
        _EVAL_134 <= _EVAL_35;
      end
    end
    if (_EVAL_159) begin
      if (_EVAL_426) begin
        _EVAL_140 <= _EVAL_6;
      end
    end
    if (_EVAL_159) begin
      if (_EVAL_426) begin
        _EVAL_215 <= _EVAL_32;
      end
    end
    if (_EVAL_42) begin
      _EVAL_302 <= 6'h0;
    end else if (_EVAL_389) begin
      if (_EVAL_97) begin
        if (_EVAL_172) begin
          _EVAL_302 <= _EVAL_479;
        end else begin
          _EVAL_302 <= 6'h0;
        end
      end else begin
        _EVAL_302 <= _EVAL_415;
      end
    end
    if (_EVAL_42) begin
      _EVAL_311 <= 6'h0;
    end else if (_EVAL_454) begin
      if (_EVAL_392) begin
        if (_EVAL_62) begin
          _EVAL_311 <= _EVAL_414;
        end else begin
          _EVAL_311 <= 6'h0;
        end
      end else begin
        _EVAL_311 <= 6'h0;
      end
    end else begin
      _EVAL_311 <= _EVAL_476;
    end
    if (_EVAL_159) begin
      if (_EVAL_426) begin
        _EVAL_331 <= _EVAL_14;
      end
    end
    if (_EVAL_159) begin
      if (_EVAL_426) begin
        _EVAL_337 <= _EVAL_18;
      end
    end
    if (_EVAL_159) begin
      if (_EVAL_426) begin
        _EVAL_358 <= _EVAL_39;
      end
    end
    if (_EVAL_42) begin
      _EVAL_363 <= 1'h0;
    end else if (_EVAL_391) begin
      _EVAL_363 <= _EVAL_392;
    end
    if (_EVAL_159) begin
      if (_EVAL_426) begin
        _EVAL_366 <= _EVAL_27;
      end
    end
    if (_EVAL_125) begin
      if (_EVAL_138) begin
        _EVAL_375 <= _EVAL_44;
      end
    end
    if (_EVAL_159) begin
      if (_EVAL_426) begin
        _EVAL_385 <= _EVAL_51;
      end
    end
    if (_EVAL_159) begin
      if (_EVAL_426) begin
        if (_EVAL_321) begin
          _EVAL_386 <= 4'h8;
        end else if (_EVAL_371) begin
          _EVAL_386 <= 4'he;
        end else if (_EVAL_277) begin
          _EVAL_386 <= 4'h6;
        end else if (_EVAL_55) begin
          _EVAL_386 <= 4'hc;
        end else begin
          _EVAL_386 <= 4'h0;
        end
      end
    end
    if (_EVAL_159) begin
      if (_EVAL_426) begin
        _EVAL_394 <= _EVAL_13;
      end
    end
    if (_EVAL_159) begin
      if (_EVAL_426) begin
        _EVAL_404 <= _EVAL_37;
      end
    end
    if (_EVAL_159) begin
      if (_EVAL_426) begin
        _EVAL_446 <= _EVAL_31;
      end
    end
    if (_EVAL_159) begin
      if (_EVAL_426) begin
        _EVAL_459 <= _EVAL_9;
      end
    end
  end
endmodule
